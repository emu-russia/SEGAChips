module ym3438 (  D0_i, D0_o, D0_d, D1_i, D1_o, D1_d, D2_i, D2_o, D2_d, D3_i, D3_o, D3_d, D4_i, D4_o, D4_d, D5_i, D5_o, D5_d, D6_i, D6_o, D6_d, D7_i, D7_o, D7_d, TEST_i, TEST_o, TEST_d, n_IC, n_IRQ, n_CS, n_WR, n_RD, A0, A1, M, MOR_sel, MOL_sel, DAC_8, DAC_7, DAC_6, DAC_5, DAC_4, DAC_3, DAC_2, DAC_1, DAC_0);

	input wire D0_i;
	output wire D0_o;
	output wire D0_d;
	input wire D1_i;
	output wire D1_o;
	output wire D1_d;
	input wire D2_i;
	output wire D2_o;
	output wire D2_d;
	input wire D3_i;
	output wire D3_o;
	output wire D3_d;
	input wire D4_i;
	output wire D4_o;
	output wire D4_d;
	input wire D5_i;
	output wire D5_o;
	output wire D5_d;
	input wire D6_i;
	output wire D6_o;
	output wire D6_d;
	input wire D7_i;
	output wire D7_o;
	output wire D7_d;
	input wire TEST_i;
	output wire TEST_o;
	output wire TEST_d;
	input wire n_IC;
	output wire n_IRQ;
	input wire n_CS;
	input wire n_WR;
	input wire n_RD;
	input wire A0;
	input wire A1;
	input wire M;
	output wire MOR_sel;
	output wire MOL_sel;
	output wire DAC_8;
	output wire DAC_7;
	output wire DAC_6;
	output wire DAC_5;
	output wire DAC_4;
	output wire DAC_3;
	output wire DAC_2;
	output wire DAC_1;
	output wire DAC_0;

	// Wires

	wire w1;
	wire w2;
	wire w3;
	wire w4;
	wire w5;
	wire w6;
	wire w7;
	wire w8;
	wire w9;
	wire w10;
	wire w11;
	wire w12;
	wire w13;
	wire w14;
	wire w15;
	wire w16;
	wire w17;
	wire w18;
	wire w19;
	wire w20;
	wire w21;
	wire w22;
	wire w23;
	wire w24;
	wire w25;
	wire w26;
	wire w27;
	wire w28;
	wire w29;
	wire w30;
	wire w31;
	wire w32;
	wire w33;
	wire w34;
	wire w35;
	wire w36;
	wire w37;
	wire w38;
	wire w39;
	wire w40;
	wire w41;
	wire w42;
	wire w43;
	wire w44;
	wire w45;
	wire w46;
	wire w47;
	wire w48;
	wire w49;
	wire w50;
	wire w51;
	wire w52;
	wire w53;
	wire w54;
	wire w55;
	wire w56;
	wire w57;
	wire w58;
	wire w59;
	wire w60;
	wire w61;
	wire w62;
	wire w63;
	wire w64;
	wire w65;
	wire w66;
	wire w67;
	wire w68;
	wire w69;
	wire w70;
	wire w71;
	wire w72;
	wire w73;
	wire w74;
	wire w75;
	wire w76;
	wire w77;
	wire w78;
	wire w79;
	wire w80;
	wire w81;
	wire w82;
	wire w83;
	wire w84;
	wire w85;
	wire w86;
	wire w87;
	wire w88;
	wire w89;
	wire w90;
	wire w91;
	wire w92;
	wire w93;
	wire w94;
	wire w95;
	wire w96;
	wire w97;
	wire w98;
	wire w99;
	wire w100;
	wire w101;
	wire w102;
	wire w103;
	wire w104;
	wire w105;
	wire w106;
	wire w107;
	wire w108;
	wire w109;
	wire w110;
	wire w111;
	wire w112;
	wire w113;
	wire w114;
	wire w115;
	wire w116;
	wire w117;
	wire w118;
	wire w119;
	wire w120;
	wire w121;
	wire w122;
	wire w123;
	wire w124;
	wire w125;
	wire w126;
	wire w127;
	wire w128;
	wire w129;
	wire w130;
	wire w131;
	wire w132;
	wire w133;
	wire w134;
	wire w135;
	wire w136;
	wire w137;
	wire w138;
	wire w139;
	wire w140;
	wire w141;
	wire w142;
	wire w143;
	wire w144;
	wire w145;
	wire w146;
	wire w147;
	wire w148;
	wire w149;
	wire w150;
	wire w151;
	wire w152;
	wire w153;
	wire w154;
	wire w155;
	wire w156;
	wire w157;
	wire w158;
	wire w159;
	wire w160;
	wire w161;
	wire w162;
	wire w163;
	wire w164;
	wire w165;
	wire w166;
	wire w167;
	wire w168;
	wire w169;
	wire w170;
	wire w171;
	wire w172;
	wire w173;
	wire w174;
	wire w175;
	wire w176;
	wire w177;
	wire w178;
	wire w179;
	wire w180;
	wire w181;
	wire w182;
	wire w183;
	wire w184;
	wire w185;
	wire w186;
	wire w187;
	wire w188;
	wire w189;
	wire w190;
	wire w191;
	wire w192;
	wire w193;
	wire w194;
	wire w195;
	wire w196;
	wire w197;
	wire w198;
	wire w199;
	wire w200;
	wire w201;
	wire w202;
	wire w203;
	wire w204;
	wire w205;
	wire w206;
	wire w207;
	wire w208;
	wire w209;
	wire w210;
	wire w211;
	wire w212;
	wire w213;
	wire w214;
	wire w215;
	wire w216;
	wire w217;
	wire w218;
	wire w219;
	wire w220;
	wire w221;
	wire w222;
	wire w223;
	wire w224;
	wire w225;
	wire w226;
	wire w227;
	wire w228;
	wire w229;
	wire w230;
	wire w231;
	wire w232;
	wire w233;
	wire w234;
	wire w235;
	wire w236;
	wire w237;
	wire w238;
	wire w239;
	wire w240;
	wire w241;
	wire w242;
	wire w243;
	wire w244;
	wire w245;
	wire w246;
	wire w247;
	wire w248;
	wire w249;
	wire w250;
	wire w251;
	wire w252;
	wire w253;
	wire w254;
	wire w255;
	wire w256;
	wire w257;
	wire w258;
	wire w259;
	wire w260;
	wire w261;
	wire w262;
	wire w263;
	wire w264;
	wire w265;
	wire w266;
	wire w267;
	wire w268;
	wire w269;
	wire w270;
	wire w271;
	wire w272;
	wire w273;
	wire w274;
	wire w275;
	wire w276;
	wire w277;
	wire w278;
	wire w279;
	wire w280;
	wire w281;
	wire w282;
	wire w283;
	wire w284;
	wire w285;
	wire w286;
	wire w287;
	wire w288;
	wire w289;
	wire w290;
	wire w291;
	wire w292;
	wire w293;
	wire w294;
	wire w295;
	wire w296;
	wire w297;
	wire w298;
	wire w299;
	wire w300;
	wire w301;
	wire w302;
	wire w303;
	wire w304;
	wire w305;
	wire w306;
	wire w307;
	wire w308;
	wire w309;
	wire w310;
	wire w311;
	wire w312;
	wire w313;
	wire w314;
	wire w315;
	wire w316;
	wire w317;
	wire w318;
	wire w319;
	wire w320;
	wire w321;
	wire w322;
	wire w323;
	wire w324;
	wire w325;
	wire w326;
	wire w327;
	wire w328;
	wire w329;
	wire w330;
	wire w331;
	wire w332;
	wire w333;
	wire w334;
	wire w335;
	wire w336;
	wire w337;
	wire w338;
	wire w339;
	wire w340;
	wire w341;
	wire w342;
	wire w343;
	wire w344;
	wire w345;
	wire w346;
	wire w347;
	wire w348;
	wire w349;
	wire w350;
	wire w351;
	wire w352;
	wire w353;
	wire w354;
	wire w355;
	wire w356;
	wire w357;
	wire w358;
	wire w359;
	wire w360;
	wire w361;
	wire w362;
	wire w363;
	wire w364;
	wire w365;
	wire w366;
	wire w367;
	wire w368;
	wire w369;
	wire w370;
	wire w371;
	wire w372;
	wire w373;
	wire w374;
	wire w375;
	wire w376;
	wire w377;
	wire w378;
	wire w379;
	wire w380;
	wire w381;
	wire w382;
	wire w383;
	wire w384;
	wire w385;
	wire w386;
	wire w387;
	wire w388;
	wire w389;
	wire w390;
	wire w391;
	wire w392;
	wire w393;
	wire w394;
	wire w395;
	wire w396;
	wire w397;
	wire w398;
	wire w399;
	wire w400;
	wire w401;
	wire w402;
	wire w403;
	wire w404;
	wire w405;
	wire w406;
	wire w407;
	wire w408;
	wire w409;
	wire w410;
	wire w411;
	wire w412;
	wire w413;
	wire w414;
	wire w415;
	wire w416;
	wire w417;
	wire w418;
	wire w419;
	wire w420;
	wire w421;
	wire w422;
	wire w423;
	wire w424;
	wire w425;
	wire w426;
	wire w427;
	wire w428;
	wire w429;
	wire w430;
	wire w431;
	wire w432;
	wire w433;
	wire w434;
	wire w435;
	wire w436;
	wire w437;
	wire w438;
	wire w439;
	wire w440;
	wire w441;
	wire w442;
	wire w443;
	wire w444;
	wire w445;
	wire w446;
	wire w447;
	wire w448;
	wire w449;
	wire w450;
	wire w451;
	wire w452;
	wire w453;
	wire w454;
	wire w455;
	wire w456;
	wire w457;
	wire w458;
	wire w459;
	wire w460;
	wire w461;
	wire w462;
	wire w463;
	wire w464;
	wire w465;
	wire w466;
	wire w467;
	wire w468;
	wire w469;
	wire w470;
	wire w471;
	wire w472;
	wire w473;
	wire w474;
	wire w475;
	wire w476;
	wire w477;
	wire w478;
	wire w479;
	wire w480;
	wire w481;
	wire w482;
	wire w483;
	wire w484;
	wire w485;
	wire w486;
	wire w487;
	wire w488;
	wire w489;
	wire w490;
	wire w491;
	wire w492;
	wire w493;
	wire w494;
	wire w495;
	wire w496;
	wire w497;
	wire w498;
	wire w499;
	wire w500;
	wire w501;
	wire w502;
	wire w503;
	wire w504;
	wire w505;
	wire w506;
	wire w507;
	wire w508;
	wire w509;
	wire w510;
	wire w511;
	wire w512;
	wire w513;
	wire w514;
	wire w515;
	wire w516;
	wire w517;
	wire w518;
	wire w519;
	wire w520;
	wire w521;
	wire w522;
	wire w523;
	wire w524;
	wire w525;
	wire w526;
	wire w527;
	wire w528;
	wire w529;
	wire w530;
	wire w531;
	wire w532;
	wire w533;
	wire w534;
	wire w535;
	wire w536;
	wire w537;
	wire w538;
	wire w539;
	wire w540;
	wire w541;
	wire w542;
	wire w543;
	wire w544;
	wire w545;
	wire w546;
	wire w547;
	wire w548;
	wire w549;
	wire w550;
	wire w551;
	wire w552;
	wire w553;
	wire w554;
	wire w555;
	wire w556;
	wire w557;
	wire w558;
	wire w559;
	wire w560;
	wire w561;
	wire w562;
	wire w563;
	wire w564;
	wire w565;
	wire w566;
	wire w567;
	wire w568;
	wire w569;
	wire w570;
	wire w571;
	wire w572;
	wire w573;
	wire w574;
	wire w575;
	wire w576;
	wire w577;
	wire w578;
	wire w579;
	wire w580;
	wire w581;
	wire w582;
	wire w583;
	wire w584;
	wire w585;
	wire w586;
	wire w587;
	wire w588;
	wire w589;
	wire w590;
	wire w591;
	wire w592;
	wire w593;
	wire w594;
	wire w595;
	wire w596;
	wire w597;
	wire w598;
	wire w599;
	wire w600;
	wire w601;
	wire w602;
	wire w603;
	wire w604;
	wire w605;
	wire w606;
	wire w607;
	wire w608;
	wire w609;
	wire w610;
	wire w611;
	wire w612;
	wire w613;
	wire w614;
	wire w615;
	wire w616;
	wire w617;
	wire w618;
	wire w619;
	wire w620;
	wire w621;
	wire w622;
	wire w623;
	wire w624;
	wire w625;
	wire w626;
	wire w627;
	wire w628;
	wire w629;
	wire w630;
	wire w631;
	wire w632;
	wire w633;
	wire w634;
	wire w635;
	wire w636;
	wire w637;
	wire w638;
	wire w639;
	wire w640;
	wire w641;
	wire w642;
	wire w643;
	wire w644;
	wire w645;
	wire w646;
	wire w647;
	wire w648;
	wire w649;
	wire w650;
	wire w651;
	wire w652;
	wire w653;
	wire w654;
	wire w655;
	wire w656;
	wire w657;
	wire w658;
	wire w659;
	wire w660;
	wire w661;
	wire w662;
	wire w663;
	wire w664;
	wire w665;
	wire w666;
	wire w667;
	wire w668;
	wire w669;
	wire w670;
	wire w671;
	wire w672;
	wire w673;
	wire w674;
	wire w675;
	wire w676;
	wire w677;
	wire w678;
	wire w679;
	wire w680;
	wire w681;
	wire w682;
	wire w683;
	wire w684;
	wire w685;
	wire w686;
	wire w687;
	wire w688;
	wire w689;
	wire w690;
	wire w691;
	wire w692;
	wire w693;
	wire w694;
	wire w695;
	wire w696;
	wire w697;
	wire w698;
	wire w699;
	wire w700;
	wire w701;
	wire w702;
	wire w703;
	wire w704;
	wire w705;
	wire w706;
	wire w707;
	wire w708;
	wire w709;
	wire w710;
	wire w711;
	wire w712;
	wire w713;
	wire w714;
	wire w715;
	wire w716;
	wire w717;
	wire w718;
	wire w719;
	wire w720;
	wire w721;
	wire w722;
	wire w723;
	wire w724;
	wire w725;
	wire w726;
	wire w727;
	wire w728;
	wire w729;
	wire w730;
	wire w731;
	wire w732;
	wire w733;
	wire w734;
	wire w735;
	wire w736;
	wire w737;
	wire w738;
	wire w739;
	wire w740;
	wire w741;
	wire w742;
	wire w743;
	wire w744;
	wire w745;
	wire w746;
	wire w747;
	wire w748;
	wire w749;
	wire w750;
	wire w751;
	wire w752;
	wire w753;
	wire w754;
	wire w755;
	wire w756;
	wire w757;
	wire w758;
	wire w759;
	wire w760;
	wire w761;
	wire w762;
	wire w763;
	wire w764;
	wire w765;
	wire w766;
	wire w767;
	wire w768;
	wire w769;
	wire w770;
	wire w771;
	wire w772;
	wire w773;
	wire w774;
	wire w775;
	wire w776;
	wire w777;
	wire w778;
	wire w779;
	wire w780;
	wire w781;
	wire w782;
	wire w783;
	wire w784;
	wire w785;
	wire w786;
	wire w787;
	wire w788;
	wire w789;
	wire w790;
	wire w791;
	wire w792;
	wire w793;
	wire w794;
	wire w795;
	wire w796;
	wire w797;
	wire w798;
	wire w799;
	wire w800;
	wire w801;
	wire w802;
	wire w803;
	wire w804;
	wire w805;
	wire w806;
	wire w807;
	wire w808;
	wire w809;
	wire w810;
	wire w811;
	wire w812;
	wire w813;
	wire w814;
	wire w815;
	wire w816;
	wire w817;
	wire w818;
	wire w819;
	wire w820;
	wire w821;
	wire w822;
	wire w823;
	wire w824;
	wire w825;
	wire w826;
	wire w827;
	wire w828;
	wire w829;
	wire w830;
	wire w831;
	wire w832;
	wire w833;
	wire w834;
	wire w835;
	wire w836;
	wire w837;
	wire w838;
	wire w839;
	wire w840;
	wire w841;
	wire w842;
	wire w843;
	wire w844;
	wire w845;
	wire w846;
	wire w847;
	wire w848;
	wire w849;
	wire w850;
	wire w851;
	wire w852;
	wire w853;
	wire w854;
	wire w855;
	wire w856;
	wire w857;
	wire w858;
	wire w859;
	wire w860;
	wire w861;
	wire w862;
	wire w863;
	wire w864;
	wire w865;
	wire w866;
	wire w867;
	wire w868;
	wire w869;
	wire w870;
	wire w871;
	wire w872;
	wire w873;
	wire w874;
	wire w875;
	wire w876;
	wire w877;
	wire w878;
	wire w879;
	wire w880;
	wire w881;
	wire w882;
	wire w883;
	wire w884;
	wire w885;
	wire w886;
	wire w887;
	wire w888;
	wire w889;
	wire w890;
	wire w891;
	wire w892;
	wire w893;
	wire w894;
	wire w895;
	wire w896;
	wire w897;
	wire w898;
	wire w899;
	wire w900;
	wire w901;
	wire w902;
	wire w903;
	wire w904;
	wire w905;
	wire w906;
	wire w907;
	wire w908;
	wire w909;
	wire w910;
	wire w911;
	wire w912;
	wire w913;
	wire w914;
	wire w915;
	wire w916;
	wire w917;
	wire w918;
	wire w919;
	wire w920;
	wire w921;
	wire w922;
	wire w923;
	wire w924;
	wire w925;
	wire w926;
	wire w927;
	wire w928;
	wire w929;
	wire w930;
	wire w931;
	wire w932;
	wire w933;
	wire w934;
	wire w935;
	wire w936;
	wire w937;
	wire w938;
	wire w939;
	wire w940;
	wire w941;
	wire w942;
	wire w943;
	wire w944;
	wire w945;
	wire w946;
	wire w947;
	wire w948;
	wire w949;
	wire w950;
	wire w951;
	wire w952;
	wire w953;
	wire w954;
	wire w955;
	wire w956;
	wire w957;
	wire w958;
	wire w959;
	wire w960;
	wire w961;
	wire w962;
	wire w963;
	wire w964;
	wire w965;
	wire w966;
	wire w967;
	wire w968;
	wire w969;
	wire w970;
	wire w971;
	wire w972;
	wire w973;
	wire w974;
	wire w975;
	wire w976;
	wire w977;
	wire w978;
	wire w979;
	wire w980;
	wire w981;
	wire w982;
	wire w983;
	wire w984;
	wire w985;
	wire w986;
	wire w987;
	wire w988;
	wire w989;
	wire w990;
	wire w991;
	wire w992;
	wire w993;
	wire w994;
	wire w995;
	wire w996;
	wire w997;
	wire w998;
	wire w999;
	wire w1000;
	wire w1001;
	wire w1002;
	wire w1003;
	wire w1004;
	wire w1005;
	wire w1006;
	wire w1007;
	wire w1008;
	wire w1009;
	wire w1010;
	wire w1011;
	wire w1012;
	wire w1013;
	wire w1014;
	wire w1015;
	wire w1016;
	wire w1017;
	wire w1018;
	wire w1019;
	wire w1020;
	wire w1021;
	wire w1022;
	wire w1023;
	wire w1024;
	wire w1025;
	wire w1026;
	wire w1027;
	wire w1028;
	wire w1029;
	wire w1030;
	wire w1031;
	wire w1032;
	wire w1033;
	wire w1034;
	wire w1035;
	wire w1036;
	wire w1037;
	wire w1038;
	wire w1039;
	wire w1040;
	wire w1041;
	wire w1042;
	wire w1043;
	wire w1044;
	wire w1045;
	wire w1046;
	wire w1047;
	wire w1048;
	wire w1049;
	wire w1050;
	wire w1051;
	wire w1052;
	wire w1053;
	wire w1054;
	wire w1055;
	wire w1056;
	wire w1057;
	wire w1058;
	wire w1059;
	wire w1060;
	wire w1061;
	wire w1062;
	wire w1063;
	wire w1064;
	wire w1065;
	wire w1066;
	wire w1067;
	wire w1068;
	wire w1069;
	wire w1070;
	wire w1071;
	wire w1072;
	wire w1073;
	wire w1074;
	wire w1075;
	wire w1076;
	wire w1077;
	wire w1078;
	wire w1079;
	wire w1080;
	wire w1081;
	wire w1082;
	wire w1083;
	wire w1084;
	wire w1085;
	wire w1086;
	wire w1087;
	wire w1088;
	wire w1089;
	wire w1090;
	wire w1091;
	wire w1092;
	wire w1093;
	wire w1094;
	wire w1095;
	wire w1096;
	wire w1097;
	wire w1098;
	wire w1099;
	wire w1100;
	wire w1101;
	wire w1102;
	wire w1103;
	wire w1104;
	wire w1105;
	wire w1106;
	wire w1107;
	wire w1108;
	wire w1109;
	wire w1110;
	wire w1111;
	wire w1112;
	wire w1113;
	wire w1114;
	wire w1115;
	wire w1116;
	wire w1117;
	wire w1118;
	wire w1119;
	wire w1120;
	wire w1121;
	wire w1122;
	wire w1123;
	wire w1124;
	wire w1125;
	wire w1126;
	wire w1127;
	wire w1128;
	wire w1129;
	wire w1130;
	wire w1131;
	wire w1132;
	wire w1133;
	wire w1134;
	wire w1135;
	wire w1136;
	wire w1137;
	wire w1138;
	wire w1139;
	wire w1140;
	wire w1141;
	wire w1142;
	wire w1143;
	wire w1144;
	wire w1145;
	wire w1146;
	wire w1147;
	wire w1148;
	wire w1149;
	wire w1150;
	wire w1151;
	wire w1152;
	wire w1153;
	wire w1154;
	wire w1155;
	wire w1156;
	wire w1157;
	wire w1158;
	wire w1159;
	wire w1160;
	wire w1161;
	wire w1162;
	wire w1163;
	wire w1164;
	wire w1165;
	wire w1166;
	wire w1167;
	wire w1168;
	wire w1169;
	wire w1170;
	wire w1171;
	wire w1172;
	wire w1173;
	wire w1174;
	wire w1175;
	wire w1176;
	wire w1177;
	wire w1178;
	wire w1179;
	wire w1180;
	wire w1181;
	wire w1182;
	wire w1183;
	wire w1184;
	wire w1185;
	wire w1186;
	wire w1187;
	wire w1188;
	wire w1189;
	wire w1190;
	wire w1191;
	wire w1192;
	wire w1193;
	wire w1194;
	wire w1195;
	wire w1196;
	wire w1197;
	wire w1198;
	wire w1199;
	wire w1200;
	wire w1201;
	wire w1202;
	wire w1203;
	wire w1204;
	wire w1205;
	wire w1206;
	wire w1207;
	wire w1208;
	wire w1209;
	wire w1210;
	wire w1211;
	wire w1212;
	wire w1213;
	wire w1214;
	wire w1215;
	wire w1216;
	wire w1217;
	wire w1218;
	wire w1219;
	wire w1220;
	wire w1221;
	wire w1222;
	wire w1223;
	wire w1224;
	wire w1225;
	wire w1226;
	wire w1227;
	wire w1228;
	wire w1229;
	wire w1230;
	wire w1231;
	wire w1232;
	wire w1233;
	wire w1234;
	wire w1235;
	wire w1236;
	wire w1237;
	wire w1238;
	wire w1239;
	wire w1240;
	wire w1241;
	wire w1242;
	wire w1243;
	wire w1244;
	wire w1245;
	wire w1246;
	wire w1247;
	wire w1248;
	wire w1249;
	wire w1250;
	wire w1251;
	wire w1252;
	wire w1253;
	wire w1254;
	wire w1255;
	wire w1256;
	wire w1257;
	wire w1258;
	wire w1259;
	wire w1260;
	wire w1261;
	wire w1262;
	wire w1263;
	wire w1264;
	wire w1265;
	wire w1266;
	wire w1267;
	wire w1268;
	wire w1269;
	wire w1270;
	wire w1271;
	wire w1272;
	wire w1273;
	wire w1274;
	wire w1275;
	wire w1276;
	wire w1277;
	wire w1278;
	wire w1279;
	wire w1280;
	wire w1281;
	wire w1282;
	wire w1283;
	wire w1284;
	wire w1285;
	wire w1286;
	wire w1287;
	wire w1288;
	wire w1289;
	wire w1290;
	wire w1291;
	wire w1292;
	wire w1293;
	wire w1294;
	wire w1295;
	wire w1296;
	wire w1297;
	wire w1298;
	wire w1299;
	wire w1300;
	wire w1301;
	wire w1302;
	wire w1303;
	wire w1304;
	wire w1305;
	wire w1306;
	wire w1307;
	wire w1308;
	wire w1309;
	wire w1310;
	wire w1311;
	wire w1312;
	wire w1313;
	wire w1314;
	wire w1315;
	wire w1316;
	wire w1317;
	wire w1318;
	wire w1319;
	wire w1320;
	wire w1321;
	wire w1322;
	wire w1323;
	wire w1324;
	wire w1325;
	wire w1326;
	wire w1327;
	wire w1328;
	wire w1329;
	wire w1330;
	wire w1331;
	wire w1332;
	wire w1333;
	wire w1334;
	wire w1335;
	wire w1336;
	wire w1337;
	wire w1338;
	wire w1339;
	wire w1340;
	wire w1341;
	wire w1342;
	wire w1343;
	wire w1344;
	wire w1345;
	wire w1346;
	wire w1347;
	wire w1348;
	wire w1349;
	wire w1350;
	wire w1351;
	wire w1352;
	wire w1353;
	wire w1354;
	wire w1355;
	wire w1356;
	wire w1357;
	wire w1358;
	wire w1359;
	wire w1360;
	wire w1361;
	wire w1362;
	wire w1363;
	wire w1364;
	wire w1365;
	wire w1366;
	wire w1367;
	wire w1368;
	wire w1369;
	wire w1370;
	wire w1371;
	wire w1372;
	wire w1373;
	wire w1374;
	wire w1375;
	wire w1376;
	wire w1377;
	wire w1378;
	wire w1379;
	wire w1380;
	wire w1381;
	wire w1382;
	wire w1383;
	wire w1384;
	wire w1385;
	wire w1386;
	wire w1387;
	wire w1388;
	wire w1389;
	wire w1390;
	wire w1391;
	wire w1392;
	wire w1393;
	wire w1394;
	wire w1395;
	wire w1396;
	wire w1397;
	wire w1398;
	wire w1399;
	wire w1400;
	wire w1401;
	wire w1402;
	wire w1403;
	wire w1404;
	wire w1405;
	wire w1406;
	wire w1407;
	wire w1408;
	wire w1409;
	wire w1410;
	wire w1411;
	wire w1412;
	wire w1413;
	wire w1414;
	wire w1415;
	wire w1416;
	wire w1417;
	wire w1418;
	wire w1419;
	wire w1420;
	wire w1421;
	wire w1422;
	wire w1423;
	wire w1424;
	wire w1425;
	wire w1426;
	wire w1427;
	wire w1428;
	wire w1429;
	wire w1430;
	wire w1431;
	wire w1432;
	wire w1433;
	wire w1434;
	wire w1435;
	wire w1436;
	wire w1437;
	wire w1438;
	wire w1439;
	wire w1440;
	wire w1441;
	wire w1442;
	wire w1443;
	wire w1444;
	wire w1445;
	wire w1446;
	wire w1447;
	wire w1448;
	wire w1449;
	wire w1450;
	wire w1451;
	wire w1452;
	wire w1453;
	wire w1454;
	wire w1455;
	wire w1456;
	wire w1457;
	wire w1458;
	wire w1459;
	wire w1460;
	wire w1461;
	wire w1462;
	wire w1463;
	wire w1464;
	wire w1465;
	wire w1466;
	wire w1467;
	wire w1468;
	wire w1469;
	wire w1470;
	wire w1471;
	wire w1472;
	wire w1473;
	wire w1474;
	wire w1475;
	wire w1476;
	wire w1477;
	wire w1478;
	wire w1479;
	wire w1480;
	wire w1481;
	wire w1482;
	wire w1483;
	wire w1484;
	wire w1485;
	wire w1486;
	wire w1487;
	wire w1488;
	wire w1489;
	wire w1490;
	wire w1491;
	wire w1492;
	wire w1493;
	wire w1494;
	wire w1495;
	wire w1496;
	wire w1497;
	wire w1498;
	wire w1499;
	wire w1500;
	wire w1501;
	wire w1502;
	wire w1503;
	wire w1504;
	wire w1505;
	wire w1506;
	wire w1507;
	wire w1508;
	wire w1509;
	wire w1510;
	wire w1511;
	wire w1512;
	wire w1513;
	wire w1514;
	wire w1515;
	wire w1516;
	wire w1517;
	wire w1518;
	wire w1519;
	wire w1520;
	wire w1521;
	wire w1522;
	wire w1523;
	wire w1524;
	wire w1525;
	wire w1526;
	wire w1527;
	wire w1528;
	wire w1529;
	wire w1530;
	wire w1531;
	wire w1532;
	wire w1533;
	wire w1534;
	wire w1535;
	wire w1536;
	wire w1537;
	wire w1538;
	wire w1539;
	wire w1540;
	wire w1541;
	wire w1542;
	wire w1543;
	wire w1544;
	wire w1545;
	wire w1546;
	wire w1547;
	wire w1548;
	wire w1549;
	wire w1550;
	wire w1551;
	wire w1552;
	wire w1553;
	wire w1554;
	wire w1555;
	wire w1556;
	wire w1557;
	wire w1558;
	wire w1559;
	wire w1560;
	wire w1561;
	wire w1562;
	wire w1563;
	wire w1564;
	wire w1565;
	wire w1566;
	wire w1567;
	wire w1568;
	wire w1569;
	wire w1570;
	wire w1571;
	wire w1572;
	wire w1573;
	wire w1574;
	wire w1575;
	wire w1576;
	wire w1577;
	wire w1578;
	wire w1579;
	wire w1580;
	wire w1581;
	wire w1582;
	wire w1583;
	wire w1584;
	wire w1585;
	wire w1586;
	wire w1587;
	wire w1588;
	wire w1589;
	wire w1590;
	wire w1591;
	wire w1592;
	wire w1593;
	wire w1594;
	wire w1595;
	wire w1596;
	wire w1597;
	wire w1598;
	wire w1599;
	wire w1600;
	wire w1601;
	wire w1602;
	wire w1603;
	wire w1604;
	wire w1605;
	wire w1606;
	wire w1607;
	wire w1608;
	wire w1609;
	wire w1610;
	wire w1611;
	wire w1612;
	wire w1613;
	wire w1614;
	wire w1615;
	wire w1616;
	wire w1617;
	wire w1618;
	wire w1619;
	wire w1620;
	wire w1621;
	wire w1622;
	wire w1623;
	wire w1624;
	wire w1625;
	wire w1626;
	wire w1627;
	wire w1628;
	wire w1629;
	wire w1630;
	wire w1631;
	wire w1632;
	wire w1633;
	wire w1634;
	wire w1635;
	wire w1636;
	wire w1637;
	wire w1638;
	wire w1639;
	wire w1640;
	wire w1641;
	wire w1642;
	wire w1643;
	wire w1644;
	wire w1645;
	wire w1646;
	wire w1647;
	wire w1648;
	wire w1649;
	wire w1650;
	wire w1651;
	wire w1652;
	wire w1653;
	wire w1654;
	wire w1655;
	wire w1656;
	wire w1657;
	wire w1658;
	wire w1659;
	wire w1660;
	wire w1661;
	wire w1662;
	wire w1663;
	wire w1664;
	wire w1665;
	wire w1666;
	wire w1667;
	wire w1668;
	wire w1669;
	wire w1670;
	wire w1671;
	wire w1672;
	wire w1673;
	wire w1674;
	wire w1675;
	wire w1676;
	wire w1677;
	wire w1678;
	wire w1679;
	wire w1680;
	wire w1681;
	wire w1682;
	wire w1683;
	wire w1684;
	wire w1685;
	wire w1686;
	wire w1687;
	wire w1688;
	wire w1689;
	wire w1690;
	wire w1691;
	wire w1692;
	wire w1693;
	wire w1694;
	wire w1695;
	wire w1696;
	wire w1697;
	wire w1698;
	wire w1699;
	wire w1700;
	wire w1701;
	wire w1702;
	wire w1703;
	wire w1704;
	wire w1705;
	wire w1706;
	wire w1707;
	wire w1708;
	wire w1709;
	wire w1710;
	wire w1711;
	wire w1712;
	wire w1713;
	wire w1714;
	wire w1715;
	wire w1716;
	wire w1717;
	wire w1718;
	wire w1719;
	wire w1720;
	wire w1721;
	wire w1722;
	wire w1723;
	wire w1724;
	wire w1725;
	wire w1726;
	wire w1727;
	wire w1728;
	wire w1729;
	wire w1730;
	wire w1731;
	wire w1732;
	wire w1733;
	wire w1734;
	wire w1735;
	wire w1736;
	wire w1737;
	wire w1738;
	wire w1739;
	wire w1740;
	wire w1741;
	wire w1742;
	wire w1743;
	wire w1744;
	wire w1745;
	wire w1746;
	wire w1747;
	wire w1748;
	wire w1749;
	wire w1750;
	wire w1751;
	wire w1752;
	wire w1753;
	wire w1754;
	wire w1755;
	wire w1756;
	wire w1757;
	wire w1758;
	wire w1759;
	wire w1760;
	wire w1761;
	wire w1762;
	wire w1763;
	wire w1764;
	wire w1765;
	wire w1766;
	wire w1767;
	wire w1768;
	wire w1769;
	wire w1770;
	wire w1771;
	wire w1772;
	wire w1773;
	wire w1774;
	wire w1775;
	wire w1776;
	wire w1777;
	wire w1778;
	wire w1779;
	wire w1780;
	wire w1781;
	wire w1782;
	wire w1783;
	wire w1784;
	wire w1785;
	wire w1786;
	wire w1787;
	wire w1788;
	wire w1789;
	wire w1790;
	wire w1791;
	wire w1792;
	wire w1793;
	wire w1794;
	wire w1795;
	wire w1796;
	wire w1797;
	wire w1798;
	wire w1799;
	wire w1800;
	wire w1801;
	wire w1802;
	wire w1803;
	wire w1804;
	wire w1805;
	wire w1806;
	wire w1807;
	wire w1808;
	wire w1809;
	wire w1810;
	wire w1811;
	wire w1812;
	wire w1813;
	wire w1814;
	wire w1815;
	wire w1816;
	wire w1817;
	wire w1818;
	wire w1819;
	wire w1820;
	wire w1821;
	wire w1822;
	wire w1823;
	wire w1824;
	wire w1825;
	wire w1826;
	wire w1827;
	wire w1828;
	wire w1829;
	wire w1830;
	wire w1831;
	wire w1832;
	wire w1833;
	wire w1834;
	wire w1835;
	wire w1836;
	wire w1837;
	wire w1838;
	wire w1839;
	wire w1840;
	wire w1841;
	wire w1842;
	wire w1843;
	wire w1844;
	wire w1845;
	wire w1846;
	wire w1847;
	wire w1848;
	wire w1849;
	wire w1850;
	wire w1851;
	wire w1852;
	wire w1853;
	wire w1854;
	wire w1855;
	wire w1856;
	wire w1857;
	wire w1858;
	wire w1859;
	wire w1860;
	wire w1861;
	wire w1862;
	wire w1863;
	wire w1864;
	wire w1865;
	wire w1866;
	wire w1867;
	wire w1868;
	wire w1869;
	wire w1870;
	wire w1871;
	wire w1872;
	wire w1873;
	wire w1874;
	wire w1875;
	wire w1876;
	wire w1877;
	wire w1878;
	wire w1879;
	wire w1880;
	wire w1881;
	wire w1882;
	wire w1883;
	wire w1884;
	wire w1885;
	wire w1886;
	wire w1887;
	wire w1888;
	wire w1889;
	wire w1890;
	wire w1891;
	wire w1892;
	wire w1893;
	wire w1894;
	wire w1895;
	wire w1896;
	wire w1897;
	wire w1898;
	wire w1899;
	wire w1900;
	wire w1901;
	wire w1902;
	wire w1903;
	wire w1904;
	wire w1905;
	wire w1906;
	wire w1907;
	wire w1908;
	wire w1909;
	wire w1910;
	wire w1911;
	wire w1912;
	wire w1913;
	wire w1914;
	wire w1915;
	wire w1916;
	wire w1917;
	wire w1918;
	wire w1919;
	wire w1920;
	wire w1921;
	wire w1922;
	wire w1923;
	wire w1924;
	wire w1925;
	wire w1926;
	wire w1927;
	wire w1928;
	wire w1929;
	wire w1930;
	wire w1931;
	wire w1932;
	wire w1933;
	wire w1934;
	wire w1935;
	wire w1936;
	wire w1937;
	wire w1938;
	wire w1939;
	wire w1940;
	wire w1941;
	wire w1942;
	wire w1943;
	wire w1944;
	wire w1945;
	wire w1946;
	wire w1947;
	wire w1948;
	wire w1949;
	wire w1950;
	wire w1951;
	wire w1952;
	wire w1953;
	wire w1954;
	wire w1955;
	wire w1956;
	wire w1957;
	wire w1958;
	wire w1959;
	wire w1960;
	wire w1961;
	wire w1962;
	wire w1963;
	wire w1964;
	wire w1965;
	wire w1966;
	wire w1967;
	wire w1968;
	wire w1969;
	wire w1970;
	wire w1971;
	wire w1972;
	wire w1973;
	wire w1974;
	wire w1975;
	wire w1976;
	wire w1977;
	wire w1978;
	wire w1979;
	wire w1980;
	wire w1981;
	wire w1982;
	wire w1983;
	wire w1984;
	wire w1985;
	wire w1986;
	wire w1987;
	wire w1988;
	wire w1989;
	wire w1990;
	wire w1991;
	wire w1992;
	wire w1993;
	wire w1994;
	wire w1995;
	wire w1996;
	wire w1997;
	wire w1998;
	wire w1999;
	wire w2000;
	wire w2001;
	wire w2002;
	wire w2003;
	wire w2004;
	wire w2005;
	wire w2006;
	wire w2007;
	wire w2008;
	wire w2009;
	wire w2010;
	wire w2011;
	wire w2012;
	wire w2013;
	wire w2014;
	wire w2015;
	wire w2016;
	wire w2017;
	wire w2018;
	wire w2019;
	wire w2020;
	wire w2021;
	wire w2022;
	wire w2023;
	wire w2024;
	wire w2025;
	wire w2026;
	wire w2027;
	wire w2028;
	wire w2029;
	wire w2030;
	wire w2031;
	wire w2032;
	wire w2033;
	wire w2034;
	wire w2035;
	wire w2036;
	wire w2037;
	wire w2038;
	wire w2039;
	wire w2040;
	wire w2041;
	wire w2042;
	wire w2043;
	wire w2044;
	wire w2045;
	wire w2046;
	wire w2047;
	wire w2048;
	wire w2049;
	wire w2050;
	wire w2051;
	wire w2052;
	wire w2053;
	wire w2054;
	wire w2055;
	wire w2056;
	wire w2057;
	wire w2058;
	wire w2059;
	wire w2060;
	wire w2061;
	wire w2062;
	wire w2063;
	wire w2064;
	wire w2065;
	wire w2066;
	wire w2067;
	wire w2068;
	wire w2069;
	wire w2070;
	wire w2071;
	wire w2072;
	wire w2073;
	wire w2074;
	wire w2075;
	wire w2076;
	wire w2077;
	wire w2078;
	wire w2079;
	wire w2080;
	wire w2081;
	wire w2082;
	wire w2083;
	wire w2084;
	wire w2085;
	wire w2086;
	wire w2087;
	wire w2088;
	wire w2089;
	wire w2090;
	wire w2091;
	wire w2092;
	wire w2093;
	wire w2094;
	wire w2095;
	wire w2096;
	wire w2097;
	wire w2098;
	wire w2099;
	wire w2100;
	wire w2101;
	wire w2102;
	wire w2103;
	wire w2104;
	wire w2105;
	wire w2106;
	wire w2107;
	wire w2108;
	wire w2109;
	wire w2110;
	wire w2111;
	wire w2112;
	wire w2113;
	wire w2114;
	wire w2115;
	wire w2116;
	wire w2117;
	wire w2118;
	wire w2119;
	wire w2120;
	wire w2121;
	wire w2122;
	wire w2123;
	wire w2124;
	wire w2125;
	wire w2126;
	wire w2127;
	wire w2128;
	wire w2129;
	wire w2130;
	wire w2131;
	wire w2132;
	wire w2133;
	wire w2134;
	wire w2135;
	wire w2136;
	wire w2137;
	wire w2138;
	wire w2139;
	wire w2140;
	wire w2141;
	wire w2142;
	wire w2143;
	wire w2144;
	wire w2145;
	wire w2146;
	wire w2147;
	wire w2148;
	wire w2149;
	wire w2150;
	wire w2151;
	wire w2152;
	wire w2153;
	wire w2154;
	wire w2155;
	wire w2156;
	wire w2157;
	wire w2158;
	wire w2159;
	wire w2160;
	wire w2161;
	wire w2162;
	wire w2163;
	wire w2164;
	wire w2165;
	wire w2166;
	wire w2167;
	wire w2168;
	wire w2169;
	wire w2170;
	wire w2171;
	wire w2172;
	wire w2173;
	wire w2174;
	wire w2175;
	wire w2176;
	wire w2177;
	wire w2178;
	wire w2179;
	wire w2180;
	wire w2181;
	wire w2182;
	wire w2183;
	wire w2184;
	wire w2185;
	wire w2186;
	wire w2187;
	wire w2188;
	wire w2189;
	wire w2190;
	wire w2191;
	wire w2192;
	wire w2193;
	wire w2194;
	wire w2195;
	wire w2196;
	wire w2197;
	wire w2198;
	wire w2199;
	wire w2200;
	wire w2201;
	wire w2202;
	wire w2203;
	wire w2204;
	wire w2205;
	wire w2206;
	wire w2207;
	wire w2208;
	wire w2209;
	wire w2210;
	wire w2211;
	wire w2212;
	wire w2213;
	wire w2214;
	wire w2215;
	wire w2216;
	wire w2217;
	wire w2218;
	wire w2219;
	wire w2220;
	wire w2221;
	wire w2222;
	wire w2223;
	wire w2224;
	wire w2225;
	wire w2226;
	wire w2227;
	wire w2228;
	wire w2229;
	wire w2230;
	wire w2231;
	wire w2232;
	wire w2233;
	wire w2234;
	wire w2235;
	wire w2236;
	wire w2237;
	wire w2238;
	wire w2239;
	wire w2240;
	wire w2241;
	wire w2242;
	wire w2243;
	wire w2244;
	wire w2245;
	wire w2246;
	wire w2247;
	wire w2248;
	wire w2249;
	wire w2250;
	wire w2251;
	wire w2252;
	wire w2253;
	wire w2254;
	wire w2255;
	wire w2256;
	wire w2257;
	wire w2258;
	wire w2259;
	wire w2260;
	wire w2261;
	wire w2262;
	wire w2263;
	wire w2264;
	wire w2265;
	wire w2266;
	wire w2267;
	wire w2268;
	wire w2269;
	wire w2270;
	wire w2271;
	wire w2272;
	wire w2273;
	wire w2274;
	wire w2275;
	wire w2276;
	wire w2277;
	wire w2278;
	wire w2279;
	wire w2280;
	wire w2281;
	wire w2282;
	wire w2283;
	wire w2284;
	wire w2285;
	wire w2286;
	wire w2287;
	wire w2288;
	wire w2289;
	wire w2290;
	wire w2291;
	wire w2292;
	wire w2293;
	wire w2294;
	wire w2295;
	wire w2296;
	wire w2297;
	wire w2298;
	wire w2299;
	wire w2300;
	wire w2301;
	wire w2302;
	wire w2303;
	wire w2304;
	wire w2305;
	wire w2306;
	wire w2307;
	wire w2308;
	wire w2309;
	wire w2310;
	wire w2311;
	wire w2312;
	wire w2313;
	wire w2314;
	wire w2315;
	wire w2316;
	wire w2317;
	wire w2318;
	wire w2319;
	wire w2320;
	wire w2321;
	wire w2322;
	wire w2323;
	wire w2324;
	wire w2325;
	wire w2326;
	wire w2327;
	wire w2328;
	wire w2329;
	wire w2330;
	wire w2331;
	wire w2332;
	wire w2333;
	wire w2334;
	wire w2335;
	wire w2336;
	wire w2337;
	wire w2338;
	wire w2339;
	wire w2340;
	wire w2341;
	wire w2342;
	wire w2343;
	wire w2344;
	wire w2345;
	wire w2346;
	wire w2347;
	wire w2348;
	wire w2349;
	wire w2350;
	wire w2351;
	wire w2352;
	wire w2353;
	wire w2354;
	wire w2355;
	wire w2356;
	wire w2357;
	wire w2358;
	wire w2359;
	wire w2360;
	wire w2361;
	wire w2362;
	wire w2363;
	wire w2364;
	wire w2365;
	wire w2366;
	wire w2367;
	wire w2368;
	wire w2369;
	wire w2370;
	wire w2371;
	wire w2372;
	wire w2373;
	wire w2374;
	wire w2375;
	wire w2376;
	wire w2377;
	wire w2378;
	wire w2379;
	wire w2380;
	wire w2381;
	wire w2382;
	wire w2383;
	wire w2384;
	wire w2385;
	wire w2386;
	wire w2387;
	wire w2388;
	wire w2389;
	wire w2390;
	wire w2391;
	wire w2392;
	wire w2393;
	wire w2394;
	wire w2395;
	wire w2396;
	wire w2397;
	wire w2398;
	wire w2399;
	wire w2400;
	wire w2401;
	wire w2402;
	wire w2403;
	wire w2404;
	wire w2405;
	wire w2406;
	wire w2407;
	wire w2408;
	wire w2409;
	wire w2410;
	wire w2411;
	wire w2412;
	wire w2413;
	wire w2414;
	wire w2415;
	wire w2416;
	wire w2417;
	wire w2418;
	wire w2419;
	wire w2420;
	wire w2421;
	wire w2422;
	wire w2423;
	wire w2424;
	wire w2425;
	wire w2426;
	wire w2427;
	wire w2428;
	wire w2429;
	wire w2430;
	wire w2431;
	wire w2432;
	wire w2433;
	wire w2434;
	wire w2435;
	wire w2436;
	wire w2437;
	wire w2438;
	wire w2439;
	wire w2440;
	wire w2441;
	wire w2442;
	wire w2443;
	wire w2444;
	wire w2445;
	wire w2446;
	wire w2447;
	wire w2448;
	wire w2449;
	wire w2450;
	wire w2451;
	wire w2452;
	wire w2453;
	wire w2454;
	wire w2455;
	wire w2456;
	wire w2457;
	wire w2458;
	wire w2459;
	wire w2460;
	wire w2461;
	wire w2462;
	wire w2463;
	wire w2464;
	wire w2465;
	wire w2466;
	wire w2467;
	wire w2468;
	wire w2469;
	wire w2470;
	wire w2471;
	wire w2472;
	wire w2473;
	wire w2474;
	wire w2475;
	wire w2476;
	wire w2477;
	wire w2478;
	wire w2479;
	wire w2480;
	wire w2481;
	wire w2482;
	wire w2483;
	wire w2484;
	wire w2485;
	wire w2486;
	wire w2487;
	wire w2488;
	wire w2489;
	wire w2490;
	wire w2491;
	wire w2492;
	wire w2493;
	wire w2494;
	wire w2495;
	wire w2496;
	wire w2497;
	wire w2498;
	wire w2499;
	wire w2500;
	wire w2501;
	wire w2502;
	wire w2503;
	wire w2504;
	wire w2505;
	wire w2506;
	wire w2507;
	wire w2508;
	wire w2509;
	wire w2510;
	wire w2511;
	wire w2512;
	wire w2513;
	wire w2514;
	wire w2515;
	wire w2516;
	wire w2517;
	wire w2518;
	wire w2519;
	wire w2520;
	wire w2521;
	wire w2522;
	wire w2523;
	wire w2524;
	wire w2525;
	wire w2526;
	wire w2527;
	wire w2528;
	wire w2529;
	wire w2530;
	wire w2531;
	wire w2532;
	wire w2533;
	wire w2534;
	wire w2535;
	wire w2536;
	wire w2537;
	wire w2538;
	wire w2539;
	wire w2540;
	wire w2541;
	wire w2542;
	wire w2543;
	wire w2544;
	wire w2545;
	wire w2546;
	wire w2547;
	wire w2548;
	wire w2549;
	wire w2550;
	wire w2551;
	wire w2552;
	wire w2553;
	wire w2554;
	wire w2555;
	wire w2556;
	wire w2557;
	wire w2558;
	wire w2559;
	wire w2560;
	wire w2561;
	wire w2562;
	wire w2563;
	wire w2564;
	wire w2565;
	wire w2566;
	wire w2567;
	wire w2568;
	wire w2569;
	wire w2570;
	wire w2571;
	wire w2572;
	wire w2573;
	wire w2574;
	wire w2575;
	wire w2576;
	wire w2577;
	wire w2578;
	wire w2579;
	wire w2580;
	wire w2581;
	wire w2582;
	wire w2583;
	wire w2584;
	wire w2585;
	wire w2586;
	wire w2587;
	wire w2588;
	wire w2589;
	wire w2590;
	wire w2591;
	wire w2592;
	wire w2593;
	wire w2594;
	wire w2595;
	wire w2596;
	wire w2597;
	wire w2598;
	wire w2599;
	wire w2600;
	wire w2601;
	wire w2602;
	wire w2603;
	wire w2604;
	wire w2605;
	wire w2606;
	wire w2607;
	wire w2608;
	wire w2609;
	wire w2610;
	wire w2611;
	wire w2612;
	wire w2613;
	wire w2614;
	wire w2615;
	wire w2616;
	wire w2617;
	wire w2618;
	wire w2619;
	wire w2620;
	wire w2621;
	wire w2622;
	wire w2623;
	wire w2624;
	wire w2625;
	wire w2626;
	wire w2627;
	wire w2628;
	wire w2629;
	wire w2630;
	wire w2631;
	wire w2632;
	wire w2633;
	wire w2634;
	wire w2635;
	wire w2636;
	wire w2637;
	wire w2638;
	wire w2639;
	wire w2640;
	wire w2641;
	wire w2642;
	wire w2643;
	wire w2644;
	wire w2645;
	wire w2646;
	wire w2647;
	wire w2648;
	wire w2649;
	wire w2650;
	wire w2651;
	wire w2652;
	wire w2653;
	wire w2654;
	wire w2655;
	wire w2656;
	wire w2657;
	wire w2658;
	wire w2659;
	wire w2660;
	wire w2661;
	wire w2662;
	wire w2663;
	wire w2664;
	wire w2665;
	wire w2666;
	wire w2667;
	wire w2668;
	wire w2669;
	wire w2670;
	wire w2671;
	wire w2672;
	wire w2673;
	wire w2674;
	wire w2675;
	wire w2676;
	wire w2677;
	wire w2678;
	wire w2679;
	wire w2680;
	wire w2681;
	wire w2682;
	wire w2683;
	wire w2684;
	wire w2685;
	wire w2686;
	wire w2687;
	wire w2688;
	wire w2689;
	wire w2690;
	wire w2691;
	wire w2692;
	wire w2693;
	wire w2694;
	wire w2695;
	wire w2696;
	wire w2697;
	wire w2698;
	wire w2699;
	wire w2700;
	wire w2701;
	wire w2702;
	wire w2703;
	wire w2704;
	wire w2705;
	wire w2706;
	wire w2707;
	wire w2708;
	wire w2709;
	wire w2710;
	wire w2711;
	wire w2712;
	wire w2713;
	wire w2714;
	wire w2715;
	wire w2716;
	wire w2717;
	wire w2718;
	wire w2719;
	wire w2720;
	wire w2721;
	wire w2722;
	wire w2723;
	wire w2724;
	wire w2725;
	wire w2726;
	wire w2727;
	wire w2728;
	wire w2729;
	wire w2730;
	wire w2731;
	wire w2732;
	wire w2733;
	wire w2734;
	wire w2735;
	wire w2736;
	wire w2737;
	wire w2738;
	wire w2739;
	wire w2740;
	wire w2741;
	wire w2742;
	wire w2743;
	wire w2744;
	wire w2745;
	wire w2746;
	wire w2747;
	wire w2748;
	wire w2749;
	wire w2750;
	wire w2751;
	wire w2752;
	wire w2753;
	wire w2754;
	wire w2755;
	wire w2756;
	wire w2757;
	wire w2758;
	wire w2759;
	wire w2760;
	wire w2761;
	wire w2762;
	wire w2763;
	wire w2764;
	wire w2765;
	wire w2766;
	wire w2767;
	wire w2768;
	wire w2769;
	wire w2770;
	wire w2771;
	wire w2772;
	wire w2773;
	wire w2774;
	wire w2775;
	wire w2776;
	wire w2777;
	wire w2778;
	wire w2779;
	wire w2780;
	wire w2781;
	wire w2782;
	wire w2783;
	wire w2784;
	wire w2785;
	wire w2786;
	wire w2787;
	wire w2788;
	wire w2789;
	wire w2790;
	wire w2791;
	wire w2792;
	wire w2793;
	wire w2794;
	wire w2795;
	wire w2796;
	wire w2797;
	wire w2798;
	wire w2799;
	wire w2800;
	wire w2801;
	wire w2802;
	wire w2803;
	wire w2804;
	wire w2805;
	wire w2806;
	wire w2807;
	wire w2808;
	wire w2809;
	wire w2810;
	wire w2811;
	wire w2812;
	wire w2813;
	wire w2814;
	wire w2815;
	wire w2816;
	wire w2817;
	wire w2818;
	wire w2819;
	wire w2820;
	wire w2821;
	wire w2822;
	wire w2823;
	wire w2824;
	wire w2825;
	wire w2826;
	wire w2827;
	wire w2828;
	wire w2829;
	wire w2830;
	wire w2831;
	wire w2832;
	wire w2833;
	wire w2834;
	wire w2835;
	wire w2836;
	wire w2837;
	wire w2838;
	wire w2839;
	wire w2840;
	wire w2841;
	wire w2842;
	wire w2843;
	wire w2844;
	wire w2845;
	wire w2846;
	wire w2847;
	wire w2848;
	wire w2849;
	wire w2850;
	wire w2851;
	wire w2852;
	wire w2853;
	wire w2854;
	wire w2855;
	wire w2856;
	wire w2857;
	wire w2858;
	wire w2859;
	wire w2860;
	wire w2861;
	wire w2862;
	wire w2863;
	wire w2864;
	wire w2865;
	wire w2866;
	wire w2867;
	wire w2868;
	wire w2869;
	wire w2870;
	wire w2871;
	wire w2872;
	wire w2873;
	wire w2874;
	wire w2875;
	wire w2876;
	wire w2877;
	wire w2878;
	wire w2879;
	wire w2880;
	wire w2881;
	wire w2882;
	wire w2883;
	wire w2884;
	wire w2885;
	wire w2886;
	wire w2887;
	wire w2888;
	wire w2889;
	wire w2890;
	wire w2891;
	wire w2892;
	wire w2893;
	wire w2894;
	wire w2895;
	wire w2896;
	wire w2897;
	wire w2898;
	wire w2899;
	wire w2900;
	wire w2901;
	wire w2902;
	wire w2903;
	wire w2904;
	wire w2905;
	wire w2906;
	wire w2907;
	wire w2908;
	wire w2909;
	wire w2910;
	wire w2911;
	wire w2912;
	wire w2913;
	wire w2914;
	wire w2915;
	wire w2916;
	wire w2917;
	wire w2918;
	wire w2919;
	wire w2920;
	wire w2921;
	wire w2922;
	wire w2923;
	wire w2924;
	wire w2925;
	wire w2926;
	wire w2927;
	wire w2928;
	wire w2929;
	wire w2930;
	wire w2931;
	wire w2932;
	wire w2933;
	wire w2934;
	wire w2935;
	wire w2936;
	wire w2937;
	wire w2938;
	wire w2939;
	wire w2940;
	wire w2941;
	wire w2942;
	wire w2943;
	wire w2944;
	wire w2945;
	wire w2946;
	wire w2947;
	wire w2948;
	wire w2949;
	wire w2950;
	wire w2951;
	wire w2952;
	wire w2953;
	wire w2954;
	wire w2955;
	wire w2956;
	wire w2957;
	wire w2958;
	wire w2959;
	wire w2960;
	wire w2961;
	wire w2962;
	wire w2963;
	wire w2964;
	wire w2965;
	wire w2966;
	wire w2967;
	wire w2968;
	wire w2969;
	wire w2970;
	wire w2971;
	wire w2972;
	wire w2973;
	wire w2974;
	wire w2975;
	wire w2976;
	wire w2977;
	wire w2978;
	wire w2979;
	wire w2980;
	wire w2981;
	wire w2982;
	wire w2983;
	wire w2984;
	wire w2985;
	wire w2986;
	wire w2987;
	wire w2988;
	wire w2989;
	wire w2990;
	wire w2991;
	wire w2992;
	wire w2993;
	wire w2994;
	wire w2995;
	wire w2996;
	wire w2997;
	wire w2998;
	wire w2999;
	wire w3000;
	wire w3001;
	wire w3002;
	wire w3003;
	wire w3004;
	wire w3005;
	wire w3006;
	wire w3007;
	wire w3008;
	wire w3009;
	wire w3010;
	wire w3011;
	wire w3012;
	wire w3013;
	wire w3014;
	wire w3015;
	wire w3016;
	wire w3017;
	wire w3018;
	wire w3019;
	wire w3020;
	wire w3021;
	wire w3022;
	wire w3023;
	wire w3024;
	wire w3025;
	wire w3026;
	wire w3027;
	wire w3028;
	wire w3029;
	wire w3030;
	wire w3031;
	wire w3032;
	wire w3033;
	wire w3034;
	wire w3035;
	wire w3036;
	wire w3037;
	wire w3038;
	wire w3039;
	wire w3040;
	wire w3041;
	wire w3042;
	wire w3043;
	wire w3044;
	wire w3045;
	wire w3046;
	wire w3047;
	wire w3048;
	wire w3049;
	wire w3050;
	wire w3051;
	wire w3052;
	wire w3053;
	wire w3054;
	wire w3055;
	wire w3056;
	wire w3057;
	wire w3058;
	wire w3059;
	wire w3060;
	wire w3061;
	wire w3062;
	wire w3063;
	wire w3064;
	wire w3065;
	wire w3066;
	wire w3067;
	wire w3068;
	wire w3069;
	wire w3070;
	wire w3071;
	wire w3072;
	wire w3073;
	wire w3074;
	wire w3075;
	wire w3076;
	wire w3077;
	wire w3078;
	wire w3079;
	wire w3080;
	wire w3081;
	wire w3082;
	wire w3083;
	wire w3084;
	wire w3085;
	wire w3086;
	wire w3087;
	wire w3088;
	wire w3089;
	wire w3090;
	wire w3091;
	wire w3092;
	wire w3093;
	wire w3094;
	wire w3095;
	wire w3096;
	wire w3097;
	wire w3098;
	wire w3099;
	wire w3100;
	wire w3101;
	wire w3102;
	wire w3103;
	wire w3104;
	wire w3105;
	wire w3106;
	wire w3107;
	wire w3108;
	wire w3109;
	wire w3110;
	wire w3111;
	wire w3112;
	wire w3113;
	wire w3114;
	wire w3115;
	wire w3116;
	wire w3117;
	wire w3118;
	wire w3119;
	wire w3120;
	wire w3121;
	wire w3122;
	wire w3123;
	wire w3124;
	wire w3125;
	wire w3126;
	wire w3127;
	wire w3128;
	wire w3129;
	wire w3130;
	wire w3131;
	wire w3132;
	wire w3133;
	wire w3134;
	wire w3135;
	wire w3136;
	wire w3137;
	wire w3138;
	wire w3139;
	wire w3140;
	wire w3141;
	wire w3142;
	wire w3143;
	wire w3144;
	wire w3145;
	wire w3146;
	wire w3147;
	wire w3148;
	wire w3149;
	wire w3150;
	wire w3151;
	wire w3152;
	wire w3153;
	wire w3154;
	wire w3155;
	wire w3156;
	wire w3157;
	wire w3158;
	wire w3159;
	wire w3160;
	wire w3161;
	wire w3162;
	wire w3163;
	wire w3164;
	wire w3165;
	wire w3166;
	wire w3167;
	wire w3168;
	wire w3169;
	wire w3170;
	wire w3171;
	wire w3172;
	wire w3173;
	wire w3174;
	wire w3175;
	wire w3176;
	wire w3177;
	wire w3178;
	wire w3179;
	wire w3180;
	wire w3181;
	wire w3182;
	wire w3183;
	wire w3184;
	wire w3185;
	wire w3186;
	wire w3187;
	wire w3188;
	wire w3189;
	wire w3190;
	wire w3191;
	wire w3192;
	wire w3193;
	wire w3194;
	wire w3195;
	wire w3196;
	wire w3197;
	wire w3198;
	wire w3199;
	wire w3200;
	wire w3201;
	wire w3202;
	wire w3203;
	wire w3204;
	wire w3205;
	wire w3206;
	wire w3207;
	wire w3208;
	wire w3209;
	wire w3210;
	wire w3211;
	wire w3212;
	wire w3213;
	wire w3214;
	wire w3215;
	wire w3216;
	wire w3217;
	wire w3218;
	wire w3219;
	wire w3220;
	wire w3221;
	wire w3222;
	wire w3223;
	wire w3224;
	wire w3225;
	wire w3226;
	wire w3227;
	wire w3228;
	wire w3229;
	wire w3230;
	wire w3231;
	wire w3232;
	wire w3233;
	wire w3234;
	wire w3235;
	wire w3236;
	wire w3237;
	wire w3238;
	wire w3239;
	wire w3240;
	wire w3241;
	wire w3242;
	wire w3243;
	wire w3244;
	wire w3245;
	wire w3246;
	wire w3247;
	wire w3248;
	wire w3249;
	wire w3250;
	wire w3251;
	wire w3252;
	wire w3253;
	wire w3254;
	wire w3255;
	wire w3256;
	wire w3257;
	wire w3258;
	wire w3259;
	wire w3260;
	wire w3261;
	wire w3262;
	wire w3263;
	wire w3264;
	wire w3265;
	wire w3266;
	wire w3267;
	wire w3268;
	wire w3269;
	wire w3270;
	wire w3271;
	wire w3272;
	wire w3273;
	wire w3274;
	wire w3275;
	wire w3276;
	wire w3277;
	wire w3278;
	wire w3279;
	wire w3280;
	wire w3281;
	wire w3282;
	wire w3283;
	wire w3284;
	wire w3285;
	wire w3286;
	wire w3287;
	wire w3288;
	wire w3289;
	wire w3290;
	wire w3291;
	wire w3292;
	wire w3293;
	wire w3294;
	wire w3295;
	wire w3296;
	wire w3297;
	wire w3298;
	wire w3299;
	wire w3300;
	wire w3301;
	wire w3302;
	wire w3303;
	wire w3304;
	wire w3305;
	wire w3306;
	wire w3307;
	wire w3308;
	wire w3309;
	wire w3310;
	wire w3311;
	wire w3312;
	wire w3313;
	wire w3314;
	wire w3315;
	wire w3316;
	wire w3317;
	wire w3318;
	wire w3319;
	wire w3320;
	wire w3321;
	wire w3322;
	wire w3323;
	wire w3324;
	wire w3325;
	wire w3326;
	wire w3327;
	wire w3328;
	wire w3329;
	wire w3330;
	wire w3331;
	wire w3332;
	wire w3333;
	wire w3334;
	wire w3335;
	wire w3336;
	wire w3337;
	wire w3338;
	wire w3339;
	wire w3340;
	wire w3341;
	wire w3342;
	wire w3343;
	wire w3344;
	wire w3345;
	wire w3346;
	wire w3347;
	wire w3348;
	wire w3349;
	wire w3350;
	wire w3351;
	wire w3352;
	wire w3353;
	wire w3354;
	wire w3355;
	wire w3356;
	wire w3357;
	wire w3358;
	wire w3359;
	wire w3360;
	wire w3361;
	wire w3362;
	wire w3363;
	wire w3364;
	wire w3365;
	wire w3366;
	wire w3367;
	wire w3368;
	wire w3369;
	wire w3370;
	wire w3371;
	wire w3372;
	wire w3373;
	wire w3374;
	wire w3375;
	wire w3376;
	wire w3377;
	wire w3378;
	wire w3379;
	wire w3380;
	wire w3381;
	wire w3382;
	wire w3383;
	wire w3384;
	wire w3385;
	wire w3386;
	wire w3387;
	wire w3388;
	wire w3389;
	wire w3390;
	wire w3391;
	wire w3392;
	wire w3393;
	wire w3394;
	wire w3395;
	wire w3396;
	wire w3397;
	wire w3398;
	wire w3399;
	wire w3400;
	wire w3401;
	wire w3402;
	wire w3403;
	wire w3404;
	wire w3405;
	wire w3406;
	wire w3407;
	wire w3408;
	wire w3409;
	wire w3410;
	wire w3411;
	wire w3412;
	wire w3413;
	wire w3414;
	wire w3415;
	wire w3416;
	wire w3417;
	wire w3418;
	wire w3419;
	wire w3420;
	wire w3421;
	wire w3422;
	wire w3423;
	wire w3424;
	wire w3425;
	wire w3426;
	wire w3427;
	wire w3428;
	wire w3429;
	wire w3430;
	wire w3431;
	wire w3432;
	wire w3433;
	wire w3434;
	wire w3435;
	wire w3436;
	wire w3437;
	wire w3438;
	wire w3439;
	wire w3440;
	wire w3441;
	wire w3442;
	wire w3443;
	wire w3444;
	wire w3445;
	wire w3446;
	wire w3447;
	wire w3448;
	wire w3449;
	wire w3450;
	wire w3451;
	wire w3452;
	wire w3453;
	wire w3454;
	wire w3455;
	wire w3456;
	wire w3457;
	wire w3458;
	wire w3459;
	wire w3460;
	wire w3461;
	wire w3462;
	wire w3463;
	wire w3464;
	wire w3465;
	wire w3466;
	wire w3467;
	wire w3468;
	wire w3469;
	wire w3470;
	wire w3471;
	wire w3472;
	wire w3473;
	wire w3474;
	wire w3475;
	wire w3476;
	wire w3477;
	wire w3478;
	wire w3479;
	wire w3480;
	wire w3481;
	wire w3482;
	wire w3483;
	wire w3484;
	wire w3485;
	wire w3486;
	wire w3487;
	wire w3488;
	wire w3489;
	wire w3490;
	wire w3491;
	wire w3492;
	wire w3493;
	wire w3494;
	wire w3495;
	wire w3496;
	wire w3497;
	wire w3498;
	wire w3499;
	wire w3500;
	wire w3501;
	wire w3502;
	wire w3503;
	wire w3504;
	wire w3505;
	wire w3506;
	wire w3507;
	wire w3508;
	wire w3509;
	wire w3510;
	wire w3511;
	wire w3512;
	wire w3513;
	wire w3514;
	wire w3515;
	wire w3516;
	wire w3517;
	wire w3518;
	wire w3519;
	wire w3520;
	wire w3521;
	wire w3522;
	wire w3523;
	wire w3524;
	wire w3525;
	wire w3526;
	wire w3527;
	wire w3528;
	wire w3529;
	wire w3530;
	wire w3531;
	wire w3532;
	wire w3533;
	wire w3534;
	wire w3535;
	wire w3536;
	wire w3537;
	wire w3538;
	wire w3539;
	wire w3540;
	wire w3541;
	wire w3542;
	wire w3543;
	wire w3544;
	wire w3545;
	wire w3546;
	wire w3547;
	wire w3548;
	wire w3549;
	wire w3550;
	wire w3551;
	wire w3552;
	wire w3553;
	wire w3554;
	wire w3555;
	wire w3556;
	wire w3557;
	wire w3558;
	wire w3559;
	wire w3560;
	wire w3561;
	wire w3562;
	wire w3563;
	wire w3564;
	wire w3565;
	wire w3566;
	wire w3567;
	wire w3568;
	wire w3569;
	wire w3570;
	wire w3571;
	wire w3572;
	wire w3573;
	wire w3574;
	wire w3575;
	wire w3576;
	wire w3577;
	wire w3578;
	wire w3579;
	wire w3580;
	wire w3581;
	wire w3582;
	wire w3583;
	wire w3584;
	wire w3585;
	wire w3586;
	wire w3587;
	wire w3588;
	wire w3589;
	wire w3590;
	wire w3591;
	wire w3592;
	wire w3593;
	wire w3594;
	wire w3595;
	wire w3596;
	wire w3597;
	wire w3598;
	wire w3599;
	wire w3600;
	wire w3601;
	wire w3602;
	wire w3603;
	wire w3604;
	wire w3605;
	wire w3606;
	wire w3607;
	wire w3608;
	wire w3609;
	wire w3610;
	wire w3611;
	wire w3612;
	wire w3613;
	wire w3614;
	wire w3615;
	wire w3616;
	wire w3617;
	wire w3618;
	wire w3619;
	wire w3620;
	wire w3621;
	wire w3622;
	wire w3623;
	wire w3624;
	wire w3625;
	wire w3626;
	wire w3627;
	wire w3628;
	wire w3629;
	wire w3630;
	wire w3631;
	wire w3632;
	wire w3633;
	wire w3634;
	wire w3635;
	wire w3636;
	wire w3637;
	wire w3638;
	wire w3639;
	wire w3640;
	wire w3641;
	wire w3642;
	wire w3643;
	wire w3644;
	wire w3645;
	wire w3646;
	wire w3647;
	wire w3648;
	wire w3649;
	wire w3650;
	wire w3651;
	wire w3652;
	wire w3653;
	wire w3654;
	wire w3655;
	wire w3656;
	wire w3657;
	wire w3658;
	wire w3659;
	wire w3660;
	wire w3661;
	wire w3662;
	wire w3663;
	wire w3664;
	wire w3665;
	wire w3666;
	wire w3667;
	wire w3668;
	wire w3669;
	wire w3670;
	wire w3671;
	wire w3672;
	wire w3673;
	wire w3674;
	wire w3675;
	wire w3676;
	wire w3677;
	wire w3678;
	wire w3679;
	wire w3680;
	wire w3681;
	wire w3682;
	wire w3683;
	wire w3684;
	wire w3685;
	wire w3686;
	wire w3687;
	wire w3688;
	wire w3689;
	wire w3690;
	wire w3691;
	wire w3692;
	wire w3693;
	wire w3694;
	wire w3695;
	wire w3696;
	wire w3697;
	wire w3698;
	wire w3699;
	wire w3700;
	wire w3701;
	wire w3702;
	wire w3703;
	wire w3704;
	wire w3705;
	wire w3706;
	wire w3707;
	wire w3708;
	wire w3709;
	wire w3710;
	wire w3711;
	wire w3712;
	wire w3713;
	wire w3714;
	wire w3715;
	wire w3716;
	wire w3717;
	wire w3718;
	wire w3719;
	wire w3720;
	wire w3721;
	wire w3722;
	wire w3723;
	wire w3724;
	wire w3725;
	wire w3726;
	wire w3727;
	wire w3728;
	wire w3729;
	wire w3730;
	wire w3731;
	wire w3732;
	wire w3733;
	wire w3734;
	wire w3735;
	wire w3736;
	wire w3737;
	wire w3738;
	wire w3739;
	wire w3740;
	wire w3741;
	wire w3742;
	wire w3743;
	wire w3744;
	wire w3745;
	wire w3746;
	wire w3747;
	wire w3748;
	wire w3749;
	wire w3750;
	wire w3751;
	wire w3752;
	wire w3753;
	wire w3754;
	wire w3755;
	wire w3756;
	wire w3757;
	wire w3758;
	wire w3759;
	wire w3760;
	wire w3761;
	wire w3762;
	wire w3763;
	wire w3764;
	wire w3765;
	wire w3766;
	wire w3767;
	wire w3768;
	wire w3769;
	wire w3770;
	wire w3771;
	wire w3772;
	wire w3773;
	wire w3774;
	wire w3775;
	wire w3776;
	wire w3777;
	wire w3778;
	wire w3779;
	wire w3780;
	wire w3781;
	wire w3782;
	wire w3783;
	wire w3784;
	wire w3785;
	wire w3786;
	wire w3787;
	wire w3788;
	wire w3789;
	wire w3790;
	wire w3791;
	wire w3792;
	wire w3793;
	wire w3794;
	wire w3795;
	wire w3796;
	wire w3797;
	wire w3798;
	wire w3799;
	wire w3800;
	wire w3801;
	wire w3802;
	wire w3803;
	wire w3804;
	wire w3805;
	wire w3806;
	wire w3807;
	wire w3808;
	wire w3809;
	wire w3810;
	wire w3811;
	wire w3812;
	wire w3813;
	wire w3814;
	wire w3815;
	wire w3816;
	wire w3817;
	wire w3818;
	wire w3819;
	wire w3820;
	wire w3821;
	wire w3822;
	wire w3823;
	wire w3824;
	wire w3825;
	wire w3826;
	wire w3827;
	wire w3828;
	wire w3829;
	wire w3830;
	wire w3831;
	wire w3832;
	wire w3833;
	wire w3834;
	wire w3835;
	wire w3836;
	wire w3837;
	wire w3838;
	wire w3839;
	wire w3840;
	wire w3841;
	wire w3842;
	wire w3843;
	wire w3844;
	wire w3845;
	wire w3846;
	wire w3847;
	wire w3848;
	wire w3849;
	wire w3850;
	wire w3851;
	wire w3852;
	wire w3853;
	wire w3854;
	wire w3855;
	wire w3856;
	wire w3857;
	wire w3858;
	wire w3859;
	wire w3860;
	wire w3861;
	wire w3862;
	wire w3863;
	wire w3864;
	wire w3865;
	wire w3866;
	wire w3867;
	wire w3868;
	wire w3869;
	wire w3870;
	wire w3871;
	wire w3872;
	wire w3873;
	wire w3874;
	wire w3875;
	wire w3876;
	wire w3877;
	wire w3878;
	wire w3879;
	wire w3880;
	wire w3881;
	wire w3882;
	wire w3883;
	wire w3884;
	wire w3885;
	wire w3886;
	wire w3887;
	wire w3888;
	wire w3889;
	wire w3890;
	wire w3891;
	wire w3892;
	wire w3893;
	wire w3894;
	wire w3895;
	wire w3896;
	wire w3897;
	wire w3898;
	wire w3899;
	wire w3900;
	wire w3901;
	wire w3902;
	wire w3903;
	wire w3904;
	wire w3905;
	wire w3906;
	wire w3907;
	wire w3908;
	wire w3909;
	wire w3910;
	wire w3911;
	wire w3912;
	wire w3913;
	wire w3914;
	wire w3915;
	wire w3916;
	wire w3917;
	wire w3918;
	wire w3919;
	wire w3920;
	wire w3921;
	wire w3922;
	wire w3923;
	wire w3924;
	wire w3925;
	wire w3926;
	wire w3927;
	wire w3928;
	wire w3929;
	wire w3930;
	wire w3931;
	wire w3932;
	wire w3933;
	wire w3934;
	wire w3935;
	wire w3936;
	wire w3937;
	wire w3938;
	wire w3939;
	wire w3940;
	wire w3941;
	wire w3942;
	wire w3943;
	wire w3944;
	wire w3945;
	wire w3946;
	wire w3947;
	wire w3948;
	wire w3949;
	wire w3950;
	wire w3951;
	wire w3952;
	wire w3953;
	wire w3954;
	wire w3955;
	wire w3956;
	wire w3957;
	wire w3958;
	wire w3959;
	wire w3960;
	wire w3961;
	wire w3962;
	wire w3963;
	wire w3964;
	wire w3965;
	wire w3966;
	wire w3967;
	wire w3968;
	wire w3969;
	wire w3970;
	wire w3971;
	wire w3972;
	wire w3973;
	wire w3974;
	wire w3975;
	wire w3976;
	wire w3977;
	wire w3978;
	wire w3979;
	wire w3980;
	wire w3981;
	wire w3982;
	wire w3983;
	wire w3984;
	wire w3985;
	wire w3986;
	wire w3987;
	wire w3988;
	wire w3989;
	wire w3990;
	wire w3991;
	wire w3992;
	wire w3993;
	wire w3994;
	wire w3995;
	wire w3996;
	wire w3997;
	wire w3998;
	wire w3999;
	wire w4000;
	wire w4001;
	wire w4002;
	wire w4003;
	wire w4004;
	wire w4005;
	wire w4006;
	wire w4007;
	wire w4008;
	wire w4009;
	wire w4010;
	wire w4011;
	wire w4012;
	wire w4013;
	wire w4014;
	wire w4015;
	wire w4016;
	wire w4017;
	wire w4018;
	wire w4019;
	wire w4020;
	wire w4021;
	wire w4022;
	wire w4023;
	wire w4024;
	wire w4025;
	wire w4026;
	wire w4027;
	wire w4028;
	wire w4029;
	wire w4030;
	wire w4031;
	wire w4032;
	wire w4033;
	wire w4034;
	wire w4035;
	wire w4036;
	wire w4037;
	wire w4038;
	wire w4039;
	wire w4040;
	wire w4041;
	wire w4042;
	wire w4043;
	wire w4044;
	wire w4045;
	wire w4046;
	wire w4047;
	wire w4048;
	wire w4049;
	wire w4050;
	wire w4051;
	wire w4052;
	wire w4053;
	wire w4054;
	wire w4055;
	wire w4056;
	wire w4057;
	wire w4058;
	wire w4059;
	wire w4060;
	wire w4061;
	wire w4062;
	wire w4063;
	wire w4064;
	wire w4065;
	wire w4066;
	wire w4067;
	wire w4068;
	wire w4069;
	wire w4070;
	wire w4071;
	wire w4072;
	wire w4073;
	wire w4074;
	wire w4075;
	wire w4076;
	wire w4077;
	wire w4078;
	wire w4079;
	wire w4080;
	wire w4081;
	wire w4082;
	wire w4083;
	wire w4084;
	wire w4085;
	wire w4086;
	wire w4087;
	wire w4088;
	wire w4089;
	wire w4090;
	wire w4091;
	wire w4092;
	wire w4093;
	wire w4094;
	wire w4095;
	wire w4096;
	wire w4097;
	wire w4098;
	wire w4099;
	wire w4100;
	wire w4101;
	wire w4102;
	wire w4103;
	wire w4104;
	wire w4105;
	wire w4106;
	wire w4107;
	wire w4108;
	wire w4109;
	wire w4110;
	wire w4111;
	wire w4112;
	wire w4113;
	wire w4114;
	wire w4115;
	wire w4116;
	wire w4117;
	wire w4118;
	wire w4119;
	wire w4120;
	wire w4121;
	wire w4122;
	wire w4123;
	wire w4124;
	wire w4125;
	wire w4126;
	wire w4127;
	wire w4128;
	wire w4129;
	wire w4130;
	wire w4131;
	wire w4132;
	wire w4133;
	wire w4134;
	wire w4135;
	wire w4136;
	wire w4137;
	wire w4138;
	wire w4139;
	wire w4140;
	wire w4141;
	wire w4142;
	wire w4143;
	wire w4144;
	wire w4145;
	wire w4146;
	wire w4147;
	wire w4148;
	wire w4149;
	wire w4150;
	wire w4151;
	wire w4152;
	wire w4153;
	wire w4154;
	wire w4155;
	wire w4156;
	wire w4157;
	wire w4158;
	wire w4159;
	wire w4160;
	wire w4161;
	wire w4162;
	wire w4163;
	wire w4164;
	wire w4165;
	wire w4166;
	wire w4167;
	wire w4168;
	wire w4169;
	wire w4170;
	wire w4171;
	wire w4172;
	wire w4173;
	wire w4174;
	wire w4175;
	wire w4176;
	wire w4177;
	wire w4178;
	wire w4179;
	wire w4180;
	wire w4181;
	wire w4182;
	wire w4183;
	wire w4184;
	wire w4185;
	wire w4186;
	wire w4187;
	wire w4188;
	wire w4189;
	wire w4190;
	wire w4191;
	wire w4192;
	wire w4193;
	wire w4194;
	wire w4195;
	wire w4196;
	wire w4197;
	wire w4198;
	wire w4199;
	wire w4200;
	wire w4201;
	wire w4202;
	wire w4203;
	wire w4204;
	wire w4205;
	wire w4206;
	wire w4207;
	wire w4208;
	wire w4209;
	wire w4210;
	wire w4211;
	wire w4212;
	wire w4213;
	wire w4214;
	wire w4215;
	wire w4216;
	wire w4217;
	wire w4218;
	wire w4219;
	wire w4220;
	wire w4221;
	wire w4222;
	wire w4223;
	wire w4224;
	wire w4225;
	wire w4226;
	wire w4227;
	wire w4228;
	wire w4229;
	wire w4230;
	wire w4231;
	wire w4232;
	wire w4233;
	wire w4234;
	wire w4235;
	wire w4236;
	wire w4237;
	wire w4238;
	wire w4239;
	wire w4240;
	wire w4241;
	wire w4242;
	wire w4243;
	wire w4244;
	wire w4245;
	wire w4246;
	wire w4247;
	wire w4248;
	wire w4249;
	wire w4250;
	wire w4251;
	wire w4252;
	wire w4253;
	wire w4254;
	wire w4255;
	wire w4256;
	wire w4257;
	wire w4258;
	wire w4259;
	wire w4260;
	wire w4261;
	wire w4262;
	wire w4263;
	wire w4264;
	wire w4265;
	wire w4266;
	wire w4267;
	wire w4268;
	wire w4269;
	wire w4270;
	wire w4271;
	wire w4272;
	wire w4273;
	wire w4274;
	wire w4275;
	wire w4276;
	wire w4277;
	wire w4278;
	wire w4279;
	wire w4280;
	wire w4281;
	wire w4282;
	wire w4283;
	wire w4284;
	wire w4285;
	wire w4286;
	wire w4287;
	wire w4288;
	wire w4289;
	wire w4290;
	wire w4291;
	wire w4292;
	wire w4293;
	wire w4294;
	wire w4295;
	wire w4296;
	wire w4297;
	wire w4298;
	wire w4299;
	wire w4300;
	wire w4301;
	wire w4302;
	wire w4303;
	wire w4304;
	wire w4305;
	wire w4306;
	wire w4307;
	wire w4308;
	wire w4309;
	wire w4310;
	wire w4311;
	wire w4312;
	wire w4313;
	wire w4314;
	wire w4315;
	wire w4316;
	wire w4317;
	wire w4318;
	wire w4319;
	wire w4320;
	wire w4321;
	wire w4322;
	wire w4323;
	wire w4324;
	wire w4325;
	wire w4326;
	wire w4327;
	wire w4328;
	wire w4329;
	wire w4330;
	wire w4331;
	wire w4332;
	wire w4333;
	wire w4334;
	wire w4335;
	wire w4336;
	wire w4337;
	wire w4338;
	wire w4339;
	wire w4340;
	wire w4341;
	wire w4342;
	wire w4343;
	wire w4344;
	wire w4345;
	wire w4346;
	wire w4347;
	wire w4348;
	wire w4349;
	wire w4350;
	wire w4351;
	wire w4352;
	wire w4353;
	wire w4354;
	wire w4355;
	wire w4356;
	wire w4357;
	wire w4358;
	wire w4359;
	wire w4360;
	wire w4361;
	wire w4362;
	wire w4363;
	wire w4364;
	wire w4365;
	wire w4366;
	wire w4367;
	wire w4368;
	wire w4369;
	wire w4370;
	wire w4371;
	wire w4372;
	wire w4373;
	wire w4374;
	wire w4375;
	wire w4376;
	wire w4377;
	wire w4378;
	wire w4379;
	wire w4380;
	wire w4381;
	wire w4382;
	wire w4383;
	wire w4384;
	wire w4385;
	wire w4386;
	wire w4387;
	wire w4388;
	wire w4389;
	wire w4390;
	wire w4391;
	wire w4392;
	wire w4393;
	wire w4394;
	wire w4395;
	wire w4396;
	wire w4397;
	wire w4398;
	wire w4399;
	wire w4400;
	wire w4401;
	wire w4402;
	wire w4403;
	wire w4404;
	wire w4405;
	wire w4406;
	wire w4407;
	wire w4408;
	wire w4409;
	wire w4410;
	wire w4411;
	wire w4412;
	wire w4413;
	wire w4414;
	wire w4415;
	wire w4416;
	wire w4417;
	wire w4418;
	wire w4419;
	wire w4420;
	wire w4421;
	wire w4422;
	wire w4423;
	wire w4424;
	wire w4425;
	wire w4426;
	wire w4427;
	wire w4428;
	wire w4429;
	wire w4430;
	wire w4431;
	wire w4432;
	wire w4433;
	wire w4434;
	wire w4435;
	wire w4436;
	wire w4437;
	wire w4438;
	wire w4439;
	wire w4440;
	wire w4441;
	wire w4442;
	wire w4443;
	wire w4444;
	wire w4445;
	wire w4446;
	wire w4447;
	wire w4448;
	wire w4449;
	wire w4450;
	wire w4451;
	wire w4452;
	wire w4453;
	wire w4454;
	wire w4455;
	wire w4456;
	wire w4457;
	wire w4458;
	wire w4459;
	wire w4460;
	wire w4461;
	wire w4462;
	wire w4463;
	wire w4464;
	wire w4465;
	wire w4466;
	wire w4467;
	wire w4468;
	wire w4469;
	wire w4470;
	wire w4471;
	wire w4472;
	wire w4473;
	wire w4474;
	wire w4475;
	wire w4476;
	wire w4477;
	wire w4478;
	wire w4479;
	wire w4480;

	assign w1074 = D0_i;
	assign D0_o = w1156;
	assign D0_d = w1076;
	assign w1311 = D1_i;
	assign D1_o = w1155;
	assign D1_d = w1076;
	assign w1312 = D2_i;
	assign D2_o = w1157;
	assign D2_d = w1076;
	assign w1317 = D3_i;
	assign D3_o = w1158;
	assign D3_d = w1076;
	assign w1075 = D4_i;
	assign D4_o = w1159;
	assign D4_d = w1076;
	assign w1077 = D5_i;
	assign D5_o = w1160;
	assign D5_d = w1076;
	assign w1313 = D6_i;
	assign D6_o = w1151;
	assign D6_d = w1076;
	assign w1314 = D7_i;
	assign D7_o = w1078;
	assign D7_d = w1076;
	assign w1153 = TEST_i;
	assign TEST_o = w847;
	assign TEST_d = w114;
	assign w1315 = n_IC;
	assign n_IRQ = w1079;
	assign w1152 = n_CS;
	assign w1316 = n_WR;
	assign w1154 = n_RD;
	assign w1090 = A0;
	assign w1318 = A1;
	assign w821 = M;
	assign MOR_sel = w862;
	assign MOL_sel = w861;
	assign DAC_8 = w853;
	assign DAC_7 = w854;
	assign DAC_6 = w855;
	assign DAC_5 = w857;
	assign DAC_4 = w858;
	assign DAC_3 = w70;
	assign DAC_2 = w860;
	assign DAC_1 = w859;
	assign DAC_0 = w856;

	// Instances

	ym3438_NOR g_1 (.Z(w1306), .A(w4095), .B(w4096) );
	ym3438_NOR g_3 (.A(w821), .Z(w1338), .B(w1307) );
	ym3438_CNT_BIT g_4 (.CI(w845), .Q(w1339), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833), .RES(w827), .CO(w1308) );
	ym3438_CNT_BIT g_5 (.CI(w1308), .Q(w844), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833), .RES(w827) );
	ym3438_OR g_6 (.A(w831), .Z(w1340), .B(w827) );
	ym3438_SR_BIT g_8 (.Q(w1342), .D(w1343), .C1(w1310), .C2(w1309), .nC1(w830), .nC2(w1341) );
	ym3438_NOT g_9 (.A(w214), .nZ(w835) );
	ym3438_SDELAY12 g_10 (.A(w835), .C1(w1310), .C2(w1309), .nC1(w830), .nC2(w1341), .C3(w1310), .C4(w1309), .C5(w1310), .C6(w1309), .C7(w1310), .C8(w1309), .C9(w1310), .C10(w1309), .C11(w1310), .C12(w1309), .C13(w1310), .C14(w1309), .C15(w1310), .C16(w1309), .C17(w1310), .C18(w1309), .C19(w1310), .C20(w1309), .C21(w1310), .C22(w1309), .C23(w1310), .C24(w1309), .nC3(w830), .nC4(w1341), .nC5(w830), .nC6(w1341), .nC7(w830), .nC8(w1341), .nC9(w830), .nC10(w1341), .nC11(w830), .nC12(w1341), .nC13(w830), .nC14(w1341), .nC15(w830), .nC16(w1341), .nC17(w830), .nC18(w1341), .nC19(w830), .nC20(w1341), .nC21(w830), .nC22(w1341), .nC23(w830), .nC24(w1341), .Q(w1345) );
	ym3438_SR_BIT g_11 (.Q(w827), .D(w1342), .C1(w1310), .C2(w1309), .nC1(w830), .nC2(w1341) );
	ym3438_SR_BIT g_12 (.Q(w1344), .D(w826), .C1(w1310), .C2(w1309), .nC1(w830), .nC2(w1341) );
	ym3438_SR_BIT g_13 (.Q(w1343), .D(w1344), .C1(w1310), .C2(w1309), .nC1(w830), .nC2(w1341) );
	ym3438_NOT g_14 (.A(w1345), .nZ(w1346) );
	ym3438_AND g_15 (.A(w835), .Z(w826), .B(w1346) );
	ym3438_NOR g_16 (.A(w836), .Z(w1347), .B(w826) );
	ym3438_SR_BIT g_17 (.Q(w825), .D(w1347), .C1(w1310), .C2(w1309), .nC1(w830), .nC2(w1341) );
	ym3438_SR_BIT g_18 (.Q(w843), .D(w825), .C1(w1310), .C2(w1309), .nC1(w830), .nC2(w1341) );
	ym3438_SR_BIT g_19 (.Q(w824), .D(w843), .C1(w1310), .C2(w1309), .nC1(w830), .nC2(w1341) );
	ym3438_OR5 g_20 (.A(w825), .Z(w836), .B(w843), .C(w824), .D(w837), .E(w842) );
	ym3438_SR_BIT g_21 (.Q(w837), .D(w824), .C1(w1310), .C2(w1309), .nC1(w830), .nC2(w1341) );
	ym3438_SR_BIT g_22 (.Q(w842), .D(w837), .C1(w1310), .C2(w1309), .nC1(w830), .nC2(w1341) );
	ym3438_SR_BIT g_23 (.Q(w841), .D(w842), .C1(w1310), .C2(w1309), .nC1(w830), .nC2(w1341) );
	ym3438_OR g_24 (.A(w837), .Z(w823), .B(w824) );
	ym3438_OR g_25 (.A(w841), .Z(w838), .B(w825) );
	ym3438_SR_BIT g_26 (.Q(w822), .D(w823), .C1(w1310), .C2(w1309), .nC1(w830), .nC2(w1341) );
	ym3438_SR_BIT g_27 (.Q(w839), .D(w838), .C1(w1310), .C2(w1309), .nC1(w830), .nC2(w1341) );
	ym3438_NOT g_28 (.A(w828), .nZ(w56) );
	ym3438_NOT g_29 (.A(w216), .nZ(w828) );
	ym3438_COMP_WE_STRONG g_30 (.A(w822), .Z(w216), .nZ(w217) );
	ym3438_NOT g_31 (.A(w217), .nZ(w832) );
	ym3438_NOT g_32 (.A(w832), .nZ(w833) );
	ym3438_NOT g_33 (.A(w829), .nZ(w57) );
	ym3438_NOT g_34 (.A(w213), .nZ(w829) );
	ym3438_COMP_WE_STRONG g_35 (.A(w839), .Z(w213), .nZ(w212) );
	ym3438_NOT g_36 (.A(w840), .nZ(w834) );
	ym3438_NOT g_37 (.A(w212), .nZ(w840) );
	ym3438_NOT g_38 (.nZ(w4095), .A(w821) );
	ym3438_BUF2 g_39 (.A(w1338), .Z(w4096) );
	ym3438_COMP_STR g_41 (.A(w1339), .Z(w1350), .nZ(w879) );
	ym3438_CNT_BIT g_42 (.CI(w1369), .Q(w831), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833), .RES(w1340) );
	ym3438_CNT_BIT g_43 (.CI(1'b1), .Q(w880), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833), .RES(w1340), .CO(w1369) );
	ym3438_COMP_STR g_44 (.A(w844), .Z(w1352), .nZ(w1348) );
	ym3438_AND5 g_45 (.A(w1355), .B(w1354), .C(w1353), .D(w879), .E(w1348) );
	ym3438_AND5 g_46 (.A(w1355), .B(w1354), .C(w1358), .D(w879), .E(w1348) );
	ym3438_AND5 g_47 (.A(w1356), .Z(w1359), .B(w1354), .C(w1353), .D(w879), .E(w1352) );
	ym3438_AND5 g_48 (.A(w1355), .Z(w1357), .B(w1365), .C(w1353), .D(w879), .E(w1352) );
	ym3438_AND5 g_49 (.A(w1356), .Z(w1360), .B(w1365), .C(w1353), .D(w879), .E(w1352) );
	ym3438_AND5 g_50 (.A(w1356), .Z(w1361), .B(w1354), .C(w1358), .D(w879), .E(w1352) );
	ym3438_AND5 g_51 (.A(w1355), .Z(w1362), .B(w1365), .C(w1358), .D(w879), .E(w1352) );
	ym3438_AND5 g_52 (.A(w1356), .Z(w1363), .B(w1365), .C(w1358), .D(w879), .E(w1352) );
	ym3438_AND5 g_53 (.A(w1356), .Z(w1364), .B(w1354), .C(w1353), .D(w1350), .E(w1348) );
	ym3438_AND5 g_54 (.A(w1355), .Z(w846), .B(w1365), .C(w1353), .D(w1350), .E(w1348) );
	ym3438_AND5 g_55 (.A(w1356), .Z(w4111), .B(w1365), .C(w1353), .D(w1350), .E(w1348) );
	ym3438_AND5 g_56 (.A(w1356), .Z(w881), .B(w1354), .C(w1358), .D(w1350), .E(w1348) );
	ym3438_AND5 g_57 (.A(w1355), .Z(w1366), .B(w1365), .C(w1358), .D(w1350), .E(w1348) );
	ym3438_AND5 g_58 (.A(w1356), .Z(w882), .B(w1365), .C(w1358), .D(w1350), .E(w1348) );
	ym3438_AND5 g_59 (.A(w1356), .Z(w883), .B(w1354), .C(w1353), .D(w879), .E(w1348) );
	ym3438_AND5 g_60 (.A(w1355), .Z(w875), .B(w1365), .C(w1353), .D(w879), .E(w1348) );
	ym3438_AND5 g_61 (.A(w1356), .Z(w1302), .B(w1365), .C(w1353), .D(w879), .E(w1348) );
	ym3438_AND5 g_62 (.A(w1356), .Z(w884), .B(w1354), .C(w1358), .D(w879), .E(w1348) );
	ym3438_AND5 g_63 (.A(w1355), .Z(w1301), .B(w1365), .C(w1358), .D(w879), .E(w1348) );
	ym3438_AND5 g_64 (.A(w1356), .Z(w874), .B(w1365), .C(w1358), .D(w879), .E(w1348) );
	ym3438_EDGE_DET g_65 (.C1(w57), .D(w884), .nC1(w834), .Q(w1367) );
	ym3438_COMP_STR g_66 (.A(w1367), .Z(w1046) );
	ym3438_COMP_STR g_67 (.A(w874), .Z(w261) );
	ym3438_COMP_STR g_68 (.A(w1301), .Z(w1175) );
	ym3438_COMP_STR g_69 (.A(w884), .Z(w726) );
	ym3438_NOT g_70 (.A(w4109), .nZ(w1381) );
	ym3438_NOR4 g_71 (.A(w1366), .Z(w4109), .B(w875), .C(w883), .D(w882) );
	ym3438_OR6 g_72 (.A(w1301), .Z(w1380), .B(w884), .C(w874), .D(w1302), .E(w875), .F(w883) );
	ym3438_NOR4 g_73 (.A(w884), .Z(w1379), .B(w881), .C(w1361), .D(w1372) );
	ym3438_NOT g_74 (.A(w1379), .nZ(w601) );
	ym3438_NOT g_75 (.A(w1378), .nZ(w1167) );
	ym3438_NOR6 g_76 (.A(w874), .Z(w1378), .B(w875), .C(w881), .D(w1363), .E(w1357), .F(w1372) );
	ym3438_NOT g_77 (.A(w1377), .nZ(w847) );
	ym3438_NOT g_78 (.A(w878), .nZ(w1377) );
	ym3438_NOT g_79 (.A(w1376), .nZ(w848) );
	ym3438_NOR6 g_80 (.A(w882), .Z(w1376), .B(w1366), .C(w881), .D(w4111), .E(w846), .F(w1364) );
	ym3438_NOR6 g_81 (.A(w1361), .Z(w4110), .B(w1362), .C(w1363), .D(w1360), .E(w1357), .F(w1359) );
	ym3438_OR6 g_82 (.A(w1361), .Z(w1375), .B(w1362), .C(w1363), .D(w1360), .E(w1357), .F(w1359) );
	ym3438_AND5 g_83 (.A(w1356), .Z(w1371), .B(w1365), .C(w1352), .D(w1350), .E(w1358) );
	ym3438_AND5 g_84 (.A(w1355), .Z(w1373), .B(w1365), .C(w1352), .D(w1358), .E(w1350) );
	ym3438_AND5 g_85 (.A(w1356), .Z(w1372), .B(w1354), .C(w1352), .D(w1358), .E(w1350) );
	ym3438_AND5 g_86 (.A(w1356), .Z(w876), .B(w1365), .C(w1352), .D(w1350), .E(w1353) );
	ym3438_AND5 g_87 (.A(w1355), .Z(w877), .B(w1365), .C(w1352), .D(w1353), .E(w1350) );
	ym3438_AND5 g_88 (.A(w1356), .Z(w878), .B(w1354), .C(w1352), .D(w1353), .E(w1350) );
	ym3438_OR6 g_89 (.A(w1373), .Z(w1374), .B(w1372), .C(w1371), .D(w876), .E(w877), .F(w878) );
	ym3438_NOR6 g_90 (.A(w1371), .Z(w1370), .B(w1372), .C(w1373), .D(w876), .E(w877), .F(w878) );
	ym3438_AND5 g_91 (.A(w1355), .B(w1354), .C(w1358), .D(w1350), .E(w1348) );
	ym3438_AND5 g_92 (.A(w1355), .B(w1354), .C(w1353), .D(w1350), .E(w1348) );
	ym3438_AND5 g_93 (.A(w1355), .B(w1354), .C(w1358), .D(w1352), .E(w879) );
	ym3438_AND5 g_94 (.A(w1355), .B(w1354), .C(w1353), .D(w1352), .E(w879) );
	ym3438_AND5 g_95 (.A(w1355), .B(w1354), .C(w1368), .D(w1358), .E(w1352) );
	ym3438_AND5 g_96 (.A(w1355), .B(w1354), .C(w1353), .D(w1350), .E(w1352) );
	ym3438_COMP_STR g_97 (.A(w880), .Z(w1355), .nZ(w1356) );
	ym3438_COMP_STR g_98 (.A(w831), .Z(w1354), .nZ(w1365) );
	ym3438_COMP_STR g_99 (.A(w1349), .Z(w1353), .nZ(w1358) );
	ym3438_EDGE_DET g_100 (.C1(w57), .D(w1167), .nC1(w834), .Q(w4025) );
	ym3438_NOR g_101 (.A(w4025), .Z(w1391), .B(w128) );
	ym3438_NOR g_102 (.A(w1166), .Z(w1390), .B(w128) );
	ym3438_COMP_STR g_103 (.A(w4108), .Z(w72), .nZ(w73) );
	ym3438_AOI21 g_104 (.A1(w1381), .Z(w4108), .B(w128), .A2(w864) );
	ym3438_NOR g_105 (.A(w848), .Z(w849), .B(w128) );
	ym3438_OR g_106 (.A(w849), .Z(w1389), .B(w128) );
	ym3438_NOT g_107 (.A(w1389), .nZ(w1388) );
	ym3438_COMP_STR g_108 (.A(w849), .Z(w86), .nZ(w87) );
	ym3438_NOT g_109 (.A(w4027), .nZ(w95) );
	ym3438_NAND g_110 (.A(w850), .Z(w4027), .B(w4026) );
	ym3438_NOT g_111 (.A(w128), .nZ(w4026) );
	ym3438_NOT g_112 (.A(w1387), .nZ(w850) );
	ym3438_AOI2222 g_113 (.A1(1'b1), .Z(w1387), .B1(w48), .A2(w1380), .B2(w1374), .C1(w47), .C2(w1375), .D1(w46), .D2(w848) );
	ym3438_NOT g_114 (.A(w4107), .nZ(w436) );
	ym3438_NOR3 g_115 (.A(w863), .Z(w4107), .B(w1374), .C(w4113) );
	ym3438_AND g_116 (.A(w1375), .Z(w4113), .B(w49) );
	ym3438_AND g_117 (.A(w50), .Z(w863), .B(w1380) );
	ym3438_NOT g_118 (.A(w4106), .nZ(w1166) );
	ym3438_AND g_119 (.A(w1370), .Z(w4106), .B(w4110) );
	ym3438_NAND g_120 (.A(w1375), .Z(w4105), .B(w41) );
	ym3438_AOI22 g_121 (.A1(w51), .Z(w4104), .B1(w1375), .A2(w848), .B2(w1382) );
	ym3438_NOT g_122 (.A(w4105), .nZ(w446) );
	ym3438_NOT g_123 (.A(w4104), .nZ(w447) );
	ym3438_COMP_STR g_124 (.A(w1374), .Z(w357) );
	ym3438_NOT g_125 (.A(w4103), .nZ(w414) );
	ym3438_AOI22 g_126 (.A1(w1375), .Z(w4103), .B1(w1380), .A2(w42), .B2(w852) );
	ym3438_NOT g_127 (.A(w4102), .nZ(w390) );
	ym3438_SR_BIT g_128 (.Q(w4102), .D(w1374), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_NOR g_129 (.A(w871), .Z(w4112), .B(w868) );
	ym3438_NAND g_130 (.A(w4112), .Z(w851), .B(w870) );
	ym3438_NOT g_131 (.A(w870), .nZ(w1385) );
	ym3438_AND3 g_132 (.A(w1385), .Z(w869), .B(w871), .C(w868) );
	ym3438_COMP_STR g_133 (.A(w851), .Z(w1383), .nZ(w1384) );
	ym3438_OR3 g_134 (.A(w39), .Z(w852), .B(w41), .C(w37) );
	ym3438_OR4 g_135 (.A(w37), .Z(w1382), .B(w42), .C(w39), .D(w43) );
	ym3438_OR5 g_136 (.A(w45), .Z(w51), .B(w44), .C(w43), .D(w42), .E(w37) );
	ym3438_OR4 g_137 (.A(w45), .Z(w48), .B(w43), .C(w44), .D(w46) );
	ym3438_OR g_138 (.A(w41), .Z(w49), .B(w44) );
	ym3438_OR g_139 (.A(w39), .Z(w50), .B(w44) );
	ym3438_COMP_WE g_140 (.A(w1171), .Z(w38), .nZ(w35) );
	ym3438_COMP_WE g_141 (.A(w1168), .Z(w40), .nZ(w36) );
	ym3438_COMP_WE g_142 (.A(w33), .Z(w34), .nZ(w32) );
	ym3438_AND3 g_143 (.A(w32), .Z(w37), .B(w36), .C(w35) );
	ym3438_AND3 g_144 (.A(w32), .Z(w39), .B(w36), .C(w38) );
	ym3438_AND3 g_145 (.A(w32), .Z(w41), .B(w40), .C(w35) );
	ym3438_AND3 g_146 (.A(w32), .Z(w42), .B(w40), .C(w38) );
	ym3438_AND3 g_147 (.A(w34), .Z(w43), .B(w36), .C(w35) );
	ym3438_AND3 g_148 (.A(w34), .Z(w44), .B(w36), .C(w38) );
	ym3438_AND3 g_149 (.A(w34), .Z(w45), .B(w40), .C(w35) );
	ym3438_AND3 g_150 (.A(w34), .Z(w46), .B(w40), .C(w38) );
	ym3438_OR3 g_151 (.A(w44), .Z(w47), .B(w45), .C(w46) );
	ym3438_COMP_STR g_152 (.A(w1391), .Z(w1393), .nZ(w1394) );
	ym3438_COMP_STR g_153 (.A(w1390), .Z(w78), .nZ(w79) );
	ym3438_AND g_154 (.A(w95), .Z(w1417), .B(w461) );
	ym3438_FA g_155 (.CO(w1416), .S(w1414), .CI(w128), .A(w1417), .B(w887) );
	ym3438_AOI21 g_156 (.A1(w1414), .Z(w1415), .B(w1384), .A2(w93) );
	ym3438_SDELAY6 g_157 (.A(w1415), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833), .C3(w57), .C4(w56), .C5(w57), .C6(w56), .C7(w57), .C8(w56), .C9(w57), .C10(w56), .C11(w57), .C12(w56), .nC3(w834), .nC4(w833), .nC5(w834), .nC6(w833), .nC7(w834), .nC8(w833), .nC9(w834), .nC10(w833), .nC11(w834), .nC12(w833), .Q(w1413) );
	ym3438_NOR g_158 (.A(w1413), .Z(w887), .B(w1388) );
	ym3438_NOT g_159 (.A(w1413), .nZ(w1412) );
	ym3438_AON22 g_160 (.A1(w86), .Z(w1410), .B2(w1412), .A2(w888), .B1(w87) );
	ym3438_SR_BIT g_161 (.Q(w1409), .D(w1410), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_162 (.Q(w1408), .D(w1409), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_163 (.Q(w1407), .D(w1408), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_164 (.Q(w1411), .D(w1407), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_165 (.Q(w1406), .D(w1411), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_166 (.Q(w888), .D(w1406), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SLATCH g_167 (.Q(w872), .nQ(w1405), .D(w4116), .nC(w1393), .C(w1394) );
	ym3438_AON22 g_168 (.A1(w1406), .Z(w4116), .B2(w888), .A2(w78), .B1(w79) );
	ym3438_AOI22 g_169 (.A1(w872), .Z(w1403), .B2(w873), .A2(w72), .B1(w73) );
	ym3438_NOT g_170 (.A(w1403), .nZ(w856) );
	ym3438_NOT g_171 (.A(w1405), .nZ(w1404) );
	ym3438_AND g_172 (.A(w95), .Z(w4119), .B(w462) );
	ym3438_FA g_173 (.CO(w1445), .S(w893), .CI(w1416), .A(w4119), .B(w890) );
	ym3438_AOI21 g_174 (.A1(w893), .Z(w1442), .B(w1384), .A2(w93) );
	ym3438_SDELAY6 g_175 (.A(w1442), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833), .C3(w57), .C4(w56), .C5(w57), .C6(w56), .C7(w57), .C8(w56), .C9(w57), .C10(w56), .C11(w57), .C12(w56), .nC3(w834), .nC4(w833), .nC5(w834), .nC6(w833), .nC7(w834), .nC8(w833), .nC9(w834), .nC10(w833), .nC11(w834), .nC12(w833), .Q(w895) );
	ym3438_NOR g_176 (.A(w895), .Z(w890), .B(w1388) );
	ym3438_NOT g_177 (.A(w895), .nZ(w1441) );
	ym3438_AON22 g_178 (.A1(w86), .Z(w1440), .B2(w1441), .A2(w891), .B1(w87) );
	ym3438_SR_BIT g_179 (.Q(w1439), .D(w1440), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_180 (.Q(w1438), .D(w1439), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_181 (.Q(w1437), .D(w1438), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_182 (.Q(w1436), .D(w1437), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_183 (.Q(w897), .D(w1436), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_184 (.Q(w891), .D(w897), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SLATCH g_185 (.Q(w899), .nQ(w1433), .D(w1435), .nC(w1393), .C(w1394) );
	ym3438_AON22 g_186 (.A1(w897), .Z(w1435), .B2(w891), .A2(w78), .B1(w79) );
	ym3438_AOI22 g_187 (.A1(w899), .Z(w1432), .B2(w113), .A2(w72), .B1(w73) );
	ym3438_NOT g_188 (.A(w1432), .nZ(w859) );
	ym3438_NOT g_189 (.A(w1433), .nZ(w1434) );
	ym3438_AND g_190 (.A(w458), .Z(w1469), .B(w95) );
	ym3438_FA g_191 (.CO(w1468), .S(w894), .CI(w1445), .A(w1469), .B(w906) );
	ym3438_AOI21 g_192 (.A1(w894), .Z(w4130), .B(w1384), .A2(w93) );
	ym3438_SDELAY6 g_193 (.A(w4130), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833), .C3(w57), .C4(w56), .C5(w57), .C6(w56), .C7(w57), .C8(w56), .C9(w57), .C10(w56), .C11(w57), .C12(w56), .nC3(w834), .nC4(w833), .nC5(w834), .nC6(w833), .nC7(w834), .nC8(w833), .nC9(w834), .nC10(w833), .nC11(w834), .nC12(w833), .Q(w896) );
	ym3438_NOR g_194 (.A(w896), .Z(w906), .B(w1388) );
	ym3438_NOT g_195 (.A(w896), .nZ(w4123) );
	ym3438_AON22 g_196 (.A1(w86), .Z(w1465), .B2(w4123), .A2(w907), .B1(w87) );
	ym3438_SR_BIT g_197 (.Q(w1464), .D(w1465), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_198 (.Q(w1463), .D(w1464), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_199 (.Q(w1462), .D(w1463), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_200 (.Q(w1466), .D(w1462), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_201 (.Q(w898), .D(w1466), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_202 (.Q(w907), .D(w898), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SLATCH g_203 (.Q(w900), .nQ(w1461), .D(w1467), .nC(w1393), .C(w1394) );
	ym3438_AON22 g_204 (.A1(w898), .Z(w1467), .B2(w907), .A2(w78), .B1(w79) );
	ym3438_AOI22 g_205 (.A1(w900), .Z(w1460), .B2(w107), .A2(w72), .B1(w73) );
	ym3438_NOT g_206 (.A(w1460), .nZ(w860) );
	ym3438_NOT g_207 (.A(w1461), .nZ(w1444) );
	ym3438_AND g_208 (.A(w96), .Z(w4129), .B(w95) );
	ym3438_FA g_209 (.CO(w97), .S(w94), .CI(w1468), .A(w4129), .B(w91) );
	ym3438_AOI21 g_210 (.A1(w94), .Z(w92), .B(w1384), .A2(w93) );
	ym3438_SDELAY6 g_211 (.A(w92), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833), .C3(w57), .C4(w56), .C5(w57), .C6(w56), .C7(w57), .C8(w56), .C9(w57), .C10(w56), .C11(w57), .C12(w56), .nC3(w834), .nC4(w833), .nC5(w834), .nC6(w833), .nC7(w834), .nC8(w833), .nC9(w834), .nC10(w833), .nC11(w834), .nC12(w833), .Q(w89) );
	ym3438_NOR g_212 (.A(w89), .Z(w91), .B(w1388) );
	ym3438_NOT g_213 (.A(w89), .nZ(w88) );
	ym3438_AON22 g_214 (.A1(w86), .Z(w84), .B2(w88), .A2(w85), .B1(w87) );
	ym3438_SR_BIT g_215 (.Q(w83), .D(w84), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_216 (.Q(w82), .D(w83), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_217 (.Q(w81), .D(w82), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_218 (.Q(w80), .D(w81), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_219 (.Q(w77), .D(w80), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_220 (.Q(w85), .D(w77), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SLATCH g_221 (.Q(w1459), .nQ(w4118), .D(w76), .nC(w1393), .C(w1394) );
	ym3438_AON22 g_222 (.A1(w77), .Z(w76), .B2(w85), .A2(w78), .B1(w79) );
	ym3438_AOI22 g_223 (.A1(w1459), .Z(w71), .B2(w74), .A2(w72), .B1(w73) );
	ym3438_NOT g_224 (.A(w71), .nZ(w70) );
	ym3438_NOT g_225 (.A(w4118), .nZ(w75) );
	ym3438_AND g_226 (.A(w457), .Z(w1481), .B(w95) );
	ym3438_FA g_227 (.CO(w1482), .S(w1480), .CI(w97), .A(w1481), .B(w915) );
	ym3438_AOI21 g_228 (.A1(w1480), .Z(w1479), .B(w1384), .A2(w93) );
	ym3438_SDELAY6 g_229 (.A(w1479), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833), .C3(w57), .C4(w56), .C5(w57), .C6(w56), .C7(w57), .C8(w56), .C9(w57), .C10(w56), .C11(w57), .C12(w56), .nC3(w834), .nC4(w833), .nC5(w834), .nC6(w833), .nC7(w834), .nC8(w833), .nC9(w834), .nC10(w833), .nC11(w834), .nC12(w833), .Q(w90) );
	ym3438_NOR g_230 (.A(w90), .Z(w915), .B(w1388) );
	ym3438_NOT g_231 (.A(w90), .nZ(w4122) );
	ym3438_AON22 g_232 (.A1(w86), .Z(w1478), .B2(w4122), .A2(w914), .B1(w87) );
	ym3438_SR_BIT g_233 (.Q(w1477), .D(w1478), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_234 (.Q(w1476), .D(w1477), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_235 (.Q(w1475), .D(w1476), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_236 (.Q(w1474), .D(w1475), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_237 (.Q(w912), .D(w1474), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_238 (.Q(w914), .D(w912), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SLATCH g_239 (.Q(w913), .nQ(w1473), .D(w4131), .nC(w1393), .C(w1394) );
	ym3438_AON22 g_240 (.A1(w912), .Z(w4131), .B2(w914), .A2(w78), .B1(w79) );
	ym3438_AOI22 g_241 (.A1(w913), .Z(w1471), .B2(w1472), .A2(w72), .B1(w73) );
	ym3438_NOT g_242 (.A(w1471), .nZ(w858) );
	ym3438_NOT g_243 (.A(w1473), .nZ(w917) );
	ym3438_AND g_244 (.A(w69), .Z(w4128), .B(w95) );
	ym3438_FA g_245 (.CO(w1458), .S(w910), .CI(w1482), .A(w4128), .B(w67) );
	ym3438_AOI21 g_246 (.A1(w910), .Z(w68), .B(w1384), .A2(w93) );
	ym3438_SDELAY6 g_247 (.A(w68), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833), .C3(w57), .C4(w56), .C5(w57), .C6(w56), .C7(w57), .C8(w56), .C9(w57), .C10(w56), .C11(w57), .C12(w56), .nC3(w834), .nC4(w833), .nC5(w834), .nC6(w833), .nC7(w834), .nC8(w833), .nC9(w834), .nC10(w833), .nC11(w834), .nC12(w833), .Q(w66) );
	ym3438_NOR g_248 (.A(w1388), .Z(w67), .B(w66) );
	ym3438_NOT g_249 (.A(w66), .nZ(w65) );
	ym3438_AON22 g_250 (.Z(w62), .B2(w65), .A2(w64), .A1(w86), .B1(w87) );
	ym3438_SR_BIT g_251 (.Q(w61), .D(w62), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_252 (.Q(w60), .D(w61), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_253 (.Q(w59), .D(w60), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_254 (.Q(w58), .D(w59), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_255 (.Q(w55), .D(w58), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_256 (.Q(w64), .D(w55), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SLATCH g_257 (.Q(w52), .nQ(w1419), .D(w1303), .nC(w1393), .C(w1394) );
	ym3438_AON22 g_258 (.Z(w1303), .B2(w64), .A2(w78), .A1(w55), .B1(w79) );
	ym3438_AOI22 g_259 (.Z(w4124), .B2(w53), .A2(w72), .A1(w52), .B1(w73) );
	ym3438_NOT g_260 (.nZ(w857), .A(w4124) );
	ym3438_NOT g_261 (.nZ(w54), .A(w1419) );
	ym3438_AND g_262 (.A(w986), .Z(w4127), .B(w95) );
	ym3438_FA g_263 (.CO(w1431), .S(w1457), .CI(w1458), .A(w4127), .B(w908) );
	ym3438_AOI21 g_264 (.A1(w93), .Z(w1456), .B(w1384), .A2(w1457) );
	ym3438_SDELAY6 g_265 (.A(w1456), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833), .C3(w57), .C4(w56), .C5(w57), .C6(w56), .C7(w57), .C8(w56), .C9(w57), .C10(w56), .C11(w57), .C12(w56), .nC3(w834), .nC4(w833), .nC5(w834), .nC6(w833), .nC7(w834), .nC8(w833), .nC9(w834), .nC10(w833), .nC11(w834), .nC12(w833), .Q(w1455) );
	ym3438_NOR g_266 (.A(w1388), .Z(w908), .B(w1455) );
	ym3438_NOT g_267 (.A(w1455), .nZ(w4125) );
	ym3438_AON22 g_268 (.Z(w1453), .B2(w4125), .A2(w909), .A1(w86), .B1(w87) );
	ym3438_SR_BIT g_269 (.Q(w1452), .D(w1453), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_270 (.Q(w1451), .D(w1452), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_271 (.Q(w1450), .D(w1451), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_272 (.Q(w1454), .D(w1450), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_273 (.Q(w904), .D(w1454), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_274 (.Q(w909), .D(w904), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SLATCH g_275 (.Q(w1447), .nQ(w1448), .D(w1449), .nC(w1393), .C(w1394) );
	ym3438_AON22 g_276 (.Z(w1449), .B2(w909), .A2(w78), .A1(w904), .B1(w79) );
	ym3438_AOI22 g_277 (.Z(w1446), .B2(w902), .A2(w72), .A1(w1447), .B1(w73) );
	ym3438_NOT g_278 (.nZ(w855), .A(w1446) );
	ym3438_NOT g_279 (.nZ(w1443), .A(w1448) );
	ym3438_AND g_280 (.A(w987), .Z(w4126), .B(w95) );
	ym3438_FA g_281 (.CO(w1402), .S(w1430), .CI(w1431), .A(w4126), .B(w892) );
	ym3438_AOI21 g_282 (.A1(w93), .Z(w1429), .B(w1384), .A2(w1430) );
	ym3438_SDELAY6 g_283 (.A(w1429), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833), .C3(w57), .C4(w56), .C5(w57), .C6(w56), .C7(w57), .C8(w56), .C9(w57), .C10(w56), .C11(w57), .C12(w56), .nC3(w834), .nC4(w833), .nC5(w834), .nC6(w833), .nC7(w834), .nC8(w833), .nC9(w834), .nC10(w833), .nC11(w834), .nC12(w833), .Q(w1428) );
	ym3438_NOR g_284 (.A(w1388), .Z(w892), .B(w1428) );
	ym3438_NOT g_285 (.A(w1428), .nZ(w1427) );
	ym3438_AON22 g_286 (.Z(w1426), .B2(w1427), .A2(w63), .A1(w86), .B1(w87) );
	ym3438_SR_BIT g_287 (.Q(w1425), .D(w1426), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_288 (.Q(w1424), .D(w1425), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_289 (.Q(w1423), .D(w1424), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_290 (.Q(w1422), .D(w1423), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_291 (.Q(w903), .D(w1422), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_292 (.Q(w63), .D(w903), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SLATCH g_293 (.Q(w905), .nQ(w1420), .D(w1421), .nC(w1393), .C(w1394) );
	ym3438_AON22 g_294 (.Z(w1421), .B2(w63), .A2(w78), .A1(w903), .B1(w79) );
	ym3438_AOI22 g_295 (.Z(w4101), .B2(w901), .A2(w72), .A1(w905), .B1(w73) );
	ym3438_NOT g_296 (.nZ(w854), .A(w4101) );
	ym3438_NOT g_297 (.nZ(w1418), .A(w1420) );
	ym3438_NOT g_298 (.nZ(w885), .A(w1169) );
	ym3438_AON22 g_299 (.Z(w4100), .B2(w885), .A2(w72), .A1(w865), .B1(w73) );
	ym3438_NOT g_300 (.nZ(w1170), .A(w1392) );
	ym3438_SLATCH g_301 (.Q(w865), .nQ(w1392), .D(w1395), .nC(w1393), .C(w1394) );
	ym3438_AON22 g_302 (.Z(w1395), .B2(w889), .A2(w78), .A1(w866), .B1(w79) );
	ym3438_SR_BIT g_303 (.Q(w889), .D(w866), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_304 (.Q(w866), .D(w1396), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_305 (.Q(w1396), .D(w1397), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_306 (.Q(w1397), .D(w1398), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_307 (.Q(w1398), .D(w1399), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_SR_BIT g_308 (.Q(w1399), .D(w1400), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833) );
	ym3438_AON22 g_309 (.Z(w1400), .B2(w1401), .A2(w889), .A1(w86), .B1(w87) );
	ym3438_NOT g_310 (.A(w867), .nZ(w1401) );
	ym3438_NOR g_311 (.A(w867), .Z(w868), .B(w1388) );
	ym3438_SDELAY6 g_312 (.A(w4117), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833), .C3(w57), .C4(w56), .C5(w57), .C6(w56), .C7(w57), .C8(w56), .C9(w57), .C10(w56), .C11(w57), .C12(w56), .nC3(w834), .nC4(w833), .nC5(w834), .nC6(w833), .nC7(w834), .nC8(w833), .nC9(w834), .nC10(w833), .nC11(w834), .nC12(w833), .Q(w867) );
	ym3438_AOI21 g_313 (.A2(w1383), .Z(w4117), .B(w869), .A1(w870) );
	ym3438_NOT g_314 (.A(w869), .nZ(w93) );
	ym3438_FA g_315 (.S(w870), .CI(w1402), .A(w871), .B(w868) );
	ym3438_AND g_316 (.A(w886), .Z(w871), .B(w95) );
	ym3438_AND g_317 (.A(w1470), .Z(w862), .B(w911) );
	ym3438_AND g_318 (.A(w1174), .Z(w861), .B(w911) );
	ym3438_OR g_319 (.A(w128), .Z(w911), .B(w916) );
	ym3438_NOT g_320 (.A(w1167), .nZ(w916) );
	ym3438_NOT g_321 (.nZ(w853), .A(w4100) );
	ym3438_NOT g_322 (.A(w216), .nZ(w1524) );
	ym3438_NOT g_323 (.A(w213), .nZ(w1523) );
	ym3438_NOT g_324 (.A(w217), .nZ(w1522) );
	ym3438_NOT g_325 (.A(w212), .nZ(w1521) );
	ym3438_NOT g_326 (.A(w1524), .nZ(w104) );
	ym3438_NOT g_327 (.A(w1523), .nZ(w103) );
	ym3438_NOT g_328 (.A(w1522), .nZ(w106) );
	ym3438_NOT g_329 (.A(w1521), .nZ(w105) );
	ym3438_SR_BIT g_330 (.Q(w920), .D(w1170), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_SR_BIT g_331 (.Q(w957), .D(w1418), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_SR_BIT g_332 (.Q(w921), .D(w1443), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_SR_BIT g_333 (.Q(w922), .D(w54), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_SR_BIT g_334 (.Q(w923), .D(w917), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_SR_BIT g_335 (.Q(w1511), .D(w4368), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_SR_BIT g_336 (.Q(w1512), .D(w1404), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_SR_BIT g_337 (.Q(w1513), .D(w1434), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_SR_BIT g_338 (.Q(w1517), .D(w1444), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_SR_BIT g_339 (.Q(w1519), .D(w75), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_SR_BIT g_340 (.Q(w1509), .D(w4369), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_SR_BIT g_341 (.Q(w124), .D(w4371), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_SR_BIT g_342 (.Q(w115), .D(w122), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_COMP_STR g_343 (.A(w1511), .Z(w873) );
	ym3438_COMP_STR g_344 (.A(w1509), .Z(w1508) );
	ym3438_COMP_STR g_345 (.A(w131), .Z(w128) );
	ym3438_SR_BIT g_346 (.Q(w131), .D(w4370), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_COMP_STR g_347 (.A(w124), .Z(w127) );
	ym3438_NOR g_348 (.A(w118), .Z(w122), .B(w102) );
	ym3438_COMP_STR g_349 (.A(w115), .Z(w114) );
	ym3438_COMP_STR g_350 (.A(w109), .Z(w113) );
	ym3438_SR_BIT g_351 (.Q(w109), .D(w4372), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_COMP_STR g_352 (.A(w99), .Z(w107) );
	ym3438_SR_BIT g_353 (.Q(w99), .D(w4373), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_COMP_STR g_354 (.A(w1506), .Z(w74) );
	ym3438_SR_BIT g_355 (.Q(w1506), .D(w4374), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_COMP_STR g_356 (.A(w1505), .Z(w1472) );
	ym3438_SR_BIT g_357 (.Q(w1505), .D(w4375), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_COMP_STR g_358 (.A(w1503), .Z(w53) );
	ym3438_SR_BIT g_359 (.Q(w1503), .D(w4376), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_COMP_STR g_360 (.A(w1502), .Z(w902) );
	ym3438_SR_BIT g_361 (.Q(w1502), .D(w4377), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_COMP_STR g_362 (.A(w1500), .Z(w901) );
	ym3438_SR_BIT g_363 (.Q(w1500), .D(w4378), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_COMP_STR g_364 (.A(w1496), .Z(w1495) );
	ym3438_SR_BIT g_365 (.Q(w1496), .D(w4379), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_COMP_STR g_366 (.A(w1494), .Z(w1139) );
	ym3438_SR_BIT g_367 (.Q(w1494), .D(w4380), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_COMP_STR g_368 (.A(w1492), .Z(w1493) );
	ym3438_SR_BIT g_369 (.Q(w1492), .D(w4381), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_COMP_STR g_370 (.A(w1490), .Z(w918) );
	ym3438_SR_BIT g_371 (.Q(w1490), .D(w4382), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_COMP_STR g_372 (.A(w1489), .Z(w919) );
	ym3438_SR_BIT g_373 (.Q(w1489), .D(w4383), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_COMP_STR g_374 (.A(w1488), .Z(w263) );
	ym3438_SR_BIT g_375 (.Q(w1488), .D(w4384), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_COMP_STR g_376 (.A(w1487), .Z(w1172) );
	ym3438_SR_BIT g_377 (.Q(w1487), .D(w4385), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_COMP_STR g_378 (.A(w1497), .Z(w864) );
	ym3438_NOR g_379 (.A(w941), .Z(w1498), .B(w102) );
	ym3438_SR_BIT g_380 (.Q(w1497), .D(w1498), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_SR_BIT g_381 (.Q(w943), .D(w1499), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_NOR g_382 (.A(w102), .Z(w1499), .B(w944) );
	ym3438_NOT g_383 (.A(w943), .nZ(w1169) );
	ym3438_NOT g_384 (.A(w100), .nZ(w942) );
	ym3438_NOT g_385 (.nZ(w102), .A(w214) );
	ym3438_AON22 g_386 (.A1(w955), .Z(w964), .B2(w458), .A2(w957), .B1(w956) );
	ym3438_AON22 g_387 (.A1(w955), .Z(w965), .B2(w462), .A2(w921), .B1(w956) );
	ym3438_AON22 g_388 (.A1(w955), .Z(w966), .B2(w461), .A2(w922), .B1(w956) );
	ym3438_AON22 g_389 (.A1(w955), .Z(w1520), .B2(w460), .A2(w923), .B1(w956) );
	ym3438_AON22 g_390 (.A1(w955), .Z(w1518), .B2(w459), .A2(w1519), .B1(w956) );
	ym3438_AON22 g_391 (.A1(w955), .Z(w1514), .B2(w454), .A2(w1512), .B1(w956) );
	ym3438_AON22 g_392 (.A1(w955), .Z(w1515), .B2(w455), .A2(w1513), .B1(w956) );
	ym3438_AON22 g_393 (.A1(w955), .Z(w1516), .B2(w456), .A2(w1517), .B1(w956) );
	ym3438_COMP_STR g_394 (.A(w1483), .Z(w1484) );
	ym3438_NOR g_395 (.A(w927), .Z(w1486), .B(w102) );
	ym3438_SR_BIT g_396 (.Q(w1483), .D(w1486), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_NOT g_397 (.A(w1485), .nZ(w926) );
	ym3438_AND3 g_398 (.A(w121), .Z(w1485), .B(w120), .C(w973) );
	ym3438_AOI22 g_399 (.A1(w926), .Z(w927), .B2(w123), .A2(w1483), .B1(w1485) );
	ym3438_NOT g_400 (.A(w1485), .nZ(w928) );
	ym3438_NOR g_401 (.A(w929), .Z(w4385), .B(w102) );
	ym3438_AOI22 g_402 (.A1(w928), .Z(w929), .B2(w961), .A2(w1487), .B1(w1485) );
	ym3438_NOT g_403 (.A(w1485), .nZ(w925) );
	ym3438_NOR g_404 (.A(w930), .Z(w4384), .B(w102) );
	ym3438_AOI22 g_405 (.A1(w925), .Z(w930), .B2(w132), .A2(w1488), .B1(w1485) );
	ym3438_AOI22 g_406 (.A1(w1491), .Z(w932), .B2(w959), .A2(w1490), .B1(w1485) );
	ym3438_AOI22 g_407 (.A1(w924), .Z(w931), .B2(w960), .A2(w1489), .B1(w1485) );
	ym3438_NOR g_409 (.A(w931), .Z(w4383), .B(w102) );
	ym3438_NOT g_410 (.A(w1485), .nZ(w1491) );
	ym3438_NOR g_411 (.A(w932), .Z(w4382), .B(w102) );
	ym3438_AOI22 g_412 (.A1(w933), .Z(w934), .B2(w958), .A2(w1492), .B1(w1485) );
	ym3438_NOT g_413 (.A(w1485), .nZ(w933) );
	ym3438_NOR g_414 (.A(w934), .Z(w4381), .B(w102) );
	ym3438_AOI22 g_415 (.A1(w935), .Z(w936), .B2(w108), .A2(w1494), .B1(w1485) );
	ym3438_NOT g_416 (.A(w1485), .nZ(w935) );
	ym3438_NOR g_417 (.A(w936), .Z(w4380), .B(w102) );
	ym3438_AOI22 g_418 (.A1(w937), .Z(w938), .B2(w112), .A2(w1496), .B1(w1485) );
	ym3438_NOT g_419 (.A(w1485), .nZ(w937) );
	ym3438_NOR g_420 (.A(w938), .Z(w4379), .B(w102) );
	ym3438_AOI22 g_421 (.A1(w1501), .Z(w945), .B2(w961), .A2(w1500), .B1(w100) );
	ym3438_NOT g_422 (.A(w100), .nZ(w1501) );
	ym3438_NOR g_423 (.A(w945), .Z(w4378), .B(w102) );
	ym3438_AOI22 g_424 (.A1(w946), .Z(w947), .B2(w132), .A2(w1502), .B1(w100) );
	ym3438_NOT g_425 (.A(w100), .nZ(w946) );
	ym3438_NOR g_426 (.A(w947), .Z(w4377), .B(w102) );
	ym3438_AOI22 g_427 (.A1(w948), .Z(w1504), .B2(w960), .A2(w1503), .B1(w100) );
	ym3438_NOT g_428 (.A(w100), .nZ(w948) );
	ym3438_NOR g_429 (.A(w1504), .Z(w4376), .B(w102) );
	ym3438_AOI22 g_430 (.A1(w949), .Z(w950), .B2(w959), .A2(w1505), .B1(w100) );
	ym3438_NOT g_431 (.A(w100), .nZ(w949) );
	ym3438_NOR g_432 (.A(w950), .Z(w4375), .B(w102) );
	ym3438_AOI22 g_433 (.A1(w951), .Z(w952), .B2(w958), .A2(w1506), .B1(w100) );
	ym3438_NOT g_434 (.A(w100), .nZ(w951) );
	ym3438_NOR g_435 (.A(w952), .Z(w4374), .B(w102) );
	ym3438_AOI22 g_436 (.A1(w101), .Z(w98), .B2(w108), .A2(w99), .B1(w100) );
	ym3438_NOT g_437 (.A(w100), .nZ(w101) );
	ym3438_NOR g_438 (.A(w98), .Z(w4373), .B(w102) );
	ym3438_AOI22 g_439 (.A1(w110), .Z(w111), .B2(w112), .A2(w109), .B1(w100) );
	ym3438_NOT g_440 (.A(w100), .nZ(w110) );
	ym3438_NOR g_441 (.A(w111), .Z(w4372), .B(w102) );
	ym3438_NOT g_442 (.A(w117), .nZ(w116) );
	ym3438_AOI22 g_443 (.A1(w125), .Z(w126), .B2(w961), .A2(w124), .B1(w117) );
	ym3438_NOT g_444 (.A(w117), .nZ(w125) );
	ym3438_NOR g_445 (.A(w126), .Z(w4371), .B(w102) );
	ym3438_AOI22 g_446 (.A1(w129), .Z(w130), .B2(w132), .A2(w131), .B1(w117) );
	ym3438_NOT g_447 (.A(w117), .nZ(w129) );
	ym3438_NOR g_448 (.A(w130), .Z(w4370), .B(w102) );
	ym3438_AOI22 g_449 (.A1(w954), .Z(w1507), .B2(w960), .A2(w1509), .B1(w117) );
	ym3438_NOT g_450 (.A(w117), .nZ(w954) );
	ym3438_NOR g_451 (.A(w1507), .Z(w4369), .B(w102) );
	ym3438_AOI22 g_452 (.A1(w953), .Z(w1510), .B2(w959), .A2(w1511), .B1(w117) );
	ym3438_NOT g_453 (.A(w117), .nZ(w953) );
	ym3438_NOR g_454 (.A(w1510), .Z(w4368), .B(w102) );
	ym3438_COMP_WE g_455 (.A(w1508), .Z(w955), .nZ(w956) );
	ym3438_AND3 g_456 (.A(w121), .Z(w117), .B(w120), .C(w119) );
	ym3438_AOI22 g_457 (.A1(w116), .Z(w118), .B2(w123), .A2(w115), .B1(w117) );
	ym3438_AND3 g_458 (.A(w121), .Z(w100), .B(w120), .C(w970) );
	ym3438_AOI22 g_459 (.A1(w942), .Z(w944), .B2(w4395), .A2(w943), .B1(w100) );
	ym3438_NOT g_460 (.A(w123), .nZ(w4395) );
	ym3438_NOT g_461 (.A(w939), .nZ(w940) );
	ym3438_AND3 g_462 (.A(w121), .Z(w939), .B(w120), .C(w972) );
	ym3438_AOI22 g_463 (.A1(w940), .Z(w941), .B2(w123), .A2(w1497), .B1(w939) );
	ym3438_NOT g_464 (.A(w1495), .nZ(w4015) );
	ym3438_AON22 g_465 (.A1(w4015), .Z(w975), .B2(w963), .A2(w962), .B1(w1495) );
	ym3438_SR_BIT g_466 (.Q(w977), .D(w102), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_CELL50 g_467 (.A(w977), .Z(w112), .B(1'b0) );
	ym3438_CELL50 g_468 (.A(w977), .Z(w108), .B(1'b0) );
	ym3438_CELL50 g_469 (.A(w977), .Z(w958), .B(1'b0) );
	ym3438_CELL50 g_470 (.A(w977), .Z(w959), .B(1'b0) );
	ym3438_CELL50 g_471 (.A(w977), .Z(w960), .B(1'b0) );
	ym3438_CELL50 g_472 (.A(w977), .Z(w132), .B(1'b0) );
	ym3438_CELL50 g_473 (.A(w977), .Z(w961), .B(1'b0) );
	ym3438_CELL50 g_474 (.A(w977), .Z(w123), .B(1'b0) );
	ym3438_AON22 g_475 (.A1(w976), .Z(w984), .B2(w964), .A2(w1538), .B1(w1539) );
	ym3438_TRI g_476 (.A(w984), .Z(w1078), .E(w967) );
	ym3438_TRI g_477 (.A(w983), .Z(w1151), .E(w967) );
	ym3438_AON22 g_478 (.A1(w975), .Z(w983), .B2(w965), .A2(w1538), .B1(w1539) );
	ym3438_AON22 g_479 (.A1(w4016), .Z(w985), .B2(w966), .A2(w1538), .B1(w1539) );
	ym3438_AON22 g_480 (.A1(w886), .Z(w4016), .B2(1'b0), .A2(w1540), .B1(w1541) );
	ym3438_TRI g_481 (.A(w985), .Z(w1160), .E(w967) );
	ym3438_AON22 g_482 (.A1(w987), .Z(w4017), .B2(1'b0), .A2(w1540), .B1(w1541) );
	ym3438_AON22 g_483 (.A1(w4017), .Z(w1545), .B2(w1520), .A2(w1538), .B1(w1539) );
	ym3438_TRI g_484 (.A(w1545), .Z(w1159), .E(w967) );
	ym3438_AON22 g_485 (.A1(w986), .Z(w4018), .B2(1'b0), .A2(w1540), .B1(w1541) );
	ym3438_AON22 g_486 (.A1(w4018), .Z(w1544), .B2(w1518), .A2(w1538), .B1(w1539) );
	ym3438_TRI g_487 (.A(w1544), .Z(w1158), .E(w967) );
	ym3438_AON22 g_488 (.A1(w69), .Z(w4019), .B2(1'b0), .A2(w1540), .B1(w1541) );
	ym3438_AON22 g_489 (.A1(w4019), .Z(w1543), .B2(w1516), .A2(w1538), .B1(w1539) );
	ym3438_TRI g_490 (.A(w1543), .Z(w1157), .E(w967) );
	ym3438_TRI g_491 (.A(w1542), .Z(w1155), .E(w967) );
	ym3438_AON22 g_492 (.A1(w4020), .Z(w1542), .B2(w1515), .A2(w1538), .B1(w1539) );
	ym3438_AON22 g_493 (.A1(w457), .Z(w4020), .B2(1'b0), .A2(w1540), .B1(w1541) );
	ym3438_AON22 g_494 (.A1(w96), .Z(w4021), .B2(w920), .A2(w1540), .B1(w1541) );
	ym3438_AON22 g_495 (.A1(w4021), .Z(w978), .B2(w1514), .A2(w1538), .B1(w1539) );
	ym3438_TRI g_496 (.A(w978), .Z(w1156), .E(w967) );
	ym3438_COMP_WE g_497 (.A(w1508), .Z(w1541), .nZ(w1540) );
	ym3438_COMP_WE g_498 (.A(w1484), .Z(w1539), .nZ(w1538) );
	ym3438_AND g_499 (.Z(w967), .B(w1088), .A(w1172) );
	ym3438_NOR5 g_500 (.Z(w1537), .B(w961), .A(w123), .C(w960), .D(w112), .E(w108) );
	ym3438_AND6 g_501 (.Z(w979), .B(w132), .A(w1537), .C(w959), .D(w958), .E(w1103), .F(w120) );
	ym3438_NOT g_502 (.A(w1536), .nZ(w119) );
	ym3438_SR_BIT g_503 (.Q(w1536), .D(w1535), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_AOI21 g_504 (.A1(w1534), .Z(w1535), .B(w979), .A2(w119) );
	ym3438_NOT g_505 (.A(w1103), .nZ(w1534) );
	ym3438_NOR5 g_506 (.Z(w969), .B(w961), .A(w123), .C(w960), .D(w958), .E(w112) );
	ym3438_AND6 g_507 (.Z(w980), .B(w132), .A(w969), .C(w959), .D(w108), .E(w120), .F(w1103) );
	ym3438_NOT g_508 (.A(w1533), .nZ(w970) );
	ym3438_SR_BIT g_509 (.Q(w1533), .D(w1532), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_AOI21 g_510 (.A1(w1531), .Z(w1532), .B(w980), .A2(w970) );
	ym3438_NOR4 g_511 (.Z(w971), .B(w961), .A(w123), .C(w960), .D(w958) );
	ym3438_NOT g_512 (.A(w1103), .nZ(w1531) );
	ym3438_AND7 g_513 (.Z(w981), .B(w132), .A(w971), .C(w959), .D(w108), .E(w112), .F(w1103), .G(w120) );
	ym3438_NOT g_514 (.A(w1530), .nZ(w972) );
	ym3438_SR_BIT g_515 (.Q(w1530), .D(w1529), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_AOI21 g_516 (.A1(w1528), .Z(w1529), .B(w981), .A2(w972) );
	ym3438_NOR6 g_517 (.Z(w974), .B(w961), .A(w123), .C(w960), .D(w959), .E(w958), .F(w108) );
	ym3438_NOT g_518 (.A(w1103), .nZ(w1528) );
	ym3438_AND5 g_519 (.Z(w982), .B(w132), .A(w974), .C(w112), .D(w120), .E(w1103) );
	ym3438_NOT g_520 (.A(w1527), .nZ(w973) );
	ym3438_SR_BIT g_521 (.Q(w1527), .D(w1526), .C1(w103), .C2(w104), .nC1(w105), .nC2(w106) );
	ym3438_AOI21 g_522 (.A1(w1525), .Z(w1526), .B(w982), .A2(w973) );
	ym3438_NOT g_523 (.A(w1103), .nZ(w1525) );
	ym3438_NOR6 g_524 (.Z(w1546), .B(w958), .A(w112), .C(w959), .D(w960), .E(w961), .F(w123) );
	ym3438_AND5 g_525 (.Z(w996), .B(w120), .A(w1103), .C(w132), .D(w108), .E(w1546) );
	ym3438_NOT g_526 (.A(w1547), .nZ(w1014) );
	ym3438_SR_BIT g_527 (.Q(w1547), .D(w4069), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_AOI21 g_528 (.A1(w1014), .Z(w4069), .B(w996), .A2(w1548) );
	ym3438_NOT g_529 (.A(w1103), .nZ(w1548) );
	ym3438_NOR5 g_530 (.Z(w1551), .B(w959), .A(w112), .C(w960), .D(w961), .E(w123) );
	ym3438_AND6 g_531 (.Z(w995), .B(w120), .A(w108), .C(w1103), .D(w958), .E(w132), .F(w1551) );
	ym3438_NOT g_532 (.A(w1549), .nZ(w1012) );
	ym3438_SR_BIT g_533 (.Q(w1549), .D(w4399), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_AOI21 g_534 (.A1(w1012), .Z(w4399), .B(w995), .A2(w1550) );
	ym3438_NOT g_535 (.A(w1103), .nZ(w1550) );
	ym3438_NOT g_536 (.A(w1552), .nZ(w1011) );
	ym3438_SR_BIT g_537 (.Q(w1552), .D(w1554), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_AOI21 g_538 (.A1(w1011), .Z(w1554), .B(w993), .A2(w1553) );
	ym3438_NOT g_539 (.A(w1103), .nZ(w1553) );
	ym3438_NOT g_540 (.A(w1556), .nZ(w1010) );
	ym3438_SR_BIT g_541 (.Q(w1556), .D(w4398), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_AOI21 g_542 (.A1(w1010), .Z(w4398), .B(w992), .A2(w1557) );
	ym3438_NOT g_543 (.A(w1103), .nZ(w1557) );
	ym3438_NOT g_544 (.A(w4400), .nZ(w1009) );
	ym3438_SR_BIT g_545 (.Q(w4400), .D(w4401), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_AOI21 g_546 (.A1(w1009), .Z(w4401), .B(w991), .A2(w1559) );
	ym3438_NOT g_547 (.A(w1103), .nZ(w1559) );
	ym3438_NOT g_548 (.A(w1562), .nZ(w1561) );
	ym3438_SR_BIT g_549 (.Q(w1562), .D(w1564), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_AOI21 g_550 (.A1(w1561), .Z(w1564), .B(w990), .A2(w1563) );
	ym3438_NOT g_551 (.A(w1103), .nZ(w1563) );
	ym3438_AND5 g_552 (.Z(w990), .B(w120), .A(w1103), .C(w959), .D(w132), .E(w1560) );
	ym3438_NOR6 g_553 (.Z(w1560), .B(w108), .A(w958), .C(w112), .D(w960), .E(w961), .F(w123) );
	ym3438_AND5 g_554 (.Z(w991), .B(w120), .A(w1103), .C(w958), .D(w132), .E(w1558) );
	ym3438_NOR6 g_555 (.Z(w1558), .B(w959), .A(w112), .C(w108), .D(w960), .E(w961), .F(w123) );
	ym3438_NOR5 g_556 (.Z(w1555), .B(w959), .A(w108), .C(w961), .D(w960), .E(w123) );
	ym3438_AND6 g_557 (.Z(w992), .B(w120), .A(w1103), .C(w112), .D(w958), .E(w132), .F(w1555) );
	ym3438_NOR4 g_558 (.Z(w994), .B(w959), .A(w960), .C(w961), .D(w123) );
	ym3438_AND7 g_559 (.Z(w993), .B(w1103), .A(w108), .C(w112), .D(w120), .E(w132), .F(w994), .G(w958) );
	ym3438_NOT g_560 (.nZ(w341), .A(w1565) );
	ym3438_CNT_BIT g_561 (.CI(w1006), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1566), .nQ(w1565) );
	ym3438_NOT g_562 (.nZ(w1177), .A(w1567) );
	ym3438_CNT_BIT g_563 (.CI(w1005), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1566), .CO(w1006), .nQ(w1567) );
	ym3438_NOT g_564 (.nZ(w1176), .A(w1568) );
	ym3438_CNT_BIT g_565 (.CI(w1007), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1566), .CO(w1005), .nQ(w1568) );
	ym3438_NOT g_566 (.nZ(w1007), .A(w1569) );
	ym3438_CNT_BIT g_567 (.CI(w1004), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w989), .nQ(w1569) );
	ym3438_NOT g_568 (.nZ(w988), .A(w1570) );
	ym3438_CNT_BIT g_569 (.CI(1'b1), .nQ(w1570), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w989), .CO(w1004) );
	ym3438_OR g_570 (.A(w847), .Z(w1566), .B(w1008) );
	ym3438_OR g_571 (.A(w1566), .Z(w989), .B(w1007) );
	ym3438_XOR g_572 (.A(w341), .Z(w1002), .B(1'b0) );
	ym3438_XOR g_573 (.A(w1177), .Z(w1571), .B(1'b0) );
	ym3438_XOR g_574 (.A(w1176), .Z(w998), .B(w1001) );
	ym3438_XOR g_575 (.A(w1007), .Z(w999), .B(w1000) );
	ym3438_XOR g_576 (.A(w988), .Z(w997), .B(w1572) );
	ym3438_AND g_577 (.A(w132), .Z(w1652), .B(w1610) );
	ym3438_AND g_578 (.A(w960), .Z(w1651), .B(w1610) );
	ym3438_NOT g_579 (.nZ(w1008), .A(w214) );
	ym3438_AOI22 g_580 (.A1(w1649), .Z(w1650), .B2(w959), .A2(w1022), .B1(w1642) );
	ym3438_NOR g_581 (.A(w1008), .Z(w4024), .B(w1650) );
	ym3438_AND3 g_582 (.Z(w1642), .B(w120), .A(w121), .C(w1014) );
	ym3438_AOI22 g_583 (.A1(w1644), .Z(w1643), .B2(w112), .A2(w1042), .B1(w1642) );
	ym3438_NOR g_584 (.A(w1008), .Z(w4023), .B(w1646) );
	ym3438_AOI22 g_585 (.A1(w1645), .Z(w1646), .B2(w108), .A2(w1043), .B1(w1642) );
	ym3438_AOI22 g_586 (.A1(w1647), .Z(w1648), .B2(w958), .A2(w1023), .B1(w1642) );
	ym3438_NOR g_587 (.A(w1008), .Z(w4067), .B(w1648) );
	ym3438_AOI22 g_588 (.A1(w1640), .Z(w1641), .B2(w112), .A2(w1024), .B1(w1624) );
	ym3438_NOR g_589 (.A(w1008), .Z(w4066), .B(w1641) );
	ym3438_AOI22 g_590 (.A1(w1638), .Z(w1639), .B2(w108), .A2(w1025), .B1(w1624) );
	ym3438_NOR g_591 (.A(w1008), .Z(w4065), .B(w1639) );
	ym3438_AOI22 g_592 (.A1(w1636), .Z(w1637), .B2(w958), .A2(w1673), .B1(w1624) );
	ym3438_NOR g_593 (.A(w1008), .Z(w4064), .B(w1637) );
	ym3438_AOI22 g_594 (.A1(w1634), .Z(w1635), .B2(w959), .A2(w1674), .B1(w1624) );
	ym3438_NOR g_595 (.A(w1008), .Z(w4063), .B(w1635) );
	ym3438_NOR5 g_596 (.Z(w4040), .B(w1571), .A(w1002), .C(w998), .D(w999), .E(w997) );
	ym3438_AND3 g_597 (.Z(w1575), .B(w1561), .A(w121), .C(w120) );
	ym3438_AOI22 g_598 (.A1(w1576), .Z(w1015), .B2(w112), .A2(w1572), .B1(w1575) );
	ym3438_AOI22 g_599 (.A1(w1578), .Z(w1016), .B2(w108), .A2(w1000), .B1(w1575) );
	ym3438_NOR g_600 (.A(w1008), .Z(w4041), .B(w1016) );
	ym3438_NOR g_601 (.A(w1008), .Z(w4042), .B(w1017) );
	ym3438_AOI22 g_602 (.A1(w1579), .Z(w1017), .B2(w958), .A2(w1001), .B1(w1575) );
	ym3438_NOR g_603 (.A(w1008), .Z(w4044), .B(w1018) );
	ym3438_AOI22 g_604 (.A1(w1580), .Z(w1018), .B2(w960), .A2(w1688), .B1(w1575) );
	ym3438_NOR g_605 (.A(w1008), .Z(w4043), .B(w1019) );
	ym3438_AOI22 g_606 (.A1(w1581), .Z(w1019), .B2(w123), .A2(w1687), .B1(w1575) );
	ym3438_NOR g_607 (.A(w1008), .Z(w4045), .B(w1020) );
	ym3438_AOI22 g_608 (.A1(w1582), .Z(w1020), .B2(w132), .A2(w1686), .B1(w1575) );
	ym3438_NOR g_609 (.A(w1008), .Z(w4046), .B(w1583) );
	ym3438_AOI22 g_610 (.A1(w1584), .Z(w1583), .B2(w961), .A2(w1684), .B1(w1575) );
	ym3438_AND3 g_611 (.Z(w1585), .B(w120), .A(w121), .C(w1009) );
	ym3438_AOI22 g_612 (.A1(w1586), .Z(w1587), .B2(w123), .A2(w1589), .B1(w1585) );
	ym3438_NOR g_613 (.A(w1008), .Z(w4049), .B(w1591) );
	ym3438_AOI22 g_614 (.A1(w1590), .Z(w1591), .B2(w961), .A2(w1032), .B1(w1585) );
	ym3438_NOR g_615 (.A(w1008), .Z(w4048), .B(w1593) );
	ym3438_AOI22 g_616 (.A1(w1592), .Z(w1593), .B2(w132), .A2(w1033), .B1(w1585) );
	ym3438_AOI22 g_617 (.A1(w1602), .Z(w1603), .B2(w112), .A2(w1031), .B1(w1585) );
	ym3438_NOR g_618 (.A(w1008), .Z(w4047), .B(w1595) );
	ym3438_AOI22 g_619 (.A1(w1594), .Z(w1595), .B2(w960), .A2(w1034), .B1(w1585) );
	ym3438_NOR g_620 (.A(w1008), .Z(w4050), .B(w1597) );
	ym3438_AOI22 g_621 (.A1(w1596), .Z(w1597), .B2(w959), .A2(w1035), .B1(w1585) );
	ym3438_NOR g_622 (.A(w1008), .Z(w4051), .B(w1599) );
	ym3438_AOI22 g_623 (.A1(w1598), .Z(w1599), .B2(w958), .A2(w1036), .B1(w1585) );
	ym3438_NOR g_624 (.A(w1008), .Z(w4052), .B(w1601) );
	ym3438_AOI22 g_625 (.A1(w1600), .Z(w1601), .B2(w108), .A2(w1037), .B1(w1585) );
	ym3438_NOR g_626 (.A(w1008), .Z(w4053), .B(w1603) );
	ym3438_AOI22 g_627 (.A1(w1631), .Z(w1632), .B2(w960), .A2(w1633), .B1(w1624) );
	ym3438_NOR g_628 (.A(w1008), .Z(w4022), .B(w1632) );
	ym3438_AOI22 g_629 (.A1(w1629), .Z(w1630), .B2(w132), .A2(w1026), .B1(w1624) );
	ym3438_NOR g_630 (.A(w1008), .Z(w4062), .B(w1630) );
	ym3438_AOI22 g_631 (.A1(w1627), .Z(w1628), .B2(w961), .A2(w1027), .B1(w1624) );
	ym3438_NOR g_632 (.A(w1008), .Z(w4091), .B(w1628) );
	ym3438_AOI22 g_633 (.A1(w1625), .Z(w1626), .B2(w123), .A2(w1028), .B1(w1624) );
	ym3438_AND3 g_634 (.Z(w1624), .B(w120), .A(w121), .C(w1012) );
	ym3438_AOI22 g_635 (.A1(w1622), .Z(w1623), .B2(w123), .A2(w1040), .B1(w1610) );
	ym3438_NOR g_636 (.A(w1008), .Z(w4060), .B(w1623) );
	ym3438_AOI22 g_637 (.A1(w1620), .Z(w1621), .B2(w961), .A2(w1039), .B1(w1610) );
	ym3438_NOR g_638 (.A(w1008), .Z(w4058), .B(w1621) );
	ym3438_AOI22 g_639 (.A1(w1618), .Z(w1619), .B2(w959), .A2(w1038), .B1(w1610) );
	ym3438_NOR g_640 (.A(w1008), .Z(w4059), .B(w1619) );
	ym3438_AOI22 g_641 (.A1(w1616), .Z(w1617), .B2(w958), .A2(w1029), .B1(w1610) );
	ym3438_NOR g_642 (.A(w1008), .Z(w4057), .B(w1617) );
	ym3438_AOI22 g_643 (.A1(w1614), .Z(w1615), .B2(w108), .A2(w1060), .B1(w1610) );
	ym3438_NOR g_644 (.A(w1008), .Z(w4056), .B(w1615) );
	ym3438_AOI22 g_645 (.A1(w1611), .Z(w1612), .B2(w112), .A2(w1054), .B1(w1610) );
	ym3438_AND3 g_646 (.Z(w1610), .B(w120), .A(w121), .C(w1011) );
	ym3438_AOI22 g_647 (.A1(w1608), .Z(w1609), .B2(w112), .A2(w1030), .B1(w1604) );
	ym3438_NOR g_648 (.A(w1008), .Z(w4055), .B(w1609) );
	ym3438_AOI22 g_649 (.A1(w1605), .Z(w1606), .B2(w108), .A2(w4054), .B1(w1604) );
	ym3438_AND3 g_650 (.Z(w1604), .B(w120), .A(w121), .C(w1010) );
	ym3438_NOT g_651 (.nZ(w1163), .A(w4037) );
	ym3438_NOT g_652 (.nZ(w4037), .A(w212) );
	ym3438_NOT g_653 (.nZ(w4036), .A(w217) );
	ym3438_COMP_STR g_654 (.Z(w1137), .A(w1023) );
	ym3438_COMP_STR g_655 (.Z(w1021), .A(w1022) );
	ym3438_SR_BIT g_656 (.Q(w1066), .D(w1652), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_SR_BIT g_657 (.Q(w1065), .D(w1651), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_SR_BIT g_658 (.Q(w1022), .D(w4024), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_SR_BIT g_659 (.Q(w1023), .D(w4067), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_SR_BIT g_660 (.Q(w1043), .D(w4023), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_SR_BIT g_661 (.Q(w1042), .D(w4068), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOR g_662 (.A(w1643), .Z(w4068), .B(w1008) );
	ym3438_NOT g_663 (.nZ(w1649), .A(w1642) );
	ym3438_NOT g_664 (.nZ(w1647), .A(w1642) );
	ym3438_NOT g_665 (.nZ(w1645), .A(w1642) );
	ym3438_NOT g_666 (.nZ(w1644), .A(w1642) );
	ym3438_SR_BIT g_667 (.Q(w1024), .D(w4066), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_668 (.nZ(w1640), .A(w1624) );
	ym3438_SR_BIT g_669 (.Q(w1025), .D(w4065), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_670 (.nZ(w1638), .A(w1624) );
	ym3438_SR_BIT g_671 (.Q(w1673), .D(w4064), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_672 (.nZ(w1636), .A(w1624) );
	ym3438_SR_BIT g_673 (.Q(w1674), .D(w4063), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_674 (.nZ(w1634), .A(w1624) );
	ym3438_SR_BIT g_675 (.Q(w1633), .D(w4022), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_676 (.nZ(w1631), .A(w1624) );
	ym3438_SR_BIT g_677 (.Q(w1026), .D(w4062), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_678 (.nZ(w1629), .A(w1624) );
	ym3438_SR_BIT g_679 (.Q(w1027), .D(w4091), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_680 (.nZ(w1627), .A(w1624) );
	ym3438_SR_BIT g_681 (.Q(w1028), .D(w4061), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOR g_682 (.A(w1626), .Z(w4061), .B(w1008) );
	ym3438_NOT g_683 (.nZ(w1625), .A(w1624) );
	ym3438_SR_BIT g_684 (.Q(w1040), .D(w4060), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_685 (.nZ(w1622), .A(w1610) );
	ym3438_SR_BIT g_686 (.Q(w1039), .D(w4058), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_687 (.nZ(w1620), .A(w1610) );
	ym3438_SR_BIT g_688 (.Q(w1038), .D(w4059), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_689 (.nZ(w1618), .A(w1610) );
	ym3438_SR_BIT g_690 (.Q(w1029), .D(w4057), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_691 (.nZ(w1616), .A(w1610) );
	ym3438_SR_BIT g_692 (.Q(w1060), .D(w4056), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_693 (.nZ(w1614), .A(w1610) );
	ym3438_SR_BIT g_694 (.Q(w1054), .D(w1613), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOR g_695 (.A(w1612), .Z(w1613), .B(w1008) );
	ym3438_NOT g_696 (.nZ(w1611), .A(w1610) );
	ym3438_SR_BIT g_697 (.Q(w1030), .D(w4055), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_SR_BIT g_698 (.Q(w4054), .D(w1607), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_699 (.nZ(w1608), .A(w1604) );
	ym3438_NOT g_700 (.nZ(w1605), .A(w1604) );
	ym3438_NOR g_701 (.A(w1606), .Z(w1607), .B(w1008) );
	ym3438_SR_BIT g_702 (.Q(w1031), .D(w4053), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_703 (.nZ(w1602), .A(w1585) );
	ym3438_SR_BIT g_704 (.Q(w1037), .D(w4052), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_705 (.nZ(w1600), .A(w1585) );
	ym3438_SR_BIT g_706 (.Q(w1036), .D(w4051), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_707 (.nZ(w1598), .A(w1585) );
	ym3438_SR_BIT g_708 (.Q(w1035), .D(w4050), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_709 (.nZ(w1596), .A(w1585) );
	ym3438_SR_BIT g_710 (.Q(w1034), .D(w4047), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_711 (.nZ(w1594), .A(w1585) );
	ym3438_SR_BIT g_712 (.Q(w1033), .D(w4048), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_713 (.nZ(w1592), .A(w1585) );
	ym3438_SR_BIT g_714 (.Q(w1032), .D(w4049), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_715 (.nZ(w1590), .A(w1585) );
	ym3438_SR_BIT g_716 (.Q(w1589), .D(w1588), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOR g_717 (.A(w1587), .Z(w1588), .B(w1008) );
	ym3438_NOT g_718 (.nZ(w1586), .A(w1585) );
	ym3438_SR_BIT g_719 (.Q(w1684), .D(w4046), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_720 (.nZ(w1584), .A(w1575) );
	ym3438_SR_BIT g_721 (.Q(w1686), .D(w4045), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_722 (.nZ(w1582), .A(w1575) );
	ym3438_SR_BIT g_723 (.Q(w1687), .D(w4043), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_724 (.nZ(w1581), .A(w1575) );
	ym3438_SR_BIT g_725 (.Q(w1688), .D(w4044), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_726 (.nZ(w1580), .A(w1575) );
	ym3438_SR_BIT g_727 (.Q(w1001), .D(w4042), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_728 (.nZ(w1579), .A(w1575) );
	ym3438_SR_BIT g_729 (.Q(w1000), .D(w4041), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_730 (.nZ(w1578), .A(w1575) );
	ym3438_SR_BIT g_731 (.Q(w1572), .D(w1577), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOR g_732 (.A(w1015), .Z(w1577), .B(w1008) );
	ym3438_NOT g_733 (.nZ(w1576), .A(w1575) );
	ym3438_COMP_WE g_734 (.Z(w1573), .A(w4040), .nZ(w1574) );
	ym3438_NOT g_735 (.nZ(w1041), .A(w4038) );
	ym3438_NOT g_736 (.nZ(w1073), .A(w4036) );
	ym3438_NOT g_737 (.nZ(w4039), .A(w1008) );
	ym3438_NOT g_738 (.nZ(w4038), .A(w216) );
	ym3438_NOT g_739 (.nZ(w1690), .A(w213) );
	ym3438_NOT g_740 (.nZ(w1072), .A(w1690) );
	ym3438_AON22 g_741 (.A1(w1574), .Z(w1052), .B2(w1573), .A2(w1682), .B1(w1684) );
	ym3438_AON22 g_742 (.A1(w1574), .Z(w1683), .B2(w1573), .A2(w1050), .B1(w1686) );
	ym3438_AON22 g_743 (.A1(w1574), .Z(w1049), .B2(w1573), .A2(w1048), .B1(w1687) );
	ym3438_AON32 g_744 (.A1(w1574), .Z(w1685), .B2(w1573), .A2(w1689), .B1(w1688), .A3(w4039) );
	ym3438_CNT_BIT_LOAD g_745 (.CI(w1670), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1680), .CO(w1681), .D(w1589), .L(w1679), .nL(w1678) );
	ym3438_CNT_BIT_LOAD g_746 (.CI(w1669), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1680), .CO(w1670), .D(w1032), .L(w1679), .nL(w1678) );
	ym3438_CNT_BIT_LOAD g_747 (.CI(w1668), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1680), .CO(w1669), .D(w1033), .L(w1679), .nL(w1678) );
	ym3438_CNT_BIT_LOAD g_748 (.CI(w1667), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1680), .CO(w1668), .D(w1034), .L(w1679), .nL(w1678) );
	ym3438_CNT_BIT_LOAD g_749 (.CI(w1666), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1680), .CO(w1667), .D(w1035), .L(w1679), .nL(w1678) );
	ym3438_CNT_BIT_LOAD g_750 (.CI(w1665), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1680), .CO(w1666), .D(w1036), .L(w1679), .nL(w1678) );
	ym3438_CNT_BIT_LOAD g_751 (.CI(w1664), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1680), .CO(w1665), .D(w1037), .L(w1679), .nL(w1678) );
	ym3438_CNT_BIT_LOAD g_752 (.CI(w1663), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1680), .CO(w1664), .D(w1031), .L(w1679), .nL(w1678) );
	ym3438_CNT_BIT_LOAD g_753 (.CI(w1662), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1680), .CO(w1663), .D(w4054), .L(w1679), .nL(w1678) );
	ym3438_CNT_BIT_LOAD g_754 (.CI(w1056), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1680), .CO(w1662), .D(w1030), .L(w1679), .nL(w1678) );
	ym3438_CNT_BIT_LOAD g_755 (.CI(w1661), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1671), .CO(w1061), .D(w1028), .nL(w1654), .L(w1653) );
	ym3438_CNT_BIT_LOAD g_756 (.CI(w1660), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1671), .CO(w1661), .D(w1027), .L(w1653), .nL(w1654) );
	ym3438_CNT_BIT_LOAD g_757 (.CI(w1659), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1671), .CO(w1660), .D(w1026), .L(w1653), .nL(w1654) );
	ym3438_CNT_BIT_LOAD g_758 (.CI(w1658), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1671), .CO(w1659), .D(w1633), .L(w1653), .nL(w1654) );
	ym3438_CNT_BIT_LOAD g_759 (.CI(w1657), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1671), .CO(w1658), .D(w1674), .L(w1653), .nL(w1654) );
	ym3438_CNT_BIT_LOAD g_760 (.CI(w1656), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1671), .CO(w1657), .D(w1673), .L(w1653), .nL(w1654) );
	ym3438_CNT_BIT_LOAD g_761 (.CI(w1655), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1671), .CO(w1656), .D(w1025), .L(w1653), .nL(w1654) );
	ym3438_CNT_BIT_LOAD g_762 (.CI(w1064), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1671), .CO(w1655), .D(w1024), .L(w1653), .nL(w1654) );
	ym3438_COMP_STR g_763 (.Z(w1045), .A(w1043) );
	ym3438_COMP_STR g_764 (.Z(w1044), .A(w1042) );
	ym3438_NOT g_765 (.nZ(w1654), .A(w1653) );
	ym3438_NOT g_766 (.nZ(w1675), .A(w1039) );
	ym3438_NOT g_767 (.nZ(w586), .A(w1676) );
	ym3438_NAND g_768 (.A(w1675), .Z(w1676), .B(w1040) );
	ym3438_NOR g_769 (.A(w1039), .Z(w1677), .B(w1040) );
	ym3438_NOT g_770 (.nZ(w1162), .A(w1677) );
	ym3438_NOT g_771 (.nZ(w1678), .A(w1679) );
	ym3438_COMP_STR g_772 (.A(w1047), .Z(w1186) );
	ym3438_AND g_773 (.A(w601), .Z(w1047), .B(w1715) );
	ym3438_NOR g_774 (.A(w1689), .Z(w1716), .B(w1047) );
	ym3438_NOT g_775 (.nZ(w745), .A(w1716) );
	ym3438_SDELAY6 g_776 (.A(w1685), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .C3(w1072), .C4(w1041), .C5(w1072), .C6(w1041), .C7(w1072), .C8(w1041), .C9(w1072), .C10(w1041), .C11(w1072), .C12(w1041), .nC3(w1163), .nC4(w1073), .nC5(w1163), .nC6(w1073), .nC7(w1163), .nC8(w1073), .nC9(w1163), .nC10(w1073), .nC11(w1163), .nC12(w1073), .Q(w1048) );
	ym3438_SDELAY6 g_777 (.A(w1049), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .C3(w1072), .C4(w1041), .C5(w1072), .C6(w1041), .C7(w1072), .C8(w1041), .C9(w1072), .C10(w1041), .C11(w1072), .C12(w1041), .nC3(w1163), .nC4(w1073), .nC5(w1163), .nC6(w1073), .nC7(w1163), .nC8(w1073), .nC9(w1163), .nC10(w1073), .nC11(w1163), .nC12(w1073), .Q(w1050) );
	ym3438_SDELAY6 g_778 (.A(w1683), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .C3(w1072), .C4(w1041), .C5(w1072), .C6(w1041), .C7(w1072), .C8(w1041), .C9(w1072), .C10(w1041), .C11(w1072), .C12(w1041), .nC3(w1163), .nC4(w1073), .nC5(w1163), .nC6(w1073), .nC7(w1163), .nC8(w1073), .nC9(w1163), .nC10(w1073), .nC11(w1163), .nC12(w1073), .Q(w1682) );
	ym3438_SDELAY6 g_779 (.A(w1052), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .C3(w1072), .C4(w1041), .C5(w1072), .C6(w1041), .C7(w1072), .C8(w1041), .C9(w1072), .C10(w1041), .C11(w1072), .C12(w1041), .nC3(w1163), .nC4(w1073), .nC5(w1163), .nC6(w1073), .nC7(w1163), .nC8(w1073), .nC9(w1163), .nC10(w1073), .nC11(w1163), .nC12(w1073), .Q(w1689) );
	ym3438_SLATCH g_780 (.Q(w1715), .D(w1051), .C(w1046), .nC(w1071) );
	ym3438_NOT g_781 (.nZ(w1071), .A(w1046) );
	ym3438_AND g_782 (.A(w586), .Z(w1051), .B(w1714) );
	ym3438_SR_BIT g_783 (.Q(w1710), .D(w1681), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_SR_BIT g_784 (.Q(w1679), .D(w1714), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_SR_BIT g_785 (.Q(w1712), .D(w1053), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_OR g_786 (.A(w1710), .Z(w1714), .B(w1070) );
	ym3438_AND g_787 (.A(w1053), .Z(w1070), .B(w1713) );
	ym3438_NOT g_788 (.nZ(w1713), .A(w1712) );
	ym3438_NOT g_789 (.nZ(w1680), .A(w1053) );
	ym3438_AND g_790 (.A(w1053), .Z(w1069), .B(w1175) );
	ym3438_OR g_791 (.A(w1069), .Z(w1056), .B(w1493) );
	ym3438_NOT g_792 (.nZ(w1068), .A(w1046) );
	ym3438_SLATCH g_793 (.Q(w1053), .D(w1054), .C(w1046), .nC(w1068) );
	ym3438_NOT g_794 (.nZ(w1711), .A(w1692) );
	ym3438_AND3 g_795 (.A(w1029), .Z(w1055), .B(w1710), .C(w1711) );
	ym3438_AOI21 g_796 (.A1(w1705), .Z(w1709), .B(w1055), .A2(w1708) );
	ym3438_NOT g_797 (.nZ(w1708), .A(w1692) );
	ym3438_NOT g_798 (.nZ(w1705), .A(w1706) );
	ym3438_SR_BIT g_799 (.Q(w1706), .D(w1709), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_800 (.nZ(w1067), .A(w1705) );
	ym3438_NOT g_801 (.nZ(w1704), .A(w1691) );
	ym3438_AOI21 g_802 (.A1(w1059), .Z(w1707), .B(w1058), .A2(w1704) );
	ym3438_SR_BIT g_803 (.Q(w1703), .D(w1707), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_NOT g_804 (.nZ(w1059), .A(w1703) );
	ym3438_NOT g_805 (.nZ(w1161), .A(w1059) );
	ym3438_AND3 g_806 (.A(w1057), .Z(w1058), .B(w1038), .C(w1702) );
	ym3438_NOT g_807 (.nZ(w1702), .A(w1691) );
	ym3438_NOT g_808 (.nZ(w1701), .A(w1046) );
	ym3438_SLATCH g_809 (.Q(w1672), .D(w1060), .C(w1046), .nC(w1701) );
	ym3438_SR_BIT g_810 (.Q(w1057), .D(w1061), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_SR_BIT g_811 (.Q(w1700), .D(w1672), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_SR_BIT g_812 (.Q(w1653), .D(w1697), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_OR g_813 (.A(w1698), .Z(w1697), .B(w1057) );
	ym3438_AND g_814 (.A(w1699), .Z(w1698), .B(w1672) );
	ym3438_NOT g_815 (.nZ(w1699), .A(w1700) );
	ym3438_CNT_BIT g_816 (.CI(w1175), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1008), .CO(w1696) );
	ym3438_CNT_BIT g_817 (.CI(w1696), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1008), .CO(w1695) );
	ym3438_CNT_BIT g_818 (.CI(w1695), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1008), .CO(w1694) );
	ym3438_CNT_BIT g_819 (.CI(w1694), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073), .RES(w1008), .CO(w1062) );
	ym3438_OR g_820 (.A(w1066), .Z(w1691), .B(w1008) );
	ym3438_OR g_821 (.A(w1008), .Z(w1692), .B(w1065) );
	ym3438_OR g_822 (.A(w1493), .Z(w1064), .B(w1693) );
	ym3438_AND g_823 (.A(w1672), .Z(w1693), .B(w1063) );
	ym3438_NOT g_824 (.nZ(w1671), .A(w1672) );
	ym3438_SR_BIT g_825 (.Q(w1063), .D(w1062), .C1(w1072), .C2(w1041), .nC1(w1163), .nC2(w1073) );
	ym3438_AND g_826 (.A(1'b1), .Z(w1), .B(w1210) );
	ym3438_AON22 g_827 (.A1(w1210), .Z(w11), .B2(1'b1), .A2(w1199), .B1(w1209) );
	ym3438_AON222 g_828 (.A1(w1210), .Z(w12), .B2(w1199), .A2(w1200), .B1(w1209), .C1(w1212), .C2(1'b1) );
	ym3438_AON2222 g_829 (.A1(w1210), .Z(w13), .B2(w1200), .A2(w1201), .B1(w1209), .C1(w1212), .C2(w1199), .D1(w1211), .D2(1'b1) );
	ym3438_AON2222 g_830 (.A1(w1210), .Z(w1218), .B2(w1201), .A2(w1202), .B1(w1209), .C1(w1212), .C2(w1200), .D1(w1211), .D2(w1199) );
	ym3438_AON2222 g_831 (.A1(w1210), .Z(w1219), .B2(w1202), .A2(w1203), .B1(w1209), .C1(w1212), .C2(w1201), .D1(w1211), .D2(w1200) );
	ym3438_AON2222 g_832 (.A1(w1210), .Z(w1220), .B2(w1203), .A2(w1204), .B1(w1209), .C1(w1212), .C2(w1202), .D1(w1211), .D2(w1201) );
	ym3438_AON2222 g_833 (.A1(w1210), .Z(w1221), .B2(w1204), .A2(w1205), .B1(w1209), .C1(w1212), .C2(w1203), .D1(w1211), .D2(w1202) );
	ym3438_AON2222 g_834 (.A1(w1210), .Z(w1224), .B2(w1205), .A2(w1206), .B1(w1209), .C1(w1212), .C2(w1204), .D1(w1211), .D2(w1203) );
	ym3438_AON2222 g_835 (.A1(w1210), .Z(w1725), .B2(w1206), .A2(w467), .B1(w1209), .C1(w1212), .C2(w1205), .D1(w1211), .D2(w1204) );
	ym3438_AON2222 g_836 (.A1(w1210), .Z(w1724), .B2(w467), .A2(w466), .B1(w1209), .C1(w1212), .C2(w1206), .D1(w1211), .D2(w1205) );
	ym3438_AON222 g_837 (.A1(w1209), .Z(w1222), .B2(w467), .A2(w466), .B1(w1212), .C1(w1211), .C2(w1206) );
	ym3438_AON22 g_838 (.A1(w1212), .Z(w1223), .B2(w467), .A2(w466), .B1(w1211) );
	ym3438_NAND g_839 (.A(w1208), .Z(w1720), .B(w1207) );
	ym3438_NAND g_840 (.A(w1718), .Z(w1721), .B(w1208) );
	ym3438_NAND g_841 (.A(w1719), .Z(w1722), .B(w1207) );
	ym3438_NAND g_842 (.A(w1718), .Z(w1723), .B(w1719) );
	ym3438_NOT g_843 (.A(w1720), .nZ(w1210) );
	ym3438_NOT g_844 (.A(w1721), .nZ(w1209) );
	ym3438_NOT g_845 (.A(w1722), .nZ(w1212) );
	ym3438_NOT g_846 (.A(w1723), .nZ(w1211) );
	ym3438_NOT g_847 (.A(w1208), .nZ(w1719) );
	ym3438_NOT g_848 (.A(w1207), .nZ(w1718) );
	ym3438_NOT g_849 (.A(w464), .nZ(w1214) );
	ym3438_NOT g_850 (.A(w465), .nZ(w1213) );
	ym3438_AND g_851 (.A(w1213), .Z(w4408), .B(w464) );
	ym3438_AND g_852 (.A(w1214), .Z(w1216), .B(w465) );
	ym3438_AND g_853 (.A(w1214), .Z(w1215), .B(w1213) );
	ym3438_AND g_854 (.A(w464), .Z(w1726), .B(w465) );
	ym3438_AON2222 g_855 (.A1(w2), .Z(w1230), .B2(w1224), .A2(w1223), .B1(w1217), .C1(w1216), .C2(w1218), .D1(w1215), .D2(w1) );
	ym3438_AON222 g_856 (.A1(w2), .Z(w1229), .B2(w1221), .A2(w1222), .B1(w1217), .C1(w1216), .C2(w13) );
	ym3438_AON222 g_857 (.A1(w2), .Z(w1228), .B2(w1220), .A2(w1724), .B1(w1217), .C1(w1216), .C2(w12) );
	ym3438_AON222 g_858 (.A1(w2), .Z(w1231), .B2(w1219), .A2(w1725), .B1(w1217), .C1(w1216), .C2(w11) );
	ym3438_AON222 g_859 (.A1(w2), .Z(w1227), .B2(w1218), .A2(w1224), .B1(w1217), .C1(w1216), .C2(w1) );
	ym3438_AON22 g_860 (.A1(w2), .Z(w1232), .B2(w13), .A2(w1221), .B1(w1217) );
	ym3438_AON22 g_861 (.A1(w2), .Z(w1331), .B2(w12), .A2(w1220), .B1(w1217) );
	ym3438_AON22 g_862 (.A1(w2), .Z(w1330), .B2(w11), .A2(w1219), .B1(w1217) );
	ym3438_AND g_863 (.A(w2), .Z(w1328), .B(w1) );
	ym3438_AND g_864 (.A(w11), .Z(w1727), .B(w2) );
	ym3438_AND g_865 (.A(w12), .Z(w1234), .B(w2) );
	ym3438_AND g_866 (.A(w13), .Z(w1329), .B(w2) );
	ym3438_AON22 g_867 (.A1(w2), .Z(w1233), .B2(w1), .A2(w1218), .B1(w1217) );
	ym3438_COMP_STR g_868 (.A(w7), .Z(w1235) );
	ym3438_COMP_STR g_869 (.A(w848), .Z(w1226), .nZ(w1225) );
	ym3438_COMP_STR g_870 (.A(w357), .Z(w356), .nZ(w358) );
	ym3438_COMP_STR g_871 (.A(w848), .Z(w363), .nZ(w361) );
	ym3438_SR_BIT g_872 (.Q(w7), .D(w8), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_873 (.Q(w8), .D(w9), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_874 (.Q(w9), .D(w10), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_COMP_STR g_875 (.A(w1726), .Z(w2) );
	ym3438_COMP_STR g_876 (.A(w4408), .Z(w1217) );
	ym3438_XOR g_877 (.A(w1230), .Z(w1741), .B(w1235) );
	ym3438_HA g_878 (.CO(w368), .S(w1743), .A(w1235), .B(w1741) );
	ym3438_SR_BIT g_879 (.Q(w1779), .D(w1743), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_AON22 g_880 (.A1(w1780), .Z(w1791), .B2(w1779), .A2(w1225), .B1(w1226) );
	ym3438_SDELAY6 g_881 (.A(w1791), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w1780) );
	ym3438_AON22 g_882 (.A1(w373), .Z(w1808), .B2(w1780), .A2(w361), .B1(w363) );
	ym3438_SDELAY6 g_883 (.A(w1808), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w373) );
	ym3438_AON22 g_884 (.A1(w427), .Z(w1824), .B2(w1779), .A2(w358), .B1(w356) );
	ym3438_SDELAY6 g_885 (.A(w1824), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w427) );
	ym3438_AON222 g_886 (.A1(w1779), .Z(w422), .B2(w427), .A2(w444), .B1(w412), .C2(w373), .C1(w439) );
	ym3438_AON22 g_887 (.A1(w1780), .Z(w423), .B2(w1779), .A2(w1828), .B1(w1827) );
	ym3438_FA g_888 (.CO(w1852), .CI(1'b0), .A(w423), .B(w422) );
	ym3438_XOR g_889 (.A(w1229), .Z(w1740), .B(w1235) );
	ym3438_HA g_890 (.CO(w366), .S(w1742), .A(w368), .B(w1740) );
	ym3438_SR_BIT g_891 (.Q(w1777), .D(w1742), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_AON22 g_892 (.A1(w1778), .Z(w1795), .B2(w1777), .A2(w1225), .B1(w1226) );
	ym3438_SDELAY6 g_893 (.A(w1795), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w1778) );
	ym3438_AON22 g_894 (.A1(w372), .Z(w1807), .B2(w1778), .A2(w361), .B1(w363) );
	ym3438_SDELAY6 g_895 (.A(w1807), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w372) );
	ym3438_AON22 g_896 (.A1(w426), .Z(w1823), .B2(w1777), .A2(w358), .B1(w356) );
	ym3438_SDELAY6 g_897 (.A(w1823), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w426) );
	ym3438_AON222 g_898 (.A1(w1777), .Z(w424), .B2(w426), .A2(w444), .B1(w412), .C2(w372), .C1(w439) );
	ym3438_AON22 g_899 (.A1(w1778), .Z(w425), .B2(w1777), .A2(w1828), .B1(w1827) );
	ym3438_FA g_900 (.CO(w1850), .S(w1851), .CI(w1852), .A(w425), .B(w424) );
	ym3438_XOR g_901 (.A(w1228), .Z(w1739), .B(w1235) );
	ym3438_HA g_902 (.CO(w367), .S(w1745), .A(w366), .B(w1739) );
	ym3438_SR_BIT g_903 (.Q(w1775), .D(w1745), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_AON22 g_904 (.A1(w1776), .Z(w1790), .B2(w1775), .A2(w1225), .B1(w1226) );
	ym3438_SDELAY6 g_905 (.A(w1790), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w1776) );
	ym3438_AON22 g_906 (.A1(w429), .Z(w1806), .B2(w1776), .A2(w361), .B1(w363) );
	ym3438_SDELAY6 g_907 (.A(w1806), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w429) );
	ym3438_AON22 g_908 (.A1(w430), .Z(w1822), .B2(w1775), .A2(w358), .B1(w356) );
	ym3438_SDELAY6 g_909 (.A(w1822), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w430) );
	ym3438_AON222 g_910 (.A1(w1775), .Z(w433), .B2(w430), .A2(w444), .B1(w412), .C2(w429), .C1(w439) );
	ym3438_AON22 g_911 (.A1(w1776), .Z(w434), .B2(w1775), .A2(w1828), .B1(w1827) );
	ym3438_FA g_912 (.CO(w1848), .S(w1849), .CI(w1850), .A(w434), .B(w433) );
	ym3438_XOR g_913 (.A(w1231), .Z(w1738), .B(w1235) );
	ym3438_HA g_914 (.CO(w365), .S(w1744), .A(w367), .B(w1738) );
	ym3438_SR_BIT g_915 (.Q(w1773), .D(w1744), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_AON22 g_916 (.A1(w1774), .Z(w1794), .B2(w1773), .A2(w1225), .B1(w1226) );
	ym3438_SDELAY6 g_917 (.A(w1794), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w1774) );
	ym3438_AON22 g_918 (.A1(w428), .Z(w1805), .B2(w1774), .A2(w361), .B1(w363) );
	ym3438_SDELAY6 g_919 (.A(w1805), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w428) );
	ym3438_AON22 g_920 (.A1(w431), .Z(w1821), .B2(w1773), .A2(w358), .B1(w356) );
	ym3438_SDELAY6 g_921 (.A(w1821), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w431) );
	ym3438_AON222 g_922 (.A1(w1773), .Z(w432), .B2(w431), .A2(w444), .B1(w412), .C2(w428), .C1(w439) );
	ym3438_AON22 g_923 (.A1(w1774), .Z(w435), .B2(w1773), .A2(w1828), .B1(w1827) );
	ym3438_FA g_924 (.CO(w1846), .S(w1847), .CI(w1848), .A(w435), .B(w432) );
	ym3438_XOR g_925 (.A(w1227), .Z(w1737), .B(w1235) );
	ym3438_HA g_926 (.CO(w364), .S(w1747), .A(w365), .B(w1737) );
	ym3438_SR_BIT g_927 (.Q(w1771), .D(w1747), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_AON22 g_928 (.A1(w1772), .Z(w1789), .B2(w1771), .A2(w1225), .B1(w1226) );
	ym3438_SDELAY6 g_929 (.A(w1789), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w1772) );
	ym3438_AON22 g_930 (.A1(w362), .Z(w1804), .B2(w1772), .A2(w361), .B1(w363) );
	ym3438_SDELAY6 g_931 (.A(w1804), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w362) );
	ym3438_AON22 g_932 (.A1(w451), .Z(w1820), .B2(w1771), .A2(w358), .B1(w356) );
	ym3438_SDELAY6 g_933 (.A(w1820), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w451) );
	ym3438_AON222 g_934 (.A1(w1771), .Z(w450), .B2(w451), .A2(w444), .B1(w412), .C2(w362), .C1(w439) );
	ym3438_AON22 g_935 (.A1(w1772), .Z(w1829), .B2(w1771), .A2(w1828), .B1(w1827) );
	ym3438_FA g_936 (.CO(w1844), .S(w1845), .CI(w1846), .A(w1829), .B(w450) );
	ym3438_XOR g_937 (.A(w1232), .Z(w1736), .B(w1235) );
	ym3438_HA g_938 (.CO(w360), .S(w1746), .A(w364), .B(w1736) );
	ym3438_SR_BIT g_939 (.Q(w1770), .D(w1746), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_AON22 g_940 (.A1(w371), .Z(w1793), .B2(w1770), .A2(w1225), .B1(w1226) );
	ym3438_SDELAY6 g_941 (.A(w1793), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w371) );
	ym3438_AON22 g_942 (.A1(w1811), .Z(w1803), .B2(w371), .A2(w361), .B1(w363) );
	ym3438_SDELAY6 g_943 (.A(w1803), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w1811) );
	ym3438_AON22 g_944 (.A1(w452), .Z(w1819), .B2(w1770), .A2(w358), .B1(w356) );
	ym3438_SDELAY6 g_945 (.A(w1819), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w452) );
	ym3438_AON222 g_946 (.A1(w1770), .Z(w448), .B2(w452), .A2(w444), .B1(w412), .C2(w1811), .C1(w439) );
	ym3438_AON22 g_947 (.A1(w371), .Z(w449), .B2(w1770), .A2(w1828), .B1(w1827) );
	ym3438_FA g_948 (.CO(w1853), .S(w1843), .CI(w1844), .A(w449), .B(w448) );
	ym3438_XOR g_949 (.A(w1331), .Z(w1735), .B(w1235) );
	ym3438_HA g_950 (.CO(w359), .S(w1749), .A(w360), .B(w1735) );
	ym3438_SR_BIT g_951 (.Q(w1768), .D(w1749), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_AON22 g_952 (.A1(w1769), .Z(w1788), .B2(w1768), .A2(w1225), .B1(w1226) );
	ym3438_SDELAY6 g_953 (.A(w1788), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w1769) );
	ym3438_AON22 g_954 (.A1(w445), .Z(w1802), .B2(w1769), .A2(w361), .B1(w363) );
	ym3438_SDELAY6 g_955 (.A(w1802), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w445) );
	ym3438_AON22 g_956 (.A1(w443), .Z(w1818), .B2(w1768), .A2(w358), .B1(w356) );
	ym3438_SDELAY6 g_957 (.A(w1818), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w443) );
	ym3438_AON222 g_958 (.A1(w1768), .Z(w440), .B2(w443), .A2(w444), .B1(w412), .C2(w445), .C1(w439) );
	ym3438_AON22 g_959 (.A1(w1769), .Z(w441), .B2(w1768), .A2(w1828), .B1(w1827) );
	ym3438_FA g_960 (.CO(w1842), .S(w1854), .CI(w1853), .A(w441), .B(w440) );
	ym3438_XOR g_961 (.A(w1330), .Z(w1734), .B(w1235) );
	ym3438_HA g_962 (.CO(w355), .S(w1748), .A(w359), .B(w1734) );
	ym3438_SR_BIT g_963 (.Q(w1766), .D(w1748), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_AON22 g_964 (.A1(w1767), .Z(w1792), .B2(w1766), .A2(w1225), .B1(w1226) );
	ym3438_SDELAY6 g_965 (.A(w1792), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w1767) );
	ym3438_AON22 g_966 (.A1(w1810), .Z(w1801), .B2(w1767), .A2(w361), .B1(w363) );
	ym3438_SDELAY6 g_967 (.A(w1801), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w1810) );
	ym3438_AON22 g_968 (.A1(w442), .Z(w1817), .B2(w1766), .A2(w358), .B1(w356) );
	ym3438_SDELAY6 g_969 (.A(w1817), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w442) );
	ym3438_AON222 g_970 (.A1(w1766), .Z(w437), .B2(w442), .A2(w444), .B1(w412), .C2(w1810), .C1(w439) );
	ym3438_AON22 g_971 (.A1(w1767), .Z(w438), .B2(w1766), .A2(w1828), .B1(w1827) );
	ym3438_FA g_972 (.CO(w1840), .S(w1841), .CI(w1842), .A(w438), .B(w437) );
	ym3438_XOR g_973 (.A(w1233), .Z(w1732), .B(w1235) );
	ym3438_HA g_974 (.CO(w354), .S(w1751), .A(w355), .B(w1732) );
	ym3438_SR_BIT g_975 (.Q(w1764), .D(w1751), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_AON22 g_976 (.A1(w1765), .Z(w1787), .B2(w1764), .A2(w1225), .B1(w1226) );
	ym3438_SDELAY6 g_977 (.A(w1787), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w1765) );
	ym3438_AON22 g_978 (.A1(w383), .Z(w1800), .B2(w1765), .A2(w361), .B1(w363) );
	ym3438_SDELAY6 g_979 (.A(w1800), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w383) );
	ym3438_AON22 g_980 (.A1(w385), .Z(w1816), .B2(w1764), .A2(w358), .B1(w356) );
	ym3438_SDELAY6 g_981 (.A(w1816), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w385) );
	ym3438_AON222 g_982 (.A1(w1764), .Z(w411), .B2(w385), .A2(w444), .B1(w412), .C2(w383), .C1(w439) );
	ym3438_AON22 g_983 (.A1(w1765), .Z(w413), .B2(w1764), .A2(w1828), .B1(w1827) );
	ym3438_FA g_984 (.CO(w1838), .S(w1839), .CI(w1840), .A(w413), .B(w411) );
	ym3438_XOR g_985 (.A(w1329), .Z(w1731), .B(w1235) );
	ym3438_HA g_986 (.CO(w353), .S(w1750), .A(w354), .B(w1731) );
	ym3438_SR_BIT g_987 (.Q(w1762), .D(w1750), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_AON22 g_988 (.A1(w1763), .Z(w1785), .B2(w1762), .A2(w1225), .B1(w1226) );
	ym3438_SDELAY6 g_989 (.A(w1785), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w1763) );
	ym3438_AON22 g_990 (.A1(w382), .Z(w1799), .B2(w1763), .A2(w361), .B1(w363) );
	ym3438_SDELAY6 g_991 (.A(w1799), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w382) );
	ym3438_AON22 g_992 (.A1(w384), .Z(w1815), .B2(w1762), .A2(w358), .B1(w356) );
	ym3438_SDELAY6 g_993 (.A(w1815), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w384) );
	ym3438_AON222 g_994 (.A1(w1762), .Z(w409), .B2(w384), .A2(w444), .B1(w412), .C2(w382), .C1(w439) );
	ym3438_AON22 g_995 (.A1(w1763), .Z(w410), .B2(w1762), .A2(w1828), .B1(w1827) );
	ym3438_FA g_996 (.CO(w1836), .S(w1837), .CI(w1838), .A(w410), .B(w409) );
	ym3438_XOR g_997 (.A(w919), .Z(w1728), .B(w1235) );
	ym3438_HA g_998 (.S(w1754), .A(w350), .B(w1728) );
	ym3438_SR_BIT g_999 (.Q(w1333), .D(w1754), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_AON22 g_1000 (.A1(w1781), .Z(w1782), .B2(w1333), .A2(w1225), .B1(w1226) );
	ym3438_SDELAY6 g_1001 (.A(w1782), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w1781) );
	ym3438_AON22 g_1002 (.A1(w369), .Z(w1809), .B2(w1781), .A2(w361), .B1(w363) );
	ym3438_SDELAY6 g_1003 (.A(w1809), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w369) );
	ym3438_AON22 g_1004 (.A1(w374), .Z(w1825), .B2(w1333), .A2(w358), .B1(w356) );
	ym3438_SDELAY6 g_1005 (.A(w1825), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w374) );
	ym3438_AON222 g_1006 (.A1(w1333), .Z(w1826), .B2(w374), .A2(w444), .B1(w412), .C2(w369), .C1(w439) );
	ym3438_AON22 g_1007 (.A1(w1781), .Z(w403), .B2(w1333), .A2(w1828), .B1(w1827) );
	ym3438_FA g_1008 (.CO(w386), .S(w1830), .CI(w1831), .A(w403), .B(w1826) );
	ym3438_XOR g_1009 (.A(w1328), .Z(w1729), .B(w1235) );
	ym3438_HA g_1010 (.CO(w350), .S(w1755), .A(w351), .B(w1729) );
	ym3438_SR_BIT g_1011 (.Q(w1756), .D(w1755), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_AON22 g_1012 (.A1(w1757), .Z(w1783), .B2(w1756), .A2(w1225), .B1(w1226) );
	ym3438_SDELAY6 g_1013 (.A(w1783), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w1757) );
	ym3438_AON22 g_1014 (.A1(w370), .Z(w1796), .B2(w1757), .A2(w361), .B1(w363) );
	ym3438_SDELAY6 g_1015 (.A(w1796), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w370) );
	ym3438_AON22 g_1016 (.A1(w375), .Z(w1812), .B2(w1756), .A2(w358), .B1(w356) );
	ym3438_SDELAY6 g_1017 (.A(w1812), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w375) );
	ym3438_AON222 g_1018 (.A1(w1756), .Z(w404), .B2(w375), .A2(w444), .B1(w412), .C2(w370), .C1(w439) );
	ym3438_AON22 g_1019 (.A1(w1757), .Z(w405), .B2(w1756), .A2(w1828), .B1(w1827) );
	ym3438_FA g_1020 (.CO(w1831), .S(w1832), .CI(w406), .A(w405), .B(w404) );
	ym3438_XOR g_1021 (.A(w1727), .Z(w1730), .B(w1235) );
	ym3438_HA g_1022 (.CO(w351), .S(w1752), .A(w352), .B(w1730) );
	ym3438_SR_BIT g_1023 (.Q(w1758), .D(w1752), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_AON22 g_1024 (.A1(w1759), .Z(w1784), .B2(w1758), .A2(w1225), .B1(w1226) );
	ym3438_SDELAY6 g_1025 (.A(w1784), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w1759) );
	ym3438_AON22 g_1026 (.A1(w376), .Z(w1797), .B2(w1759), .A2(w361), .B1(w363) );
	ym3438_SDELAY6 g_1027 (.A(w1797), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w376) );
	ym3438_AON22 g_1028 (.A1(w378), .Z(w1813), .B2(w1758), .A2(w358), .B1(w356) );
	ym3438_SDELAY6 g_1029 (.A(w1813), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w378) );
	ym3438_AON222 g_1030 (.A1(w1758), .Z(w407), .B2(w378), .A2(w444), .B1(w412), .C2(w376), .C1(w439) );
	ym3438_AON22 g_1031 (.A1(w1759), .Z(w380), .B2(w1758), .A2(w1828), .B1(w1827) );
	ym3438_FA g_1032 (.CO(w406), .S(w1833), .CI(w1834), .A(w380), .B(w407) );
	ym3438_XOR g_1033 (.A(w1234), .Z(w1733), .B(w1235) );
	ym3438_HA g_1034 (.CO(w352), .S(w1753), .A(w353), .B(w1733) );
	ym3438_SR_BIT g_1035 (.Q(w1760), .D(w1753), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_AON22 g_1036 (.A1(w1761), .Z(w1786), .B2(w1760), .A2(w1225), .B1(w1226) );
	ym3438_SDELAY6 g_1037 (.A(w1786), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w1761) );
	ym3438_AON22 g_1038 (.A1(w377), .Z(w1798), .B2(w1761), .A2(w361), .B1(w363) );
	ym3438_SDELAY6 g_1039 (.A(w1798), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w377) );
	ym3438_AON22 g_1040 (.A1(w379), .Z(w1814), .B2(w1760), .A2(w358), .B1(w356) );
	ym3438_SDELAY6 g_1041 (.A(w1814), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .C11(w6), .C12(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .nC11(w4), .nC12(w3), .Q(w379) );
	ym3438_AON222 g_1042 (.A1(w1760), .Z(w408), .B2(w379), .A2(w444), .B1(w412), .C2(w377), .C1(w439) );
	ym3438_AON22 g_1043 (.A1(w1761), .Z(w381), .B2(w1760), .A2(w1828), .B1(w1827) );
	ym3438_FA g_1044 (.CO(w1834), .S(w1835), .CI(w1836), .A(w381), .B(w408) );
	ym3438_COMP_STR g_1045 (.A(w436), .Z(w1828) );
	ym3438_COMP_STR g_1046 (.Z(w1827), .A(w447) );
	ym3438_COMP_STR g_1047 (.Z(w444), .A(w446) );
	ym3438_COMP_STR g_1048 (.A(w357), .Z(w439) );
	ym3438_COMP_STR g_1049 (.Z(w412), .A(w414) );
	ym3438_SR_BIT g_1050 (.Q(w401), .D(w1830), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1051 (.Q(w1332), .D(w1832), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BIT g_1052 (.Q(w453), .D(w1833), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1053 (.Q(w1264), .D(w1835), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BIT g_1054 (.Q(w1260), .D(w1837), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1055 (.Q(w1261), .D(w1839), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BIT g_1056 (.Q(w420), .D(w1841), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1057 (.Q(w419), .D(w1854), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BIT g_1058 (.Q(w418), .D(w1843), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1059 (.Q(w417), .D(w1845), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BIT g_1060 (.Q(w416), .D(w1847), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1061 (.Q(w415), .D(w1849), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BIT g_1062 (.Q(w1249), .D(w1851), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_COMP_STR g_1063 (.A(w1779), .Z(w454) );
	ym3438_COMP_STR g_1064 (.Z(w455), .A(w1777) );
	ym3438_COMP_STR g_1065 (.Z(w456), .A(w1775) );
	ym3438_COMP_STR g_1066 (.Z(w459), .A(w1773) );
	ym3438_COMP_STR g_1067 (.Z(w460), .A(w1771) );
	ym3438_COMP_STR g_1068 (.Z(w461), .A(w1770) );
	ym3438_COMP_STR g_1069 (.Z(w462), .A(w1768) );
	ym3438_COMP_STR g_1070 (.Z(w458), .A(w1766) );
	ym3438_COMP_STR g_1071 (.Z(w96), .A(w1764) );
	ym3438_COMP_STR g_1072 (.Z(w457), .A(w1762) );
	ym3438_COMP_STR g_1073 (.Z(w69), .A(w1760) );
	ym3438_COMP_STR g_1074 (.Z(w986), .A(w1758) );
	ym3438_COMP_STR g_1075 (.Z(w987), .A(w1756) );
	ym3438_FA g_1076 (.S(w4035), .CI(w386), .A(w403), .B(w1826) );
	ym3438_SR_BIT g_1077 (.Q(w402), .D(w4035), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_COMP_STR g_1078 (.A(w1333), .Z(w886) );
	ym3438_COMP_WE g_1079 (.nZ(w387), .A(w388), .Z(w394) );
	ym3438_COMP_WE g_1080 (.nZ(w393), .A(w389), .Z(w395) );
	ym3438_COMP_WE g_1081 (.nZ(w1862), .A(w1187), .Z(w392) );
	ym3438_NOT g_1082 (.nZ(w396), .A(w1861) );
	ym3438_NOT g_1083 (.nZ(w397), .A(w1860) );
	ym3438_NOT g_1084 (.nZ(w1266), .A(w1859) );
	ym3438_NOT g_1085 (.nZ(w398), .A(w1858) );
	ym3438_NOT g_1086 (.nZ(w399), .A(w1855) );
	ym3438_NOT g_1087 (.nZ(w400), .A(w1856) );
	ym3438_NAND4 g_1088 (.Z(w1855), .B(w395), .A(w394), .C(w392), .D(w391) );
	ym3438_NAND4 g_1089 (.Z(w1856), .B(w395), .A(w387), .C(w392), .D(w391) );
	ym3438_NAND4 g_1090 (.Z(w1857), .B(w393), .A(w394), .C(w392), .D(w391) );
	ym3438_NAND4 g_1091 (.Z(w1858), .B(w393), .A(w387), .C(w392), .D(w391) );
	ym3438_NOT g_1092 (.nZ(w463), .A(w1857) );
	ym3438_NOT g_1093 (.nZ(w391), .A(w390) );
	ym3438_NAND4 g_1094 (.Z(w1861), .B(w393), .A(w394), .C(w1862), .D(w391) );
	ym3438_NAND4 g_1095 (.Z(w1860), .B(w395), .A(w387), .C(w1862), .D(w391) );
	ym3438_NAND4 g_1096 (.Z(w1859), .B(w395), .A(w394), .C(w1862), .D(w391) );
	ym3438_AON22222222 g_1097 (.A1(w399), .Z(w1259), .B2(w417), .A2(w416), .B1(w400), .C1(w463), .C2(w418), .D1(w398), .D2(w419), .E1(w1266), .E2(w420), .F1(w397), .F2(w1261), .G1(w396), .G2(w1260), .H1(w390), .H2(w1249) );
	ym3438_AON22222222 g_1098 (.A1(w399), .Z(w1871), .B2(w419), .A2(w418), .B1(w400), .C1(w463), .C2(w420), .D1(w398), .D2(w1261), .E1(w1266), .E2(w1260), .F1(w397), .F2(w1264), .G1(w396), .G2(w453), .H1(w390), .H2(w416) );
	ym3438_AON22222222 g_1099 (.A1(w399), .Z(w1870), .B2(w1261), .A2(w420), .B1(w400), .C1(w463), .C2(w1260), .D1(w398), .D2(w1264), .E1(w1266), .E2(w453), .F1(w397), .F2(w1332), .G1(w396), .G2(w401), .H1(w390), .H2(w418) );
	ym3438_AOI2222 g_1100 (.A1(w399), .Z(w4426), .B2(w1332), .A2(w453), .B1(w400), .C1(w463), .C2(w401), .D1(w390), .D2(w1260) );
	ym3438_AOI22 g_1101 (.A1(w397), .Z(w1262), .B2(w1265), .A2(w1265), .B1(w396) );
	ym3438_AOI2222 g_1102 (.A1(w398), .Z(w1863), .B2(w1265), .A2(w1265), .B1(w1266), .C1(w397), .C2(w1265), .D1(w396), .D2(w1265) );
	ym3438_AOI222222 g_1103 (.A1(w420), .Z(w233), .B2(w1266), .A2(w390), .B1(w401), .C1(w1332), .C2(w398), .D1(w453), .D2(w463), .E1(w1264), .E2(w400), .F1(w1260), .F2(w399) );
	ym3438_NAND g_1104 (.A(w233), .Z(w1867), .B(w1262) );
	ym3438_AON22222222 g_1108 (.A1(w399), .Z(w1872), .B2(w418), .A2(w417), .B1(w400), .C1(w463), .C2(w419), .D1(w398), .D2(w420), .E1(w1266), .E2(w1261), .F1(w397), .F2(w1260), .G1(w396), .G2(w1264), .H1(w390), .H2(w415) );
	ym3438_AON22222222 g_1109 (.A1(w399), .Z(w1873), .B2(w420), .A2(w419), .B1(w400), .C1(w463), .C2(w1261), .D1(w398), .D2(w1260), .E1(w1266), .E2(w1264), .F1(w397), .F2(w453), .G1(w396), .G2(w1332), .H1(w390), .H2(w417) );
	ym3438_AON22222222 g_1110 (.A1(w399), .Z(w1869), .B2(w1260), .A2(w1261), .B1(w400), .C1(w463), .C2(w1264), .D1(w398), .D2(w453), .E1(w1266), .E2(w1332), .F1(w397), .F2(w401), .G1(w396), .G2(w1265), .H1(w390), .H2(w419) );
	ym3438_NAND g_1111 (.A(w1262), .Z(w1868), .B(w1263) );
	ym3438_AOI222222 g_1112 (.A1(w1261), .Z(w1263), .B2(w1266), .A2(w390), .B1(w1265), .C1(w401), .C2(w398), .D1(w1332), .D2(w463), .E1(w453), .E2(w400), .F1(w1264), .F2(w399) );
	ym3438_NAND g_1113 (.A(w1863), .Z(w1866), .B(w1864) );
	ym3438_AOI2222 g_1114 (.A1(w399), .Z(w1864), .B2(w401), .A2(w1332), .B1(w400), .C1(w463), .C2(w1265), .D1(w390), .D2(w1264) );
	ym3438_SR_BIT g_1132 (.Q(w1874), .D(w1259), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1133 (.Q(w1876), .D(w1872), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1134 (.Q(w1875), .D(w1871), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1135 (.Q(w1877), .D(w1873), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1136 (.Q(w1878), .D(w1870), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1137 (.Q(w4090), .D(w1869), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1138 (.Q(w1880), .D(w1867), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1139 (.Q(w4089), .D(w1868), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1140 (.Q(w1879), .D(w1865), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1141 (.Q(w4088), .D(w1866), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_COMP_STR g_1142 (.A(w402), .Z(w1265) );
	ym3438_SDELAY5 g_1143 (.A(w4088), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .Q(w1256) );
	ym3438_SDELAY5 g_1144 (.A(w4089), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .Q(w1257) );
	ym3438_SDELAY5 g_1145 (.A(w4090), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .Q(w1255) );
	ym3438_SDELAY5 g_1146 (.A(w1877), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .Q(w1254) );
	ym3438_SDELAY5 g_1147 (.A(w1876), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3), .Q(w1251) );
	ym3438_SDELAY5 g_1148 (.A(w1874), .Q(w1250), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3) );
	ym3438_SDELAY5 g_1149 (.A(w1875), .Q(w1252), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3) );
	ym3438_SDELAY5 g_1150 (.A(w1878), .Q(w1253), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3) );
	ym3438_SDELAY5 g_1151 (.A(w1880), .Q(w1258), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3) );
	ym3438_SDELAY5 g_1152 (.A(w1879), .Q(w1267), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3), .C3(w6), .C4(w5), .C5(w6), .C6(w5), .C7(w6), .C8(w5), .C9(w6), .C10(w5), .nC3(w4), .nC4(w3), .nC5(w4), .nC6(w3), .nC7(w4), .nC8(w3), .nC9(w4), .nC10(w3) );
	ym3438_NOT g_1153 (.A(w1319), .nZ(w3) );
	ym3438_NOT g_1154 (.A(w1320), .nZ(w4) );
	ym3438_NOT g_1155 (.A(w1321), .nZ(w6) );
	ym3438_NOT g_1156 (.A(w1322), .nZ(w5) );
	ym3438_NOT g_1157 (.A(w217), .nZ(w1319) );
	ym3438_NOT g_1158 (.A(w212), .nZ(w1320) );
	ym3438_NOT g_1159 (.A(w213), .nZ(w1321) );
	ym3438_NOT g_1160 (.A(w216), .nZ(w1322) );
	ym3438_EXPONENT_TABLE g_1161 (.D12(w1894), .D11(w1895), .D10(w1896), .D9(w1897), .D8(w1898), .D7(w1899), .D6(w1900), .D5(w1901), .D4(w1902), .D3(w1903), .D2(w1892), .D1(w1893), .D0(w1891), .CA3(w473), .CA2(w472), .CA1(w471), .CA0(w468), .RA1(w1905), .RA0(w1904), .RA3(w1298), .RA2(w1906), .RA4(w1907) );
	ym3438_SINE_TABLE g_1162 (.D10(w490), .D9(w479), .D8(w480), .D11(w489), .D3(w1943), .D2(w1944), .D1(w1945), .D0(w1946), .D7(w4391), .D6(w1942), .D5(w4393), .D4(w4392), .D12(w488), .D13(w487), .D14(w486), .D15(w485), .D16(w484), .D17(w483), .D18(w482), .CA3(w1296), .CA2(w1292), .CA1(w1293), .CA0(w1947), .RA1(w1291), .RA0(w1286), .RA3(w1289), .RA2(w1290), .RA4(w1285) );
	ym3438_HA g_1163 (.S(w1199), .A(w1882), .B(w1881) );
	ym3438_HA g_1164 (.CO(w1882), .S(w1200), .A(w1883), .B(w1238) );
	ym3438_HA g_1165 (.CO(w1883), .S(w1201), .A(w1884), .B(w1239) );
	ym3438_HA g_1166 (.CO(w1884), .S(w1202), .A(w1885), .B(w1245) );
	ym3438_HA g_1167 (.CO(w1885), .S(w1203), .A(w1886), .B(w1244) );
	ym3438_HA g_1168 (.CO(w1886), .S(w1204), .A(w1887), .B(w1240) );
	ym3438_HA g_1169 (.CO(w1887), .S(w1205), .A(w1888), .B(w1237) );
	ym3438_FA g_1170 (.CO(w1888), .S(w1206), .CI(w1236), .A(w1247), .B(w1248) );
	ym3438_SR_BITi g_1171 (.nQ(w1881), .D(w1894), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1172 (.nQ(w1238), .D(w1895), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1173 (.nQ(w1239), .D(w1896), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1174 (.nQ(w1245), .D(w1897), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1175 (.nQ(w1244), .D(w1898), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1176 (.nQ(w1240), .D(w1899), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1177 (.nQ(w1237), .D(w1900), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1178 (.nQ(w1246), .D(w1901), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1179 (.nQ(w1247), .D(w1902), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1180 (.nQ(w1242), .D(w1903), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1181 (.nQ(w1241), .D(w1892), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1182 (.nQ(w1243), .D(w1893), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1183 (.nQ(w470), .D(w1891), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_AND g_1184 (.A(w1246), .Z(w1248), .B(w474) );
	ym3438_AND g_1185 (.A(w1243), .Z(w469), .B(w474) );
	ym3438_AND g_1186 (.A(w1242), .Z(w475), .B(w474) );
	ym3438_FA g_1187 (.CO(w1236), .S(w467), .A(w1241), .B(w475), .CI(w4445) );
	ym3438_FA g_1188 (.CI(1'b0), .CO(w4445), .S(w466), .A(w470), .B(w469) );
	ym3438_SR_BIT g_1189 (.Q(w474), .D(w1299), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_NOT g_1190 (.A(w1890), .nZ(w476) );
	ym3438_NOR g_1191 (.A(w476), .Z(w473), .B(w477) );
	ym3438_NOR g_1192 (.A(w1890), .Z(w472), .B(w477) );
	ym3438_NOT g_1193 (.A(w478), .nZ(w477) );
	ym3438_NOR g_1194 (.A(w476), .Z(w471), .B(w478) );
	ym3438_NOR g_1195 (.A(w1890), .Z(w468), .B(w478) );
	ym3438_SR_BIT g_1196 (.Q(w1909), .D(w1908), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1197 (.Q(w1910), .D(w1300), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1198 (.Q(w464), .D(w1911), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1199 (.Q(w1912), .D(w4389), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1200 (.Q(w465), .D(w1913), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1201 (.Q(w1914), .D(w4387), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1202 (.Q(w1208), .D(w1915), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1203 (.Q(w1916), .D(w4388), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1204 (.Q(w1917), .D(w4390), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1205 (.Q(w1207), .D(w1297), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_COMP_STR g_1206 (.A(w1909), .Z(w14) );
	ym3438_NOR g_1207 (.A(w14), .Z(w1911), .B(w1910) );
	ym3438_NOR g_1208 (.A(w14), .Z(w1913), .B(w1912) );
	ym3438_NOR g_1209 (.A(w14), .Z(w1915), .B(w1914) );
	ym3438_NOR g_1210 (.A(w14), .Z(w1297), .B(w1916) );
	ym3438_NOR g_1211 (.A(w14), .Z(w478), .B(w1917) );
	ym3438_NOR g_1212 (.A(w14), .Z(w1907), .B(w15) );
	ym3438_NOR g_1213 (.A(w14), .Z(w1890), .B(w538) );
	ym3438_FA g_1214 (.CO(w1908), .S(w1300), .CI(w1918), .A(w506), .B(w539) );
	ym3438_FA g_1215 (.CO(w1918), .S(w4389), .CI(w1919), .A(w537), .B(w541) );
	ym3438_FA g_1216 (.CO(w1919), .S(w4387), .CI(w1920), .A(w509), .B(w4442) );
	ym3438_FA g_1217 (.CO(w1920), .S(w4388), .CI(w1921), .A(w544), .B(w1922) );
	ym3438_FA g_1218 (.CO(w1921), .S(w4390), .CI(w536), .A(w543), .B(w1923) );
	ym3438_NOR g_1219 (.A(w14), .Z(w1904), .B(w1924) );
	ym3438_NOR g_1220 (.A(w14), .Z(w1905), .B(w1925) );
	ym3438_NOR g_1221 (.A(w14), .Z(w1906), .B(w1926) );
	ym3438_NOR g_1222 (.A(w14), .Z(w1298), .B(w1927) );
	ym3438_NOR g_1223 (.A(w14), .Z(w1299), .B(w542) );
	ym3438_SR_BIT g_1224 (.Q(w538), .D(w4074), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1225 (.Q(w4073), .D(w533), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1226 (.Q(w539), .D(w540), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1227 (.Q(w15), .D(w4071), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1228 (.Q(w4072), .D(w481), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1229 (.Q(w541), .D(w698), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1230 (.Q(w4442), .D(w674), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1231 (.Q(w534), .D(w535), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1232 (.Q(w1922), .D(w669), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1233 (.Q(w1928), .D(w555), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1234 (.Q(w1923), .D(w634), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1235 (.Q(w4441), .D(w551), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1236 (.Q(w1924), .D(w520), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1237 (.Q(w542), .D(w521), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_FA g_1238 (.CO(w536), .S(w4074), .CI(w1929), .A(w505), .B(w4073) );
	ym3438_FA g_1239 (.CO(w1929), .S(w4071), .CI(w1930), .A(w1933), .B(w4072) );
	ym3438_FA g_1240 (.CO(w1930), .S(w529), .CI(w1931), .A(w530), .B(w534) );
	ym3438_FA g_1241 (.CO(w1931), .S(w527), .CI(w1932), .A(w531), .B(w1928) );
	ym3438_FA g_1242 (.CO(w1932), .S(w528), .CI(1'b0), .A(w532), .B(w4441) );
	ym3438_SR_BIT g_1243 (.Q(w1925), .D(w528), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BIT g_1244 (.Q(w1926), .D(w527), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BIT g_1245 (.Q(w1927), .D(w529), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1246 (.nQ(w1934), .D(w482), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1247 (.nQ(w504), .D(w483), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1248 (.nQ(w16), .D(w484), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1249 (.nQ(w507), .D(w485), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1250 (.nQ(w510), .D(w486), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1251 (.nQ(w496), .D(w490), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1252 (.nQ(w497), .D(w489), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1253 (.nQ(w502), .D(w488), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1254 (.nQ(w503), .D(w487), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_HA g_1255 (.CO(w506), .S(w537), .A(w1935), .B(w1934) );
	ym3438_HA g_1256 (.CO(w1935), .S(w509), .A(w1936), .B(w504) );
	ym3438_FA g_1257 (.CO(w1936), .S(w544), .CI(w508), .A(w16), .B(w512) );
	ym3438_FA g_1258 (.CO(w1938), .S(w505), .CI(w515), .A(w503), .B(w511) );
	ym3438_FA g_1259 (.CO(w508), .S(w543), .CI(w1938), .A(w507), .B(w512) );
	ym3438_AND g_1260 (.Z(w512), .B(w510), .A(w523) );
	ym3438_AND g_1261 (.Z(w511), .B(w502), .A(w523) );
	ym3438_FA g_1262 (.CO(w515), .S(w1933), .CI(w1939), .A(w497), .B(w513) );
	ym3438_FA g_1263 (.CO(w1939), .S(w530), .CI(w517), .A(w491), .B(w514) );
	ym3438_AND g_1264 (.Z(w513), .B(w496), .A(w523) );
	ym3438_AND g_1265 (.Z(w514), .B(w498), .A(w523) );
	ym3438_AND g_1266 (.Z(w516), .B(w492), .A(w523) );
	ym3438_AND g_1267 (.Z(w518), .B(w499), .A(w523) );
	ym3438_FA g_1268 (.CO(w1940), .S(w532), .CI(w519), .A(w501), .B(w516) );
	ym3438_FA g_1269 (.CO(w517), .S(w531), .CI(w1940), .A(w495), .B(w518) );
	ym3438_FA g_1270 (.CO(w519), .S(w520), .CI(w1941), .A(w500), .B(w522) );
	ym3438_FA g_1271 (.CO(w1941), .S(w521), .CI(1'b0), .A(w494), .B(w524) );
	ym3438_AND g_1272 (.Z(w522), .B(w493), .A(w523) );
	ym3438_AND g_1273 (.Z(w524), .B(w1937), .A(w523) );
	ym3438_not g_1274 (.nZ(w523), .A(w4075) );
	ym3438_SR_BIT g_1275 (.Q(w4075), .D(w526), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BITi g_1276 (.nQ(w1937), .D(w1946), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1277 (.nQ(w494), .D(w1945), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1278 (.nQ(w493), .D(w1944), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1279 (.nQ(w500), .D(w1943), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1280 (.nQ(w492), .D(w4392), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1281 (.nQ(w501), .D(w4393), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1282 (.nQ(w499), .D(w1942), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1283 (.nQ(w495), .D(w4391), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1284 (.nQ(w498), .D(w480), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_SR_BITi g_1285 (.nQ(w491), .D(w479), .nC1(w4), .nC2(w3), .C1(w6), .C2(w5) );
	ym3438_NOR g_1286 (.Z(w1947), .B(w1294), .A(w1295) );
	ym3438_NOR g_1287 (.Z(w1293), .B(w1294), .A(w1287) );
	ym3438_NOR g_1288 (.Z(w1292), .B(w1288), .A(w1295) );
	ym3438_NOR g_1289 (.Z(w1296), .B(w1288), .A(w1287) );
	ym3438_NOT g_1290 (.nZ(w1295), .A(w1287) );
	ym3438_NOT g_1291 (.nZ(w1294), .A(w1288) );
	ym3438_SR_BIT g_1292 (.Q(w10), .D(w1278), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1293 (.Q(w1284), .D(w1279), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_XOR g_1294 (.A(w1948), .Z(w1288), .B(w1284) );
	ym3438_SR_BIT g_1295 (.Q(w1948), .D(w1280), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_XOR g_1296 (.A(w1951), .Z(w1287), .B(w1284) );
	ym3438_SR_BIT g_1297 (.Q(w1951), .D(w1281), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_XOR g_1298 (.A(w1959), .Z(w1285), .B(w1284) );
	ym3438_XOR g_1299 (.A(w1960), .Z(w1289), .B(w1284) );
	ym3438_XOR g_1300 (.A(w1961), .Z(w1290), .B(w1284) );
	ym3438_XOR g_1301 (.A(w1962), .Z(w1291), .B(w1284) );
	ym3438_XOR g_1302 (.A(w1284), .Z(w1286), .B(w1283) );
	ym3438_XOR g_1303 (.A(w1284), .Z(w526), .B(w1282) );
	ym3438_SR_BIT g_1304 (.Q(w1282), .D(w1272), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1305 (.Q(w1283), .D(w1271), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1306 (.Q(w1962), .D(w1269), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1307 (.Q(w1961), .D(w1268), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1308 (.Q(w1960), .D(w1273), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_SR_BIT g_1309 (.Q(w1959), .D(w1274), .C1(w6), .C2(w5), .nC1(w4), .nC2(w3) );
	ym3438_FA g_1310 (.CO(w1952), .S(w1281), .CI(w1275), .A(w1270), .B(w1258) );
	ym3438_FA g_1311 (.CO(w1950), .S(w1280), .CI(w1952), .A(w1276), .B(w1257) );
	ym3438_FA g_1312 (.CO(w1949), .S(w1279), .CI(w1950), .A(w1324), .B(w1267) );
	ym3438_FA g_1313 (.S(w1278), .CI(w1949), .A(w1277), .B(w1256) );
	ym3438_FA g_1314 (.CO(w1275), .S(w1274), .CI(w1958), .A(w1323), .B(w1255) );
	ym3438_FA g_1315 (.CO(w1958), .S(w1273), .CI(w1957), .A(w1188), .B(w1253) );
	ym3438_FA g_1316 (.CO(w1957), .S(w1268), .CI(w1956), .A(w1189), .B(w1254) );
	ym3438_FA g_1317 (.CO(w1956), .S(w1269), .CI(w1955), .A(w1190), .B(w1252) );
	ym3438_FA g_1318 (.CO(w1955), .S(w1271), .CI(w1954), .A(w1191), .B(w1251) );
	ym3438_FA g_1319 (.CO(w1954), .S(w1272), .CI(1'b0), .A(w1192), .B(w1250) );
	ym3438_DLATCH_INV g_1320 (.nQ(w574), .D(w1335), .C(w17), .nC(w248) );
	ym3438_AOI21 g_1321 (.Z(w2024), .A2(w1980), .A1(w2072), .B(w733) );
	ym3438_NOT g_1322 (.A(w2024), .nZ(w589) );
	ym3438_DLATCH_INV g_1323 (.D(w589), .C(w17), .nC(w248), .nQ(w2025) );
	ym3438_FA g_1324 (.CI(1'b1), .CO(w2026), .S(w575), .A(w2025), .B(w574) );
	ym3438_DLATCH_INV g_1325 (.D(w575), .C(w18), .nC(w545), .nQ(w2029) );
	ym3438_SDELAY23 g_1326 (.A(w2029), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545), .C3(w17), .C4(w18), .C5(w17), .C6(w18), .C7(w17), .C8(w18), .C9(w17), .C10(w18), .C11(w17), .C12(w18), .C13(w17), .C14(w18), .C15(w17), .C16(w18), .C17(w17), .C18(w18), .C19(w17), .C20(w18), .C21(w17), .C22(w18), .C23(w17), .C24(w18), .nC3(w248), .nC4(w545), .nC5(w248), .nC6(w545), .nC7(w248), .nC8(w545), .nC9(w248), .nC10(w545), .nC11(w248), .nC12(w545), .nC13(w248), .nC14(w545), .nC15(w248), .nC16(w545), .nC17(w248), .nC18(w545), .nC19(w248), .nC20(w545), .nC21(w248), .nC22(w545), .nC23(w248), .nC24(w545), .Q(w19), .C25(w17), .C26(w18), .C27(w17), .C28(w18), .C29(w17), .C30(w18), .nC25(w248), .nC26(w545), .nC27(w248), .nC28(w545), .nC29(w248), .nC30(w545), .C36(w18), .nC36(w545), .C35(w17), .nC35(w248), .C34(w18), .nC34(w545), .C33(w17), .nC33(w248), .C32(w18), .nC32(w545), .C31(w17), .nC31(w248), .C42(w18), .nC42(w545), .C41(w17), .nC41(w248), .C40(w18), .nC40(w545), .C39(w17), .nC39(w248), .C38(w18), .nC38(w545), .C37(w17), .nC37(w248), .C44(w18), .nC44(w545), .C43(w17), .nC43(w248), .C46(w18), .nC46(w545), .C45(w17), .nC45(w248), .Q42(w572) );
	ym3438_AON22 g_1327 (.A1(w20), .Z(w1980), .B2(w19), .A2(w731), .B1(w732) );
	ym3438_SR_BIT g_1328 (.Q(w568), .D(w572), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_DLATCH_INV g_1329 (.D(w572), .C(w17), .nC(w248), .nQ(w570) );
	ym3438_HA g_1330 (.CO(w2044), .S(w566), .A(1'b1), .B(w570) );
	ym3438_DLATCH_INV g_1331 (.D(w566), .C(w18), .nC(w545), .nQ(w2030) );
	ym3438_AON22 g_1332 (.A1(w568), .Z(w564), .B2(w2030), .A2(w2042), .B1(w2043) );
	ym3438_SR_BIT g_1333 (.Q(w20), .D(w564), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_AND g_1334 (.Z(w559), .B(w564), .A(w2031) );
	ym3438_AOI2222 g_1335 (.A1(w548), .Z(w561), .A2(w581), .B1(1'b0), .C1(w546), .D2(1'b0), .C2(w580), .D1(w610), .B2(w547) );
	ym3438_DLATCH_INV g_1336 (.nQ(w576), .D(w302), .C(w17), .nC(w248) );
	ym3438_AOI21 g_1337 (.Z(w2046), .A2(w303), .A1(w2072), .B(w733) );
	ym3438_NOT g_1338 (.A(w2046), .nZ(w590) );
	ym3438_DLATCH_INV g_1339 (.nQ(w2028), .D(w590), .C(w17), .nC(w248) );
	ym3438_FA g_1340 (.CI(w2026), .CO(w2049), .S(w2027), .A(w2028), .B(w576) );
	ym3438_DLATCH_INV g_1341 (.nQ(w2045), .D(w2027), .C(w18), .nC(w545) );
	ym3438_SDELAY23 g_1342 (.A(w2045), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545), .C3(w17), .C4(w18), .C5(w17), .C6(w18), .C7(w17), .C8(w18), .C9(w17), .C10(w18), .C11(w17), .C12(w18), .C13(w17), .C14(w18), .C15(w17), .C16(w18), .C17(w17), .C18(w18), .C19(w17), .C20(w18), .C21(w17), .C22(w18), .C23(w17), .C24(w18), .nC3(w248), .nC4(w545), .nC5(w248), .nC6(w545), .nC7(w248), .nC8(w545), .nC9(w248), .nC10(w545), .nC11(w248), .nC12(w545), .nC13(w248), .nC14(w545), .nC15(w248), .nC16(w545), .nC17(w248), .nC18(w545), .nC19(w248), .nC20(w545), .nC21(w248), .nC22(w545), .nC23(w248), .nC24(w545), .Q(w2050), .C25(w17), .C26(w18), .C27(w17), .C28(w18), .C29(w17), .C30(w18), .nC25(w248), .nC26(w545), .nC27(w248), .nC28(w545), .nC29(w248), .nC30(w545), .C36(w18), .nC36(w545), .C35(w17), .nC35(w248), .C34(w18), .nC34(w545), .C33(w17), .nC33(w248), .C32(w18), .nC32(w545), .C31(w17), .nC31(w248), .C42(w18), .nC42(w545), .C41(w17), .nC41(w248), .C40(w18), .nC40(w545), .C39(w17), .nC39(w248), .C38(w18), .nC38(w545), .C37(w17), .nC37(w248), .C44(w18), .nC44(w545), .C43(w17), .nC43(w248), .C46(w18), .nC46(w545), .C45(w17), .nC45(w248), .Q42(w573) );
	ym3438_AON22 g_1343 (.A1(w577), .Z(w303), .B2(w2050), .A2(w731), .B1(w732) );
	ym3438_SR_BIT g_1344 (.Q(w569), .D(w573), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_DLATCH_INV g_1345 (.D(w573), .nC(w248), .C(w17), .nQ(w571) );
	ym3438_HA g_1346 (.CO(w2052), .S(w567), .A(w2044), .B(w571) );
	ym3438_DLATCH_INV g_1347 (.D(w567), .nC(w545), .C(w18), .nQ(w2053) );
	ym3438_AON22 g_1348 (.A1(w569), .Z(w565), .B2(w2053), .A2(w2042), .B1(w2043) );
	ym3438_SR_BIT g_1349 (.Q(w577), .D(w565), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_AND g_1350 (.Z(w560), .B(w565), .A(w2031) );
	ym3438_AOI2222 g_1351 (.A1(w2055), .Z(w562), .B2(w548), .A2(w581), .B1(1'b0), .C1(w547), .D2(w546), .C2(w580), .D1(w610) );
	ym3438_DLATCH_INV g_1352 (.nQ(w591), .D(w1979), .C(w17), .nC(w248) );
	ym3438_AOI21 g_1353 (.Z(w2047), .A2(w305), .A1(w2072), .B(w733) );
	ym3438_NOT g_1354 (.A(w2047), .nZ(w2048) );
	ym3438_DLATCH_INV g_1355 (.D(w2048), .C(w17), .nC(w248), .nQ(w2073) );
	ym3438_FA g_1356 (.CI(w2049), .CO(w2075), .S(w592), .A(w2073), .B(w591) );
	ym3438_DLATCH_INV g_1357 (.D(w592), .C(w18), .nC(w545), .nQ(w2076) );
	ym3438_SDELAY23 g_1358 (.A(w2076), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545), .C3(w17), .C4(w18), .C5(w17), .C6(w18), .C7(w17), .C8(w18), .C9(w17), .C10(w18), .C11(w17), .C12(w18), .C13(w17), .C14(w18), .C15(w17), .C16(w18), .C17(w17), .C18(w18), .C19(w17), .C20(w18), .C21(w17), .C22(w18), .C23(w17), .C24(w18), .nC3(w248), .nC4(w545), .nC5(w248), .nC6(w545), .nC7(w248), .nC8(w545), .nC9(w248), .nC10(w545), .nC11(w248), .nC12(w545), .nC13(w248), .nC14(w545), .nC15(w248), .nC16(w545), .nC17(w248), .nC18(w545), .nC19(w248), .nC20(w545), .nC21(w248), .nC22(w545), .nC23(w248), .nC24(w545), .Q(w2051), .C25(w17), .C26(w18), .C27(w17), .C28(w18), .C29(w17), .C30(w18), .nC25(w248), .nC26(w545), .nC27(w248), .nC28(w545), .nC29(w248), .nC30(w545), .C36(w18), .nC36(w545), .C35(w17), .nC35(w248), .C34(w18), .nC34(w545), .C33(w17), .nC33(w248), .C32(w18), .nC32(w545), .C31(w17), .nC31(w248), .C42(w18), .nC42(w545), .C41(w17), .nC41(w248), .C40(w18), .nC40(w545), .C39(w17), .nC39(w248), .C38(w18), .nC38(w545), .C37(w17), .nC37(w248), .C44(w18), .nC44(w545), .C43(w17), .nC43(w248), .C46(w18), .nC46(w545), .C45(w17), .nC45(w248), .Q42(w595) );
	ym3438_AON22 g_1359 (.A1(w578), .Z(w305), .B2(w2051), .A2(w731), .B1(w732) );
	ym3438_SR_BIT g_1360 (.Q(w596), .D(w595), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_DLATCH_INV g_1361 (.D(w595), .C(w17), .nC(w248), .nQ(w599) );
	ym3438_HA g_1362 (.CO(w2066), .S(w597), .A(w2052), .B(w599) );
	ym3438_DLATCH_INV g_1363 (.D(w597), .C(w18), .nC(w545), .nQ(w2054) );
	ym3438_AON22 g_1364 (.A1(w596), .Z(w615), .B2(w2054), .A2(w2042), .B1(w2043) );
	ym3438_SR_BIT g_1365 (.Q(w578), .D(w615), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_AND g_1366 (.Z(w608), .B(w615), .A(w2031) );
	ym3438_AOI2222 g_1367 (.A1(w614), .Z(w579), .B2(w2055), .A2(w581), .B1(1'b0), .C1(w548), .D2(w547), .C2(w580), .D1(w610) );
	ym3438_NOT g_1368 (.A(w2081), .nZ(w630) );
	ym3438_DLATCH_INV g_1369 (.nQ(w2074), .D(w630), .C(w17), .nC(w248) );
	ym3438_FA g_1370 (.CI(w2075), .CO(w2083), .S(w594), .A(w2074), .B(w593) );
	ym3438_DLATCH_INV g_1371 (.nQ(w2077), .D(w594), .C(w18), .nC(w545) );
	ym3438_SDELAY23 g_1372 (.A(w2077), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545), .C3(w17), .C4(w18), .C5(w17), .C6(w18), .C7(w17), .C8(w18), .C9(w17), .C10(w18), .C11(w17), .C12(w18), .C13(w17), .C14(w18), .C15(w17), .C16(w18), .C17(w17), .C18(w18), .C19(w17), .C20(w18), .C21(w17), .C22(w18), .C23(w17), .C24(w18), .nC3(w248), .nC4(w545), .nC5(w248), .nC6(w545), .nC7(w248), .nC8(w545), .nC9(w248), .nC10(w545), .nC11(w248), .nC12(w545), .nC13(w248), .nC14(w545), .nC15(w248), .nC16(w545), .nC17(w248), .nC18(w545), .nC19(w248), .nC20(w545), .nC21(w248), .nC22(w545), .nC23(w248), .nC24(w545), .Q(w2112), .C25(w17), .C26(w18), .C27(w17), .C28(w18), .C29(w17), .C30(w18), .nC25(w248), .nC26(w545), .nC27(w248), .nC28(w545), .nC29(w248), .nC30(w545), .C36(w18), .nC36(w545), .C35(w17), .nC35(w248), .C34(w18), .nC34(w545), .C33(w17), .nC33(w248), .C32(w18), .nC32(w545), .C31(w17), .nC31(w248), .C42(w18), .nC42(w545), .C41(w17), .nC41(w248), .C40(w18), .nC40(w545), .C39(w17), .nC39(w248), .C38(w18), .nC38(w545), .C37(w17), .nC37(w248), .C44(w18), .nC44(w545), .C43(w17), .nC43(w248), .C46(w18), .nC46(w545), .C45(w17), .nC45(w248), .Q42(w618) );
	ym3438_AON22 g_1373 (.A1(w627), .Z(w304), .B2(w2112), .A2(w731), .B1(w732) );
	ym3438_SR_BIT g_1374 (.Q(w617), .D(w618), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_DLATCH_INV g_1375 (.D(w618), .nC(w248), .C(w17), .nQ(w600) );
	ym3438_HA g_1376 (.CO(w2118), .S(w598), .A(w2066), .B(w600) );
	ym3438_DLATCH_INV g_1377 (.D(w598), .nC(w545), .C(w18), .nQ(w2119) );
	ym3438_AON22 g_1378 (.A1(w617), .Z(w616), .B2(w2119), .A2(w2042), .B1(w2043) );
	ym3438_SR_BIT g_1379 (.Q(w627), .D(w616), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_AND g_1380 (.Z(w612), .B(w616), .A(w2031) );
	ym3438_AOI2222 g_1381 (.A1(w643), .Z(w613), .B2(w614), .A2(w581), .B1(1'b0), .C1(w2055), .D2(w548), .C2(w580), .D1(w610) );
	ym3438_NOT g_1382 (.A(w303), .nZ(w280) );
	ym3438_NOT g_1383 (.A(w305), .nZ(w283) );
	ym3438_AOI221 g_1384 (.Z(w2081), .B2(w2072), .B1(w304), .A(w733), .C2(w2078), .C1(w2079) );
	ym3438_DLATCH_INV g_1385 (.nQ(w593), .D(w301), .C(w17), .nC(w248) );
	ym3438_NOT g_1386 (.A(w2082), .nZ(w629) );
	ym3438_DLATCH_INV g_1387 (.D(w629), .C(w17), .nQ(w2084), .nC(w248) );
	ym3438_FA g_1388 (.CI(w2083), .CO(w2086), .S(w665), .A(w2084), .B(w664) );
	ym3438_DLATCH_INV g_1389 (.D(w665), .C(w18), .nC(w545), .nQ(w2087) );
	ym3438_SDELAY23 g_1390 (.A(w2087), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545), .C3(w17), .C4(w18), .C5(w17), .C6(w18), .C7(w17), .C8(w18), .C9(w17), .C10(w18), .C11(w17), .C12(w18), .C13(w17), .C14(w18), .C15(w17), .C16(w18), .C17(w17), .C18(w18), .C19(w17), .C20(w18), .C21(w17), .C22(w18), .C23(w17), .C24(w18), .nC3(w248), .nC4(w545), .nC5(w248), .nC6(w545), .nC7(w248), .nC8(w545), .nC9(w248), .nC10(w545), .nC11(w248), .nC12(w545), .nC13(w248), .nC14(w545), .nC15(w248), .nC16(w545), .nC17(w248), .nC18(w545), .nC19(w248), .nC20(w545), .nC21(w248), .nC22(w545), .nC23(w248), .nC24(w545), .Q(w2113), .C25(w17), .C26(w18), .C27(w17), .C28(w18), .C29(w17), .C30(w18), .nC25(w248), .nC26(w545), .nC27(w248), .nC28(w545), .nC29(w248), .nC30(w545), .C36(w18), .nC36(w545), .C35(w17), .nC35(w248), .C34(w18), .nC34(w545), .C33(w17), .nC33(w248), .C32(w18), .nC32(w545), .C31(w17), .nC31(w248), .C42(w18), .nC42(w545), .C41(w17), .nC41(w248), .C40(w18), .nC40(w545), .C39(w17), .nC39(w248), .C38(w18), .nC38(w545), .C37(w17), .nC37(w248), .C44(w18), .nC44(w545), .C43(w17), .nC43(w248), .C46(w18), .nC46(w545), .C45(w17), .nC45(w248), .Q42(w653) );
	ym3438_AON22 g_1391 (.A1(w628), .Z(w306), .B2(w2113), .A2(w731), .B1(w732) );
	ym3438_SR_BIT g_1392 (.Q(w647), .D(w653), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_DLATCH_INV g_1393 (.D(w653), .C(w17), .nC(w248), .nQ(w651) );
	ym3438_HA g_1394 (.CO(w2067), .S(w648), .A(w2118), .B(w651) );
	ym3438_DLATCH_INV g_1395 (.D(w648), .C(w18), .nC(w545), .nQ(w2120) );
	ym3438_AON22 g_1396 (.A1(w647), .Z(w645), .B2(w2120), .A2(w2042), .B1(w2043) );
	ym3438_SR_BIT g_1397 (.Q(w628), .D(w645), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_AND g_1398 (.Z(w640), .B(w645), .A(w2031) );
	ym3438_AOI2222 g_1399 (.A1(1'b0), .Z(w642), .B2(w643), .A2(w581), .B1(1'b0), .C1(w614), .D2(w2055), .C2(w580), .D1(w610) );
	ym3438_AOI221 g_1400 (.Z(w2082), .B2(w2072), .B1(w306), .A(w733), .C2(w2078), .C1(w2080) );
	ym3438_DLATCH_INV g_1401 (.nQ(w664), .D(w308), .C(w17), .nC(w248) );
	ym3438_DLATCH_INV g_1402 (.nQ(w667), .D(w310), .C(w17), .nC(w248) );
	ym3438_NOT g_1403 (.A(w2099), .nZ(w234) );
	ym3438_DLATCH_INV g_1404 (.nQ(w2085), .D(w234), .C(w17), .nC(w248) );
	ym3438_FA g_1405 (.CI(w2086), .CO(w2101), .S(w666), .A(w2085), .B(w667) );
	ym3438_DLATCH_INV g_1406 (.nQ(w2088), .D(w666), .C(w18), .nC(w545) );
	ym3438_SDELAY23 g_1407 (.A(w2088), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545), .C3(w17), .C4(w18), .C5(w17), .C6(w18), .C7(w17), .C8(w18), .C9(w17), .C10(w18), .C11(w17), .C12(w18), .C13(w17), .C14(w18), .C15(w17), .C16(w18), .C17(w17), .C18(w18), .C19(w17), .C20(w18), .C21(w17), .C22(w18), .C23(w17), .C24(w18), .nC3(w248), .nC4(w545), .nC5(w248), .nC6(w545), .nC7(w248), .nC8(w545), .nC9(w248), .nC10(w545), .nC11(w248), .nC12(w545), .nC13(w248), .nC14(w545), .nC15(w248), .nC16(w545), .nC17(w248), .nC18(w545), .nC19(w248), .nC20(w545), .nC21(w248), .nC22(w545), .nC23(w248), .nC24(w545), .Q(w2114), .C25(w17), .C26(w18), .C27(w17), .C28(w18), .C29(w17), .C30(w18), .nC25(w248), .nC26(w545), .nC27(w248), .nC28(w545), .nC29(w248), .nC30(w545), .C36(w18), .nC36(w545), .C35(w17), .nC35(w248), .C34(w18), .nC34(w545), .C33(w17), .nC33(w248), .C32(w18), .nC32(w545), .C31(w17), .nC31(w248), .C42(w18), .nC42(w545), .C41(w17), .nC41(w248), .C40(w18), .nC40(w545), .C39(w17), .nC39(w248), .C38(w18), .nC38(w545), .C37(w17), .nC37(w248), .C44(w18), .nC44(w545), .C43(w17), .nC43(w248), .C46(w18), .nC46(w545), .C45(w17), .nC45(w248), .Q42(w654) );
	ym3438_AON22 g_1408 (.A1(w662), .Z(w309), .B2(w2114), .A2(w731), .B1(w732) );
	ym3438_SR_BIT g_1409 (.Q(w650), .D(w654), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_DLATCH_INV g_1410 (.D(w654), .nC(w248), .C(w17), .nQ(w652) );
	ym3438_HA g_1411 (.CO(w2121), .S(w649), .A(w2067), .B(w652) );
	ym3438_DLATCH_INV g_1412 (.D(w649), .nC(w545), .C(w18), .nQ(w2122) );
	ym3438_AON22 g_1413 (.A1(w650), .Z(w646), .B2(w2122), .A2(w2042), .B1(w2043) );
	ym3438_AOI221 g_1414 (.Z(w2099), .B2(w2072), .B1(w309), .A(w733), .C2(w2078), .C1(w2107) );
	ym3438_SR_BIT g_1415 (.Q(w662), .D(w646), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_AND g_1416 (.Z(w641), .B(w646), .A(w2031) );
	ym3438_AOI22 g_1417 (.A1(w643), .Z(w644), .B2(w614), .A2(w580), .B1(w610) );
	ym3438_DLATCH_INV g_1418 (.nQ(w690), .D(w1337), .C(w17), .nC(w248) );
	ym3438_NOT g_1419 (.A(w2100), .nZ(w235) );
	ym3438_DLATCH_INV g_1420 (.D(w235), .C(w17), .nQ(w2089), .nC(w248) );
	ym3438_FA g_1421 (.CI(w2101), .CO(w2091), .S(w689), .A(w2089), .B(w690) );
	ym3438_DLATCH_INV g_1422 (.D(w689), .C(w18), .nC(w545), .nQ(w2092) );
	ym3438_SDELAY23 g_1423 (.A(w2092), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545), .C3(w17), .C4(w18), .C5(w17), .C6(w18), .C7(w17), .C8(w18), .C9(w17), .C10(w18), .C11(w17), .C12(w18), .C13(w17), .C14(w18), .C15(w17), .C16(w18), .C17(w17), .C18(w18), .C19(w17), .C20(w18), .C21(w17), .C22(w18), .C23(w17), .C24(w18), .nC3(w248), .nC4(w545), .nC5(w248), .nC6(w545), .nC7(w248), .nC8(w545), .nC9(w248), .nC10(w545), .nC11(w248), .nC12(w545), .nC13(w248), .nC14(w545), .nC15(w248), .nC16(w545), .nC17(w248), .nC18(w545), .nC19(w248), .nC20(w545), .nC21(w248), .nC22(w545), .nC23(w248), .nC24(w545), .Q(w2115), .C25(w17), .C26(w18), .C27(w17), .C28(w18), .C29(w17), .C30(w18), .nC25(w248), .nC26(w545), .nC27(w248), .nC28(w545), .nC29(w248), .nC30(w545), .C36(w18), .nC36(w545), .C35(w17), .nC35(w248), .C34(w18), .nC34(w545), .C33(w17), .nC33(w248), .C32(w18), .nC32(w545), .C31(w17), .nC31(w248), .C42(w18), .nC42(w545), .C41(w17), .nC41(w248), .C40(w18), .nC40(w545), .C39(w17), .nC39(w248), .C38(w18), .nC38(w545), .C37(w17), .nC37(w248), .C44(w18), .nC44(w545), .C43(w17), .nC43(w248), .C46(w18), .nC46(w545), .C45(w17), .nC45(w248), .Q42(w687) );
	ym3438_AON22 g_1424 (.A1(w663), .Z(w300), .B2(w2115), .A2(w731), .B1(w732) );
	ym3438_SR_BIT g_1425 (.Q(w682), .D(w687), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_DLATCH_INV g_1426 (.D(w687), .C(w17), .nC(w248), .nQ(w686) );
	ym3438_HA g_1427 (.CO(w2068), .S(w683), .A(w2121), .B(w686) );
	ym3438_DLATCH_INV g_1428 (.D(w683), .C(w18), .nC(w545), .nQ(w2123) );
	ym3438_AON22 g_1429 (.A1(w682), .Z(w2127), .B2(w2123), .A2(w2042), .B1(w2043) );
	ym3438_AOI221 g_1430 (.Z(w2100), .B2(w2072), .B1(w300), .A(w733), .C2(w2078), .C1(w2108) );
	ym3438_SR_BIT g_1431 (.Q(w663), .D(w2127), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_AND g_1432 (.Z(w677), .B(w2127), .A(w2031) );
	ym3438_AOI22 g_1433 (.A1(1'b0), .Z(w679), .B2(w643), .A2(w580), .B1(w610) );
	ym3438_DLATCH_INV g_1434 (.nQ(w691), .D(w313), .C(w17), .nC(w248) );
	ym3438_NOT g_1435 (.A(w2102), .nZ(w704) );
	ym3438_DLATCH_INV g_1436 (.nQ(w2090), .D(w704), .C(w17), .nC(w248) );
	ym3438_FA g_1437 (.CI(w2091), .CO(w2104), .S(w692), .A(w2090), .B(w691) );
	ym3438_DLATCH_INV g_1438 (.nQ(w2093), .D(w692), .C(w18), .nC(w545) );
	ym3438_SDELAY23 g_1439 (.A(w2093), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545), .C3(w17), .C4(w18), .C5(w17), .C6(w18), .C7(w17), .C8(w18), .C9(w17), .C10(w18), .C11(w17), .C12(w18), .C13(w17), .C14(w18), .C15(w17), .C16(w18), .C17(w17), .C18(w18), .C19(w17), .C20(w18), .C21(w17), .C22(w18), .C23(w17), .C24(w18), .nC3(w248), .nC4(w545), .nC5(w248), .nC6(w545), .nC7(w248), .nC8(w545), .nC9(w248), .nC10(w545), .nC11(w248), .nC12(w545), .nC13(w248), .nC14(w545), .nC15(w248), .nC16(w545), .nC17(w248), .nC18(w545), .nC19(w248), .nC20(w545), .nC21(w248), .nC22(w545), .nC23(w248), .nC24(w545), .Q(w2116), .C25(w17), .C26(w18), .C27(w17), .C28(w18), .C29(w17), .C30(w18), .nC25(w248), .nC26(w545), .nC27(w248), .nC28(w545), .nC29(w248), .nC30(w545), .C36(w18), .nC36(w545), .C35(w17), .nC35(w248), .C34(w18), .nC34(w545), .C33(w17), .nC33(w248), .C32(w18), .nC32(w545), .C31(w17), .nC31(w248), .C42(w18), .nC42(w545), .C41(w17), .nC41(w248), .C40(w18), .nC40(w545), .C39(w17), .nC39(w248), .C38(w18), .nC38(w545), .C37(w17), .nC37(w248), .C44(w18), .nC44(w545), .C43(w17), .nC43(w248), .C46(w18), .nC46(w545), .C45(w17), .nC45(w248), .Q42(w688) );
	ym3438_AON22 g_1440 (.A1(w696), .Z(w307), .B2(w2116), .A2(w731), .B1(w732) );
	ym3438_SR_BIT g_1441 (.Q(w2069), .D(w688), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_DLATCH_INV g_1442 (.D(w688), .nC(w248), .C(w17), .nQ(w685) );
	ym3438_HA g_1443 (.CO(w2124), .S(w684), .A(w2068), .B(w685) );
	ym3438_DLATCH_INV g_1444 (.D(w684), .nC(w545), .C(w18), .nQ(w2125) );
	ym3438_AON22 g_1445 (.A1(w2069), .Z(w681), .B2(w2125), .A2(w2042), .B1(w2043) );
	ym3438_AOI221 g_1446 (.Z(w2102), .B2(w2072), .B1(w307), .A(w733), .C2(w2078), .C1(w2109) );
	ym3438_SR_BIT g_1447 (.Q(w696), .D(w681), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_AND g_1448 (.Z(w678), .B(w681), .A(w2031) );
	ym3438_DLATCH_INV g_1449 (.nQ(w722), .D(w272), .C(w17), .nC(w248) );
	ym3438_NOT g_1450 (.A(w2103), .nZ(w705) );
	ym3438_DLATCH_INV g_1451 (.D(w705), .C(w17), .nQ(w2094), .nC(w248) );
	ym3438_FA g_1452 (.CI(w2104), .CO(w2096), .S(w721), .A(w2094), .B(w722) );
	ym3438_DLATCH_INV g_1453 (.D(w721), .C(w18), .nC(w545), .nQ(w2097) );
	ym3438_SDELAY23 g_1454 (.A(w2097), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545), .C3(w17), .C4(w18), .C5(w17), .C6(w18), .C7(w17), .C8(w18), .C9(w17), .C10(w18), .C11(w17), .C12(w18), .C13(w17), .C14(w18), .C15(w17), .C16(w18), .C17(w17), .C18(w18), .C19(w17), .C20(w18), .C21(w17), .C22(w18), .C23(w17), .C24(w18), .nC3(w248), .nC4(w545), .nC5(w248), .nC6(w545), .nC7(w248), .nC8(w545), .nC9(w248), .nC10(w545), .nC11(w248), .nC12(w545), .nC13(w248), .nC14(w545), .nC15(w248), .nC16(w545), .nC17(w248), .nC18(w545), .nC19(w248), .nC20(w545), .nC21(w248), .nC22(w545), .nC23(w248), .nC24(w545), .Q(w2117), .C25(w17), .C26(w18), .C27(w17), .C28(w18), .C29(w17), .C30(w18), .nC25(w248), .nC26(w545), .nC27(w248), .nC28(w545), .nC29(w248), .nC30(w545), .C36(w18), .nC36(w545), .C35(w17), .nC35(w248), .C34(w18), .nC34(w545), .C33(w17), .nC33(w248), .C32(w18), .nC32(w545), .C31(w17), .nC31(w248), .C42(w18), .nC42(w545), .C41(w17), .nC41(w248), .C40(w18), .nC40(w545), .C39(w17), .nC39(w248), .C38(w18), .nC38(w545), .C37(w17), .nC37(w248), .C44(w18), .nC44(w545), .C43(w17), .nC43(w248), .C46(w18), .nC46(w545), .C45(w17), .nC45(w248), .Q42(w720) );
	ym3438_AON22 g_1455 (.A1(w697), .Z(w318), .B2(w2117), .A2(w731), .B1(w732) );
	ym3438_SR_BIT g_1456 (.Q(w718), .D(w720), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_DLATCH_INV g_1457 (.D(w720), .C(w17), .nC(w248), .nQ(w2071) );
	ym3438_HA g_1458 (.CO(w2070), .S(w717), .A(w2124), .B(w2071) );
	ym3438_DLATCH_INV g_1459 (.D(w717), .C(w18), .nC(w545), .nQ(w2126) );
	ym3438_AON22 g_1460 (.A1(w718), .Z(w714), .B2(w2126), .A2(w2042), .B1(w2043) );
	ym3438_AOI221 g_1461 (.Z(w2103), .B2(w2072), .B1(w318), .A(w733), .C2(w2078), .C1(w2110) );
	ym3438_SR_BIT g_1462 (.Q(w697), .D(w714), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_AND g_1463 (.Z(w713), .B(w714), .A(w2031) );
	ym3438_DLATCH_INV g_1464 (.nQ(w734), .D(w236), .C(w17), .nC(w248) );
	ym3438_NOT g_1465 (.A(w2105), .nZ(w2106) );
	ym3438_DLATCH_INV g_1466 (.nQ(w2095), .D(w2106), .C(w17), .nC(w248) );
	ym3438_FA g_1467 (.CI(w2096), .S(w735), .A(w2095), .B(w734) );
	ym3438_DLATCH_INV g_1468 (.nQ(w2098), .D(w735), .nC(w545), .C(w18) );
	ym3438_SDELAY23 g_1469 (.A(w2098), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545), .C3(w17), .C4(w18), .C5(w17), .C6(w18), .C7(w17), .C8(w18), .C9(w17), .C10(w18), .C11(w17), .C12(w18), .C13(w17), .C14(w18), .C15(w17), .C16(w18), .C17(w17), .C18(w18), .C19(w17), .C20(w18), .C21(w17), .C22(w18), .C23(w17), .C24(w18), .nC3(w248), .nC4(w545), .nC5(w248), .nC6(w545), .nC7(w248), .nC8(w545), .nC9(w248), .nC10(w545), .nC11(w248), .nC12(w545), .nC13(w248), .nC14(w545), .nC15(w248), .nC16(w545), .nC17(w248), .nC18(w545), .nC19(w248), .nC20(w545), .nC21(w248), .nC22(w545), .nC23(w248), .nC24(w545), .Q(w2162), .C25(w17), .C26(w18), .C27(w17), .C28(w18), .C29(w17), .C30(w18), .nC25(w248), .nC26(w545), .nC27(w248), .nC28(w545), .nC29(w248), .nC30(w545), .C36(w18), .nC36(w545), .C35(w17), .nC35(w248), .C34(w18), .nC34(w545), .C33(w17), .nC33(w248), .C32(w18), .nC32(w545), .C31(w17), .nC31(w248), .C42(w18), .nC42(w545), .C41(w17), .nC41(w248), .C40(w18), .nC40(w545), .C39(w17), .nC39(w248), .C38(w18), .nC38(w545), .C37(w17), .nC37(w248), .C44(w18), .nC44(w545), .C43(w17), .nC43(w248), .C46(w18), .nC46(w545), .C45(w17), .nC45(w248), .Q42(w2111) );
	ym3438_AON22 g_1470 (.A1(w2163), .Z(w317), .B2(w2162), .A2(w731), .B1(w732) );
	ym3438_SR_BIT g_1471 (.Q(w719), .D(w2111), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_DLATCH_INV g_1472 (.D(w2111), .nC(w248), .C(w17), .nQ(w1305) );
	ym3438_AON22 g_1473 (.A1(w719), .Z(w715), .B2(w4087), .A2(w2042), .B1(w2043) );
	ym3438_AOI221 g_1474 (.Z(w2105), .B2(w2072), .A(w733), .C2(w2078), .C1(w2159), .B1(w317) );
	ym3438_SR_BIT g_1475 (.Q(w2163), .D(w715), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_AND g_1476 (.Z(w729), .B(w715), .A(w2031) );
	ym3438_DLATCH_INV g_1477 (.D(w730), .nC(w545), .C(w18), .nQ(w4086) );
	ym3438_SLATCH g_1478 (.Q(w793), .D(w249), .C(w238), .nC(w237) );
	ym3438_SLATCH g_1479 (.Q(w1325), .D(w1963), .C(w238), .nC(w237) );
	ym3438_SR_BIT g_1480 (.Q(w244), .D(w250), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SR_BIT g_1481 (.Q(w239), .D(w244), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SR_BIT g_1482 (.Q(w247), .D(w239), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SR_BIT g_1483 (.Q(w240), .D(w247), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SR_BIT g_1484 (.Q(w251), .D(w240), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_OR5 g_1485 (.Z(w1964), .B(w239), .A(w244), .C(w247), .D(w240), .E(w251) );
	ym3438_SLATCH g_1486 (.Q(w1326), .D(w1964), .C(w238), .nC(w237) );
	ym3438_SR_BIT g_1487 (.Q(w253), .D(w251), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SR_BIT g_1488 (.Q(w241), .D(w253), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SR_BIT g_1489 (.Q(w242), .D(w241), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SLATCH g_1490 (.Q(w1327), .D(w1965), .C(w238), .nC(w237) );
	ym3438_OR5 g_1491 (.Z(w1965), .B(w253), .A(w244), .C(w241), .D(w242), .E(w245) );
	ym3438_SR_BIT g_1492 (.Q(w245), .D(w242), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SLATCH g_1493 (.Q(w786), .D(w1970), .C(w238), .nC(w237) );
	ym3438_OR6 g_1494 (.Z(w1970), .B(w247), .A(w253), .C(w239), .D(w241), .E(w246), .F(w243) );
	ym3438_SR_BIT g_1495 (.Q(w246), .D(w245), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SR_BIT g_1496 (.Q(w243), .D(w246), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SR_BIT g_1497 (.Q(w1971), .D(w243), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_OR6 g_1498 (.Z(w1972), .B(w240), .A(w253), .C(w239), .D(w242), .E(w246), .F(w1971) );
	ym3438_SLATCH g_1499 (.Q(w1164), .D(w1972), .C(w238), .nC(w237) );
	ym3438_COMP_WE g_1500 (.Z(w238), .A(w1334), .nZ(w237) );
	ym3438_SDELAY12 g_1501 (.A(w255), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545), .C3(w17), .C4(w18), .C5(w17), .C6(w18), .C7(w17), .C8(w18), .C9(w17), .C10(w18), .C11(w17), .C12(w18), .C13(w17), .C14(w18), .C15(w17), .C16(w18), .C17(w17), .C18(w18), .C19(w17), .C20(w18), .C21(w17), .C22(w18), .C23(w17), .C24(w18), .nC3(w248), .nC4(w545), .nC5(w248), .nC6(w545), .nC7(w248), .nC8(w545), .nC9(w248), .nC10(w545), .nC11(w248), .nC12(w545), .nC13(w248), .nC14(w545), .nC15(w248), .nC16(w545), .nC17(w248), .nC18(w545), .nC19(w248), .nC20(w545), .nC21(w248), .nC22(w545), .nC23(w248), .nC24(w545), .Q(w249), .Q22(w1963) );
	ym3438_SR_BIT g_1502 (.Q(w256), .D(w1966), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_HA g_1503 (.CO(w1966), .S(w254), .A(w1967), .B(w249) );
	ym3438_NOT g_1504 (.A(w1968), .nZ(w1967) );
	ym3438_AOI21 g_1505 (.A1(w252), .Z(w1968), .B(w256), .A2(w781) );
	ym3438_NOT g_1506 (.A(w258), .nZ(w257) );
	ym3438_AND g_1507 (.Z(w250), .B(w259), .A(w257) );
	ym3438_OR g_1508 (.Z(w259), .B(w782), .A(w255) );
	ym3438_AND g_1509 (.Z(w255), .B(w1969), .A(w254) );
	ym3438_NOR g_1510 (.Z(w1969), .B(w262), .A(w263) );
	ym3438_OR g_1511 (.Z(w1975), .B(w259), .A(w258) );
	ym3438_SR_BIT g_1512 (.Q(w258), .D(w1976), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_AND g_1513 (.Z(w1976), .B(w1974), .A(w1975) );
	ym3438_NOR3 g_1514 (.Z(w1974), .B(w261), .A(w262), .C(w1973) );
	ym3438_SDELAY12 g_1515 (.A(w261), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545), .C3(w17), .C4(w18), .C5(w17), .C6(w18), .C7(w17), .C8(w18), .C9(w17), .C10(w18), .C11(w17), .C12(w18), .C13(w17), .C14(w18), .C15(w17), .C16(w18), .C17(w17), .C18(w18), .C19(w17), .C20(w18), .C21(w17), .C22(w18), .C23(w17), .C24(w18), .nC3(w248), .nC4(w545), .nC5(w248), .nC6(w545), .nC7(w248), .nC8(w545), .nC9(w248), .nC10(w545), .nC11(w248), .nC12(w545), .nC13(w248), .nC14(w545), .nC15(w248), .nC16(w545), .nC17(w248), .nC18(w545), .nC19(w248), .nC20(w545), .nC21(w248), .nC22(w545), .nC23(w248), .nC24(w545), .Q(w1973) );
	ym3438_SR_BIT g_1516 (.Q(w252), .D(w261), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_AOI33 g_1517 (.A1(w265), .Z(w279), .B2(w264), .A2(w268), .B1(w280), .A3(w266), .B3(w267) );
	ym3438_AOI333 g_1518 (.A1(w268), .Z(w278), .B2(w264), .A2(w264), .B1(w778), .A3(w281), .B3(w269), .C2(w264), .C1(w779), .C3(w283) );
	ym3438_AOI33 g_1519 (.A1(w265), .Z(w1977), .B2(w264), .A2(w778), .B1(w283), .A3(w266), .B3(w267) );
	ym3438_AOI333 g_1520 (.A1(w268), .Z(w282), .B2(w264), .A2(w264), .B1(w778), .A3(w286), .B3(w281), .C2(w264), .C1(w779), .C3(w269) );
	ym3438_AOI333 g_1521 (.A1(w267), .Z(w277), .B2(w779), .A2(w264), .B1(w266), .A3(w269), .B3(w265), .C2(w268), .C1(w270), .C3(w265) );
	ym3438_AOI333 g_1522 (.A1(w268), .Z(w276), .B2(w264), .A2(w264), .B1(w778), .A3(w291), .B3(w286), .C2(w264), .C1(w779), .C3(w281) );
	ym3438_AOI333 g_1523 (.A1(w267), .Z(w288), .B2(w267), .A2(w264), .B1(w266), .A3(w281), .B3(w265), .C2(w778), .C1(w270), .C3(w265) );
	ym3438_AOI333 g_1524 (.A1(w268), .Z(w287), .B2(w264), .A2(w264), .B1(w778), .A3(w290), .B3(w291), .C2(w264), .C1(w779), .C3(w286) );
	ym3438_AOI33 g_1525 (.A1(w265), .Z(w285), .B2(w264), .A2(w779), .B1(w286), .A3(w270), .B3(w267) );
	ym3438_AOI333 g_1526 (.A1(w268), .Z(w284), .B2(w264), .A2(w264), .B1(w778), .A3(w293), .B3(w290), .C2(w264), .C1(w779), .C3(w291) );
	ym3438_AOI33 g_1527 (.A1(w265), .Z(w273), .B2(w264), .A2(w267), .B1(w291), .A3(w270), .B3(w267) );
	ym3438_AOI333 g_1528 (.A1(w268), .Z(w275), .B2(w264), .A2(w264), .B1(w778), .A3(w294), .B3(w293), .C2(w264), .C1(w779), .C3(w290) );
	ym3438_AOI33 g_1529 (.A1(w294), .Z(w260), .B2(w779), .A2(w264), .B1(w264), .A3(w267), .B3(1'b1) );
	ym3438_NAND g_1530 (.Z(w272), .B(w260), .A(w319) );
	ym3438_AON2222 g_1531 (.A1(w268), .Z(w236), .B2(w778), .A2(w264), .B1(w264), .D1(w267), .D2(w264), .C2(w779), .C1(w264) );
	ym3438_AND g_1532 (.Z(w271), .B(w289), .A(w274) );
	ym3438_NAND g_1533 (.Z(w1335), .B(w278), .A(w279) );
	ym3438_NAND g_1534 (.Z(w302), .B(w282), .A(w1977) );
	ym3438_NAND g_1535 (.Z(w1979), .B(w276), .A(w277) );
	ym3438_NOT g_1536 (.A(w304), .nZ(w269) );
	ym3438_NOR5 g_1537 (.Z(w289), .B(w303), .A(w1980), .C(w305), .D(w304), .E(w306) );
	ym3438_NAND g_1538 (.Z(w301), .B(w287), .A(w288) );
	ym3438_NOT g_1539 (.A(w306), .nZ(w281) );
	ym3438_NAND g_1540 (.Z(w308), .B(w284), .A(w285) );
	ym3438_NOT g_1541 (.A(w309), .nZ(w286) );
	ym3438_XOR g_1542 (.Z(w315), .B(w311), .A(w309) );
	ym3438_NOT g_1543 (.A(w300), .nZ(w291) );
	ym3438_NAND g_1544 (.Z(w310), .B(w275), .A(w273) );
	ym3438_XOR g_1545 (.Z(w320), .B(w312), .A(w300) );
	ym3438_NOT g_1546 (.A(w307), .nZ(w290) );
	ym3438_AON3333 g_1547 (.A1(1'b1), .Z(w1337), .B2(w264), .A2(w268), .B1(w778), .A3(w264), .B3(w294), .C1(w779), .D2(w264), .C2(w264), .D1(w267), .C3(w293), .D3(w290) );
	ym3438_XOR g_1548 (.Z(w1981), .B(w295), .A(w307) );
	ym3438_NOR5 g_1549 (.Z(w274), .B(w300), .A(w309), .C(w307), .D(w318), .E(w317) );
	ym3438_AND6 g_1550 (.Z(w299), .B(w309), .A(w300), .C(w306), .D(w317), .E(w307), .F(w318) );
	ym3438_NOR6 g_1551 (.Z(w314), .B(w320), .A(w306), .C(w315), .D(w1981), .E(w292), .F(w297) );
	ym3438_AOI22 g_1552 (.A1(w268), .Z(w319), .B2(w264), .A2(w264), .B1(w778) );
	ym3438_AOI33 g_1553 (.A1(w293), .Z(w298), .B2(w264), .A2(w264), .B1(w294), .A3(w267), .B3(w779) );
	ym3438_NAND g_1554 (.Z(w313), .B(w319), .A(w298) );
	ym3438_XOR g_1555 (.Z(w292), .B(w316), .A(w318) );
	ym3438_XOR g_1556 (.Z(w297), .B(w296), .A(w317) );
	ym3438_NOT g_1557 (.A(w318), .nZ(w293) );
	ym3438_NOT g_1558 (.A(w317), .nZ(w294) );
	ym3438_FA g_1559 (.CO(w2038), .S(w557), .CI(1'b0), .A(w2040), .B(w559) );
	ym3438_FA g_1560 (.CO(w2057), .S(w558), .CI(w2038), .A(w2039), .B(w560) );
	ym3438_FA g_1561 (.CO(w611), .S(w607), .CI(w2057), .A(w2056), .B(w608) );
	ym3438_FA g_1562 (.CO(w2128), .S(w609), .CI(w611), .A(w2065), .B(w612) );
	ym3438_FA g_1563 (.CO(w2134), .S(w638), .CI(w2128), .A(w2135), .B(w640) );
	ym3438_FA g_1564 (.CO(w2138), .S(w639), .CI(w2134), .A(w2136), .B(w641) );
	ym3438_FA g_1565 (.CO(w2143), .S(w675), .CI(w2138), .A(w2144), .B(w677) );
	ym3438_FA g_1566 (.CO(w2147), .S(w676), .CI(w2143), .A(1'b0), .B(w678) );
	ym3438_FA g_1567 (.CO(w2150), .S(w712), .CI(w2147), .A(1'b0), .B(w713) );
	ym3438_FA g_1568 (.CO(w711), .S(w728), .CI(w2150), .A(1'b0), .B(w729) );
	ym3438_FA g_1569 (.CO(w2130), .S(w606), .CI(1'b1), .A(w2064), .B(w622) );
	ym3438_FA g_1570 (.CO(w2131), .S(w637), .CI(w2130), .A(w2132), .B(w621) );
	ym3438_FA g_1571 (.CO(w2139), .S(w636), .CI(w2131), .A(w2133), .B(w656) );
	ym3438_FA g_1572 (.CO(w2140), .S(w671), .CI(w2139), .A(w2141), .B(w657) );
	ym3438_FA g_1573 (.CO(w2146), .S(w672), .CI(w2140), .A(w2142), .B(w695) );
	ym3438_FA g_1574 (.CO(w2151), .S(w708), .CI(w2146), .A(w2152), .B(w701) );
	ym3438_DLATCH_INV g_1575 (.D(w613), .nC(w545), .C(w18), .nQ(w2065) );
	ym3438_DLATCH_INV g_1576 (.D(w642), .C(w18), .nC(w545), .nQ(w2135) );
	ym3438_DLATCH_INV g_1577 (.D(w644), .nC(w545), .C(w18), .nQ(w2136) );
	ym3438_DLATCH_INV g_1578 (.D(w679), .C(w18), .nC(w545), .nQ(w2144) );
	ym3438_DLATCH_INV g_1579 (.D(w1196), .nC(w248), .C(w17), .nQ(w2145) );
	ym3438_DLATCH_INV g_1580 (.D(w711), .nC(w248), .C(w17), .nQ(w2148) );
	ym3438_NOT g_1581 (.nZ(w700), .A(w2149) );
	ym3438_SR_BIT g_1582 (.Q(w2078), .D(w4463), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_NAND g_1583 (.Z(w2149), .B(w710), .A(w2148) );
	ym3438_SR_BIT g_1584 (.Q(w4463), .D(w1186), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_NOT g_1585 (.nZ(w643), .A(w2145) );
	ym3438_AND g_1586 (.Z(w580), .B(w588), .A(w583) );
	ym3438_AND g_1587 (.Z(w581), .B(w2041), .A(w582) );
	ym3438_AND g_1588 (.Z(w610), .B(w583), .A(w582) );
	ym3438_DLATCH_INV g_1589 (.D(w579), .C(w18), .nC(w545), .nQ(w2056) );
	ym3438_DLATCH_INV g_1590 (.D(w562), .nC(w545), .C(w18), .nQ(w2039) );
	ym3438_DLATCH_INV g_1591 (.D(w561), .C(w18), .nC(w545), .nQ(w2040) );
	ym3438_DLATCH_INV g_1592 (.D(w549), .C(w17), .nC(w248), .nQ(w2033) );
	ym3438_DLATCH_INV g_1593 (.D(w1198), .C(w17), .nC(w248), .nQ(w2032) );
	ym3438_NOT g_1594 (.nZ(w546), .A(w2032) );
	ym3438_NOT g_1595 (.nZ(w547), .A(w2033) );
	ym3438_NOT g_1596 (.nZ(w588), .A(w582) );
	ym3438_NOT g_1597 (.nZ(w2041), .A(w583) );
	ym3438_AND g_1598 (.B(w2041), .A(w588) );
	ym3438_NOT g_1599 (.nZ(w548), .A(w2034) );
	ym3438_DLATCH_INV g_1600 (.D(w550), .C(w17), .nC(w248), .nQ(w2034) );
	ym3438_DLATCH_INV g_1601 (.D(w557), .C(w17), .nC(w248), .nQ(w2036) );
	ym3438_DLATCH_INVS g_1602 (.D(w552), .C(w18), .nC(w545), .nQ(w551) );
	ym3438_AND g_1603 (.Z(w552), .B(w2036), .A(w700) );
	ym3438_AON21SR g_1604 (.Q(w554), .nC2(w545), .C2(w18), .nC1(w248), .C1(w17), .B(1'b0), .A2(w551), .A1(w4464) );
	ym3438_AON21SR g_1605 (.Q(w587), .C2(w18), .nC2(w545), .C1(w17), .nC1(w248), .B(w554), .A2(w555), .A1(w4464) );
	ym3438_AON21SR g_1606 (.Q(w603), .nC2(w545), .C2(w18), .nC1(w248), .C1(w17), .B(w587), .A2(w535), .A1(w4464) );
	ym3438_AON21SR g_1607 (.Q(w619), .C2(w18), .nC2(w545), .C1(w17), .nC1(w248), .B(w603), .A2(w481), .A1(w4464) );
	ym3438_AON21SR g_1608 (.Q(w633), .nC2(w545), .C2(w18), .nC1(w248), .C1(w17), .B(w619), .A2(w533), .A1(w4464) );
	ym3438_AON21SR g_1609 (.Q(w655), .C2(w18), .nC2(w545), .C1(w17), .nC1(w248), .B(w633), .A2(w634), .A1(w4464) );
	ym3438_AON21SR g_1610 (.Q(w668), .nC2(w545), .C2(w18), .nC1(w248), .C1(w17), .B(w655), .A2(w669), .A1(w4464) );
	ym3438_AON21SR g_1611 (.Q(w699), .C2(w18), .nC2(w545), .C1(w17), .nC1(w248), .B(w668), .A2(w674), .A1(w4464) );
	ym3438_AON21SR g_1612 (.Q(w706), .nC2(w545), .C2(w18), .nC1(w248), .C1(w17), .B(w699), .A2(w698), .A1(w4464) );
	ym3438_AON21SR g_1613 (.Q(w963), .C2(w18), .nC2(w545), .C1(w17), .nC1(w248), .B(w706), .A2(w540), .A1(w4464) );
	ym3438_NOT g_1614 (.nZ(w2031), .A(w263) );
	ym3438_DLATCH_INV g_1615 (.D(w585), .C(w17), .nC(w248), .nQ(w2129) );
	ym3438_DLATCH_INV g_1616 (.D(w1197), .nC(w248), .C(w17), .nQ(w4034) );
	ym3438_NOT g_1617 (.nZ(w2055), .A(w2129) );
	ym3438_NOT g_1618 (.nZ(w4033), .A(w213) );
	ym3438_NOT g_1619 (.nZ(w614), .A(w4034) );
	ym3438_NOT g_1620 (.nZ(w17), .A(w4033) );
	ym3438_NOT g_1621 (.nZ(w4032), .A(w212) );
	ym3438_NOT g_1622 (.nZ(w248), .A(w4032) );
	ym3438_DLATCH_INVS g_1623 (.D(w2035), .nC(w545), .C(w18), .nQ(w555) );
	ym3438_DLATCH_INVS g_1624 (.D(w605), .C(w18), .nC(w545), .nQ(w535) );
	ym3438_DLATCH_INVS g_1625 (.D(w604), .nC(w545), .C(w18), .nQ(w481) );
	ym3438_DLATCH_INVS g_1626 (.D(w632), .C(w18), .nC(w545), .nQ(w533) );
	ym3438_DLATCH_INVS g_1627 (.D(w635), .nC(w545), .C(w18), .nQ(w634) );
	ym3438_DLATCH_INVS g_1628 (.D(w670), .C(w18), .nC(w545), .nQ(w669) );
	ym3438_DLATCH_INVS g_1629 (.D(w673), .nC(w545), .C(w18), .nQ(w674) );
	ym3438_DLATCH_INV g_1630 (.D(w558), .nC(w248), .C(w17), .nQ(w2037) );
	ym3438_DLATCH_INV g_1631 (.D(w607), .C(w17), .nC(w248), .nQ(w2060) );
	ym3438_DLATCH_INV g_1632 (.D(w553), .nC(w248), .C(w17), .nQ(w2059) );
	ym3438_DLATCH_INV g_1633 (.D(w584), .nC(w248), .C(w17), .nQ(w2058) );
	ym3438_SR_BIT g_1634 (.Q(w2061), .D(w601), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1635 (.Q(w2079), .D(w626), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SR_BIT g_1636 (.Q(w626), .D(w602), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_DLATCH_INV g_1637 (.D(w623), .nC(w248), .C(w17), .nQ(w622) );
	ym3438_DLATCH_INV g_1638 (.D(w609), .nC(w248), .C(w17), .nQ(w2064) );
	ym3438_DLATCH_INV g_1639 (.D(w638), .C(w17), .nC(w248), .nQ(w2132) );
	ym3438_DLATCH_INV g_1640 (.D(w624), .C(w17), .nC(w248), .nQ(w621) );
	ym3438_SR_BIT g_1641 (.Q(w2080), .D(w625), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1642 (.Q(w625), .D(w631), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1643 (.Q(w2107), .D(w660), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SR_BIT g_1644 (.Q(w660), .D(w349), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_DLATCH_INV g_1645 (.D(w659), .nC(w248), .C(w17), .nQ(w656) );
	ym3438_DLATCH_INV g_1646 (.D(w639), .nC(w248), .C(w17), .nQ(w2133) );
	ym3438_DLATCH_INVS g_1647 (.D(w707), .C(w18), .nC(w545), .nQ(w698) );
	ym3438_DLATCH_INVS g_1648 (.D(w709), .nC(w545), .C(w18), .nQ(w540) );
	ym3438_DLATCH_INV g_1649 (.D(w658), .C(w17), .nC(w248), .nQ(w657) );
	ym3438_DLATCH_INV g_1650 (.D(w675), .C(w17), .nC(w248), .nQ(w2141) );
	ym3438_DLATCH_INV g_1651 (.D(w676), .nC(w248), .C(w17), .nQ(w2142) );
	ym3438_DLATCH_INV g_1652 (.D(w694), .nC(w248), .C(w17), .nQ(w695) );
	ym3438_DLATCH_INV g_1653 (.D(w702), .C(w17), .nC(w248), .nQ(w701) );
	ym3438_DLATCH_INV g_1654 (.D(w712), .C(w17), .nC(w248), .nQ(w2152) );
	ym3438_DLATCH_INV g_1655 (.D(w728), .nC(w248), .C(w17), .nQ(w2153) );
	ym3438_DLATCH_INV g_1656 (.D(w2166), .nC(w248), .C(w17), .nQ(w724) );
	ym3438_FA g_1657 (.CO(w710), .S(w723), .CI(w2151), .A(w2153), .B(w724) );
	ym3438_AND g_1658 (.Z(w709), .B(w723), .A(w700) );
	ym3438_AND g_1659 (.Z(w707), .B(w708), .A(w700) );
	ym3438_AND g_1660 (.Z(w673), .B(w672), .A(w700) );
	ym3438_AND g_1661 (.Z(w670), .B(w671), .A(w700) );
	ym3438_AND g_1662 (.Z(w635), .B(w636), .A(w700) );
	ym3438_AND g_1663 (.Z(w632), .B(w637), .A(w700) );
	ym3438_AND g_1664 (.Z(w604), .B(w606), .A(w700) );
	ym3438_AND g_1665 (.Z(w605), .B(w2060), .A(w700) );
	ym3438_AND g_1666 (.Z(w2035), .B(w2037), .A(w700) );
	ym3438_NOT g_1667 (.nZ(w583), .A(w2058) );
	ym3438_NOT g_1668 (.nZ(w582), .A(w2059) );
	ym3438_NOT g_1669 (.nZ(w2063), .A(w2062) );
	ym3438_AND g_1670 (.Z(w2062), .B(w2061), .A(w586) );
	ym3438_AND g_1671 (.Z(w623), .B(w626), .A(w2063) );
	ym3438_AND g_1672 (.Z(w624), .B(w625), .A(w2063) );
	ym3438_AND g_1673 (.Z(w659), .B(w660), .A(w2063) );
	ym3438_AND g_1674 (.Z(w658), .B(w661), .A(w2063) );
	ym3438_AND g_1675 (.Z(w694), .B(w693), .A(w2063) );
	ym3438_AND g_1676 (.Z(w702), .B(w703), .A(w2063) );
	ym3438_AND g_1677 (.Z(w2166), .B(w725), .A(w2063) );
	ym3438_SR_BIT g_1678 (.Q(w661), .D(w348), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1679 (.Q(w2108), .D(w661), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1680 (.Q(w2109), .D(w693), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SR_BIT g_1681 (.Q(w693), .D(w347), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SR_BIT g_1682 (.Q(w2110), .D(w703), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1683 (.Q(w703), .D(w346), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1684 (.Q(w2159), .D(w725), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SR_BIT g_1685 (.Q(w725), .D(w345), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_EDGE_DET g_1686 (.D(w780), .nC1(w248), .C1(w17), .Q(w1334) );
	ym3438_CNT_BIT g_1687 (.CI(w4480), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545), .RES(w794), .Q(w781) );
	ym3438_CNT_BIT g_1688 (.CI(w261), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545), .RES(w794), .CO(w4480) );
	ym3438_AND g_1689 (.Z(w780), .B(w1982), .A(w252) );
	ym3438_AOI21 g_1690 (.A1(w261), .Z(w1983), .B(w262), .A2(w781) );
	ym3438_AND g_1691 (.Z(w782), .B(w127), .A(w1153) );
	ym3438_NOT g_1692 (.A(w1983), .nZ(w794) );
	ym3438_NOT g_1693 (.A(w1984), .nZ(w795) );
	ym3438_NOT g_1694 (.A(w1325), .nZ(w787) );
	ym3438_DLATCH_INV g_1695 (.D(w781), .nC(w248), .C(w17), .nQ(w1984) );
	ym3438_SR_BIT g_1696 (.Q(w1982), .D(w781), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SR_BIT g_1697 (.Q(w4479), .D(w1985), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_COMP_STR g_1698 (.Z(w962), .A(w4479) );
	ym3438_OR4 g_1699 (.Z(w1985), .B(w779), .A(w268), .C(w778), .D(w267) );
	ym3438_AND4 g_1700 (.Z(w796), .B(w793), .A(w1999), .C(w787), .D(w1998) );
	ym3438_DLATCH_INV g_1701 (.D(w1987), .C(w18), .nC(w545), .nQ(w1986) );
	ym3438_AND4 g_1702 (.Z(w788), .B(w798), .A(w1999), .C(w787), .D(w2010) );
	ym3438_AND g_1703 (.Z(w1987), .B(w1988), .A(w795) );
	ym3438_NOT g_1704 (.A(w1986), .nZ(w267) );
	ym3438_NOT g_1705 (.A(w1989), .nZ(w1988) );
	ym3438_AOI21 g_1706 (.A1(w1991), .Z(w1989), .B(w1990), .A2(w800) );
	ym3438_NOT g_1707 (.A(w1992), .nZ(w779) );
	ym3438_NOT g_1708 (.A(w793), .nZ(w798) );
	ym3438_AND g_1709 (.Z(w799), .B(w4028), .A(w795) );
	ym3438_AON22 g_1710 (.A1(w800), .Z(w4028), .B2(w1991), .A2(w776), .B1(w777) );
	ym3438_AND g_1711 (.Z(w1993), .B(w766), .A(w795) );
	ym3438_AON22 g_1712 (.A1(w800), .Z(w802), .B2(w776), .A2(w1994), .B1(w777) );
	ym3438_AND g_1713 (.Z(w4472), .B(w802), .A(w795) );
	ym3438_NOT g_1714 (.A(w4471), .nZ(w778) );
	ym3438_NOT g_1715 (.A(w4473), .nZ(w268) );
	ym3438_NOT g_1716 (.A(w1998), .nZ(w2010) );
	ym3438_DLATCH_INV g_1717 (.D(w799), .C(w18), .nC(w545), .nQ(w1992) );
	ym3438_DLATCH_INV g_1718 (.D(w4472), .C(w18), .nC(w545), .nQ(w4471) );
	ym3438_DLATCH_INV g_1719 (.D(w797), .C(w17), .nC(w248), .nQ(w800) );
	ym3438_DLATCH_INV g_1720 (.D(w1993), .C(w18), .nC(w545), .nQ(w4473) );
	ym3438_DLATCH_INV g_1721 (.D(w792), .C(w17), .nC(w248), .nQ(w801) );
	ym3438_AND g_1722 (.Z(w2011), .B(w1998), .A(w798) );
	ym3438_NOR3 g_1723 (.Z(w797), .B(w788), .A(w796), .C(w2011) );
	ym3438_NOR3 g_1724 (.Z(w792), .B(w817), .A(w789), .C(w2012) );
	ym3438_AND7 g_1725 (.Z(w2012), .B(w2014), .A(w2013), .C(w790), .D(w803), .E(w2015), .F(w804), .G(w1999) );
	ym3438_AND7 g_1726 (.Z(w789), .B(w2014), .A(w2013), .C(w790), .D(w803), .E(w791), .F(w804), .G(w4474) );
	ym3438_NOT g_1727 (.A(w1995), .nZ(w766) );
	ym3438_AOI21 g_1728 (.A1(w777), .Z(w1995), .B(w801), .A2(w1994) );
	ym3438_NOT g_1729 (.A(w800), .nZ(w777) );
	ym3438_DLATCH_INV g_1730 (.D(w765), .nC(w248), .C(w17), .nQ(w776) );
	ym3438_DLATCH_INV g_1731 (.D(w775), .nC(w248), .C(w17), .nQ(w1994) );
	ym3438_OR6 g_1732 (.Z(w4474), .B(w820), .A(w819), .C(w1996), .D(w1997), .E(w1998), .F(w1999) );
	ym3438_NAND4 g_1733 (.Z(w775), .B(w820), .A(w819), .C(w774), .D(w4029) );
	ym3438_NAND4 g_1734 (.Z(w765), .B(w1997), .A(w820), .C(w819), .D(w4029) );
	ym3438_DLATCH_INV g_1735 (.D(w818), .nC(w248), .C(w17), .nQ(w1991) );
	ym3438_NOT g_1736 (.A(w1996), .nZ(w4029) );
	ym3438_NAND4 g_1737 (.Z(w818), .B(w819), .A(w1996), .C(w820), .D(w774) );
	ym3438_NOT g_1738 (.A(w1997), .nZ(w774) );
	ym3438_DLATCH_INV g_1739 (.D(w773), .nC(w248), .C(w17), .nQ(w1990) );
	ym3438_NAND4 g_1740 (.Z(w773), .B(w819), .A(w1996), .C(w820), .D(w1997) );
	ym3438_NAND5 g_1741 (.Z(w2000), .B(w820), .A(w819), .C(w1997), .D(w1996), .E(w1998) );
	ym3438_NOT g_1742 (.A(w2016), .nZ(w804) );
	ym3438_AND7 g_1743 (.Z(w817), .B(w2014), .A(w2013), .C(w790), .D(w803), .E(w791), .F(w2016), .G(w1998) );
	ym3438_NOT g_1744 (.A(w2015), .nZ(w791) );
	ym3438_FA g_1745 (.S(w790), .CI(w4478), .A(w819), .B(w1326) );
	ym3438_FA g_1746 (.CO(w4478), .S(w803), .CI(w4477), .A(w820), .B(w1327) );
	ym3438_FA g_1747 (.CO(w4477), .S(w2015), .CI(w4476), .A(w1996), .B(w786) );
	ym3438_FA g_1748 (.CO(w4476), .S(w2016), .CI(1'b0), .A(w1997), .B(w1164) );
	ym3438_NAND g_1749 (.Z(w2014), .B(w820), .A(w819) );
	ym3438_AND3 g_1750 (.A(w2021), .B(w2020), .C(w1145), .Z(w2019) );
	ym3438_AON33 g_1751 (.A1(w2021), .Z(w816), .B2(w2022), .A2(w2020), .B1(w2021), .A3(w806), .B3(w1145) );
	ym3438_DLATCH_INV g_1752 (.D(w2019), .C(w17), .nC(w248), .nQ(w4082) );
	ym3438_DLATCH_INV g_1753 (.D(w210), .C(w17), .nC(w248), .nQ(w805) );
	ym3438_DLATCH_INV g_1754 (.D(w209), .C(w17), .nC(w248), .nQ(w4475) );
	ym3438_SR_BIT g_1755 (.Q(w2013), .D(w2018), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_DLATCH_INV g_1756 (.D(w816), .C(w17), .nC(w248), .nQ(w815) );
	ym3438_DLATCH_INV g_1757 (.D(w208), .C(w17), .nC(w248), .nQ(w814) );
	ym3438_AON333 g_1758 (.A1(w2021), .Z(w813), .B2(w2022), .A2(w2020), .B1(w2021), .A3(w808), .B3(w806), .C1(w785), .C2(w2020), .C3(w1145) );
	ym3438_DLATCH_INV g_1759 (.D(w813), .C(w17), .nC(w248), .nQ(w811) );
	ym3438_DLATCH_INV g_1760 (.D(w207), .C(w17), .nC(w248), .nQ(w812) );
	ym3438_AON3333 g_1761 (.A1(w2020), .Z(w2023), .B2(w2022), .A2(w2021), .B1(w2021), .A3(w783), .B3(w808), .C1(w785), .D2(w2022), .C2(w2020), .D1(w785), .C3(w806), .D3(w1145) );
	ym3438_DLATCH_INV g_1762 (.D(w2023), .C(w17), .nC(w248), .nQ(w810) );
	ym3438_DLATCH_INV g_1763 (.D(w206), .C(w17), .nC(w248), .nQ(w809) );
	ym3438_AON3333 g_1764 (.A1(w2020), .Z(w807), .B2(w2022), .A2(w2021), .B1(w2021), .A3(w1144), .B3(w783), .C1(w785), .D2(w2022), .C2(w2020), .D1(w785), .C3(w808), .D3(w806) );
	ym3438_OR5 g_1765 (.Z(w2018), .B(w207), .A(w206), .C(w208), .D(w210), .E(w209) );
	ym3438_DLATCH_INV g_1766 (.D(w807), .C(w17), .nC(w248), .nQ(w4083) );
	ym3438_COMP_WE g_1767 (.nZ(w785), .A(w784), .Z(w2021) );
	ym3438_COMP_WE g_1768 (.nZ(w2022), .A(w200), .Z(w2020) );
	ym3438_NOT g_1769 (.nZ(w545), .A(w4084) );
	ym3438_NOT g_1770 (.nZ(w4084), .A(w217) );
	ym3438_FA g_1771 (.CO(w761), .S(w760), .CI(1'b1), .A(1'b1), .B(w4083) );
	ym3438_DLATCH_INV g_1772 (.D(w760), .nC(w545), .C(w18), .nQ(w2009) );
	ym3438_OR g_1773 (.Z(w1999), .B(w2009), .A(w2001) );
	ym3438_FA g_1774 (.CO(w762), .S(w2008), .CI(w761), .A(w809), .B(w810) );
	ym3438_FA g_1775 (.CO(w764), .S(w763), .CI(w762), .A(w812), .B(w811) );
	ym3438_FA g_1776 (.CO(w768), .S(w767), .CI(w764), .A(w814), .B(w815) );
	ym3438_FA g_1777 (.CO(w770), .S(w769), .CI(w768), .A(w805), .B(w4082) );
	ym3438_FA g_1778 (.CO(w772), .S(w771), .CI(w770), .A(w4475), .B(1'b1) );
	ym3438_DLATCH_INV g_1779 (.D(w2008), .nC(w545), .C(w18), .nQ(w2007) );
	ym3438_OR g_1780 (.Z(w1998), .B(w2007), .A(w2001) );
	ym3438_DLATCH_INV g_1781 (.D(w763), .nC(w545), .C(w18), .nQ(w2006) );
	ym3438_OR g_1782 (.Z(w1997), .B(w2006), .A(w2001) );
	ym3438_OR g_1783 (.Z(w1996), .B(w2005), .A(w2001) );
	ym3438_OR g_1784 (.Z(w820), .B(w2004), .A(w2001) );
	ym3438_OR g_1785 (.Z(w819), .B(w2002), .A(w2001) );
	ym3438_DLATCH_INV g_1786 (.D(w772), .nC(w545), .C(w18), .nQ(w2001) );
	ym3438_DLATCH_INV g_1787 (.D(w771), .nC(w545), .C(w18), .nQ(w2002) );
	ym3438_DLATCH_INV g_1788 (.D(w769), .nC(w545), .C(w18), .nQ(w2004) );
	ym3438_DLATCH_INV g_1789 (.D(w767), .nC(w545), .C(w18), .nQ(w2005) );
	ym3438_SDELAY24 g_1790 (.A(w759), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545), .C3(w17), .C4(w18), .C5(w17), .C6(w18), .C7(w17), .C8(w18), .C9(w17), .C10(w18), .C11(w17), .C12(w18), .C13(w17), .C14(w18), .C15(w17), .C16(w18), .C17(w17), .C18(w18), .C19(w17), .C20(w18), .C21(w17), .C22(w18), .C23(w17), .C24(w18), .nC3(w248), .nC4(w545), .nC5(w248), .nC6(w545), .nC7(w248), .nC8(w545), .nC9(w248), .nC10(w545), .nC11(w248), .nC12(w545), .nC13(w248), .nC14(w545), .nC15(w248), .nC16(w545), .nC17(w248), .nC18(w545), .nC19(w248), .nC20(w545), .nC21(w248), .nC22(w545), .nC23(w248), .nC24(w545), .Q(w2191), .C25(w17), .C26(w18), .C27(w17), .C28(w18), .C29(w17), .C30(w18), .nC25(w248), .nC26(w545), .nC27(w248), .nC28(w545), .nC29(w248), .nC30(w545), .C36(w18), .nC36(w545), .C35(w17), .nC35(w248), .C34(w18), .nC34(w545), .C33(w17), .nC33(w248), .C32(w18), .nC32(w545), .C31(w17), .nC31(w248), .C42(w18), .nC42(w545), .C41(w17), .nC41(w248), .C40(w18), .nC40(w545), .C39(w17), .nC39(w248), .C38(w18), .nC38(w545), .C37(w17), .nC37(w248), .C44(w18), .nC44(w545), .C43(w17), .nC43(w248), .C46(w18), .nC46(w545), .C45(w17), .nC45(w248), .Q44(w758), .C48(w18), .nC48(w545), .C47(w17), .nC47(w248) );
	ym3438_SDELAY24 g_1791 (.A(w748), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545), .C3(w17), .C4(w18), .C5(w17), .C6(w18), .C7(w17), .C8(w18), .C9(w17), .C10(w18), .C11(w17), .C12(w18), .C13(w17), .C14(w18), .C15(w17), .C16(w18), .C17(w17), .C18(w18), .C19(w17), .C20(w18), .C21(w17), .C22(w18), .C23(w17), .C24(w18), .nC3(w248), .nC4(w545), .nC5(w248), .nC6(w545), .nC7(w248), .nC8(w545), .nC9(w248), .nC10(w545), .nC11(w248), .nC12(w545), .nC13(w248), .nC14(w545), .nC15(w248), .nC16(w545), .nC17(w248), .nC18(w545), .nC19(w248), .nC20(w545), .nC21(w248), .nC22(w545), .nC23(w248), .nC24(w545), .Q(w749), .C25(w17), .C26(w18), .C27(w17), .C28(w18), .C29(w17), .C30(w18), .nC25(w248), .nC26(w545), .nC27(w248), .nC28(w545), .nC29(w248), .nC30(w545), .C36(w18), .nC36(w545), .C35(w17), .nC35(w248), .C34(w18), .nC34(w545), .C33(w17), .nC33(w248), .C32(w18), .nC32(w545), .C31(w17), .nC31(w248), .C42(w18), .nC42(w545), .C41(w17), .nC41(w248), .C40(w18), .nC40(w545), .C39(w17), .nC39(w248), .C38(w18), .nC38(w545), .C37(w17), .nC37(w248), .C44(w18), .nC44(w545), .C43(w17), .nC43(w248), .C46(w18), .nC46(w545), .C45(w17), .nC45(w248), .C48(w18), .nC48(w545), .C47(w17), .nC47(w248), .Q44(w746) );
	ym3438_SDELAY24 g_1792 (.A(w2169), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545), .C3(w17), .C4(w18), .C5(w17), .C6(w18), .C7(w17), .C8(w18), .C9(w17), .C10(w18), .C11(w17), .C12(w18), .C13(w17), .C14(w18), .C15(w17), .C16(w18), .C17(w17), .C18(w18), .C19(w17), .C20(w18), .C21(w17), .C22(w18), .C23(w17), .C24(w18), .nC3(w248), .nC4(w545), .nC5(w248), .nC6(w545), .nC7(w248), .nC8(w545), .nC9(w248), .nC10(w545), .nC11(w248), .nC12(w545), .nC13(w248), .nC14(w545), .nC15(w248), .nC16(w545), .nC17(w248), .nC18(w545), .nC19(w248), .nC20(w545), .nC21(w248), .nC22(w545), .nC23(w248), .nC24(w545), .Q(w752), .C25(w17), .C26(w18), .C27(w17), .C28(w18), .C29(w17), .C30(w18), .nC25(w248), .nC26(w545), .nC27(w248), .nC28(w545), .nC29(w248), .nC30(w545), .C36(w18), .nC36(w545), .C35(w17), .nC35(w248), .C34(w18), .nC34(w545), .C33(w17), .nC33(w248), .C32(w18), .nC32(w545), .C31(w17), .nC31(w248), .C42(w18), .nC42(w545), .C41(w17), .nC41(w248), .C40(w18), .nC40(w545), .C39(w17), .nC39(w248), .C38(w18), .nC38(w545), .C37(w17), .nC37(w248), .C44(w18), .nC44(w545), .C43(w17), .nC43(w248), .C46(w18), .nC46(w545), .C45(w17), .nC45(w248), .C48(w18), .nC48(w545), .C47(w17), .nC47(w248), .Q44(w744) );
	ym3438_SDELAY24 g_1793 (.A(w743), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545), .C3(w17), .C4(w18), .C5(w17), .C6(w18), .C7(w17), .C8(w18), .C9(w17), .C10(w18), .C11(w17), .C12(w18), .C13(w17), .C14(w18), .C15(w17), .C16(w18), .C17(w17), .C18(w18), .C19(w17), .C20(w18), .C21(w17), .C22(w18), .C23(w17), .C24(w18), .nC3(w248), .nC4(w545), .nC5(w248), .nC6(w545), .nC7(w248), .nC8(w545), .nC9(w248), .nC10(w545), .nC11(w248), .nC12(w545), .nC13(w248), .nC14(w545), .nC15(w248), .nC16(w545), .nC17(w248), .nC18(w545), .nC19(w248), .nC20(w545), .nC21(w248), .nC22(w545), .nC23(w248), .nC24(w545), .C25(w17), .C26(w18), .C27(w17), .C28(w18), .C29(w17), .C30(w18), .nC25(w248), .nC26(w545), .nC27(w248), .nC28(w545), .nC29(w248), .nC30(w545), .C36(w18), .nC36(w545), .C35(w17), .nC35(w248), .C34(w18), .nC34(w545), .C33(w17), .nC33(w248), .C32(w18), .nC32(w545), .C31(w17), .nC31(w248), .C42(w18), .nC42(w545), .C41(w17), .nC41(w248), .C40(w18), .nC40(w545), .C39(w17), .nC39(w248), .C38(w18), .nC38(w545), .C37(w17), .nC37(w248), .C44(w18), .nC44(w545), .C43(w17), .nC43(w248), .C46(w18), .nC46(w545), .C45(w17), .nC45(w248), .C48(w18), .nC48(w545), .C47(w17), .nC47(w248), .Q(w2179) );
	ym3438_NOT g_1794 (.nZ(w18), .A(w4031) );
	ym3438_AND g_1795 (.Z(w328), .B(w2192), .A(w746) );
	ym3438_AND g_1796 (.Z(w192), .B(w758), .A(w2192) );
	ym3438_NOT g_1797 (.nZ(w4031), .A(w216) );
	ym3438_COMP_STR g_1798 (.Z(w4464), .A(w726) );
	ym3438_NAND3 g_1799 (.Z(w2154), .B(w27), .A(w1184), .C(w745) );
	ym3438_SR_BIT g_1800 (.Q(w2158), .D(w2157), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1801 (.Q(w2157), .D(w27), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1802 (.Q(w2169), .D(w2156), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1803 (.Q(w2156), .D(w745), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1804 (.Q(w2180), .D(w2155), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1805 (.Q(w2155), .D(w2154), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_AND g_1806 (.Z(w742), .B(w1185), .A(w2111) );
	ym3438_AND g_1807 (.Z(w2190), .B(w1179), .A(w2111) );
	ym3438_XOR g_1808 (.Z(w2165), .B(w2179), .A(w2190) );
	ym3438_OR g_1809 (.Z(w2189), .B(w742), .A(w2165) );
	ym3438_AND3 g_1810 (.Z(w743), .B(w27), .A(w2189), .C(w744) );
	ym3438_XOR g_1811 (.Z(w2188), .B(w1173), .A(w2179) );
	ym3438_AND g_1812 (.Z(w2187), .B(w744), .A(w2188) );
	ym3438_SR_BIT g_1813 (.Q(w2164), .D(w2187), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_NOT g_1814 (.nZ(w741), .A(w2169) );
	ym3438_NOT g_1815 (.nZ(w4087), .A(w4086) );
	ym3438_COMP_STR g_1816 (.nZ(w2042), .A(w2164), .Z(w2043) );
	ym3438_AON22 g_1817 (.A1(w266), .Z(w736), .B2(w270), .A2(w299), .B1(w317) );
	ym3438_COMP_WE g_1818 (.A(w2158), .nZ(w266), .Z(w270) );
	ym3438_NOT g_1819 (.A(w2160), .nZ(w2072) );
	ym3438_AOI21 g_1820 (.A1(w2174), .Z(w2160), .B(w737), .A2(w2161) );
	ym3438_NOT g_1821 (.A(w737), .nZ(w2161) );
	ym3438_NOT g_1822 (.A(w736), .nZ(w2170) );
	ym3438_NOT g_1823 (.A(w314), .nZ(w2171) );
	ym3438_SR_BIT g_1824 (.Q(w738), .D(w2172), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1825 (.Q(w2172), .D(w2175), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_AND3 g_1826 (.Z(w2175), .B(w2111), .A(w27), .C(w727) );
	ym3438_AND3 g_1827 (.Z(w2177), .B(w2111), .A(w1178), .C(w27) );
	ym3438_NOT g_1828 (.A(w4085), .nZ(w733) );
	ym3438_NOT g_1829 (.A(w2169), .nZ(w4448) );
	ym3438_COMP_STR g_1830 (.Z(w731), .A(w2178), .nZ(w732) );
	ym3438_AOI22 g_1831 (.A1(w2186), .Z(w2192), .B2(w2177), .A2(w745), .B1(w744) );
	ym3438_AND4 g_1832 (.Z(w4030), .B(w2191), .A(w2171), .C(w2200), .D(w2174) );
	ym3438_OR6 g_1833 (.Z(w748), .B(w750), .A(w754), .C(w733), .D(w747), .F(w2196), .E(w2185) );
	ym3438_NOR g_1834 (.Z(w4085), .B(w2196), .A(w740) );
	ym3438_AND g_1835 (.Z(w2178), .B(w752), .A(w4448) );
	ym3438_AND4 g_1836 (.Z(w740), .B(w2174), .A(w736), .C(w2180), .D(w2198) );
	ym3438_AND g_1837 (.Z(w2181), .B(w2200), .A(w2199) );
	ym3438_NOT g_1838 (.A(w2181), .nZ(w2198) );
	ym3438_NOT g_1839 (.A(w2182), .nZ(w264) );
	ym3438_NAND5 g_1840 (.Z(w2182), .B(w737), .A(w755), .C(w2199), .D(w2169), .E(w2200) );
	ym3438_NOT g_1841 (.A(w2183), .nZ(w265) );
	ym3438_NOR g_1842 (.Z(w2183), .B(w2184), .A(w751) );
	ym3438_AND3 g_1843 (.Z(w2184), .B(w2170), .A(w749), .C(w2174) );
	ym3438_AND5 g_1844 (.Z(w751), .B(w2171), .A(w2170), .C(w2191), .D(w2200), .E(w2174) );
	ym3438_AND g_1845 (.Z(w750), .B(w741), .A(w2174) );
	ym3438_AND3 g_1846 (.Z(w754), .B(w749), .A(w2191), .C(w2174) );
	ym3438_AND3 g_1847 (.Z(w747), .B(w749), .A(w2199), .C(w2174) );
	ym3438_AND4 g_1848 (.Z(w2185), .B(w2174), .A(w2200), .C(w314), .D(w2191) );
	ym3438_NOT g_1849 (.nZ(w2186), .A(w744) );
	ym3438_NOT g_1850 (.nZ(w2199), .A(w2191) );
	ym3438_NOT g_1851 (.nZ(w2200), .A(w749) );
	ym3438_AND4 g_1852 (.Z(w2201), .B(w2199), .A(w2174), .C(w271), .D(w2200) );
	ym3438_OR6 g_1853 (.Z(w759), .B(w733), .A(w750), .C(w754), .D(w4030), .E(w2196), .F(w2201) );
	ym3438_SR_BIT g_1854 (.Q(w312), .D(w4447), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1855 (.Q(w296), .D(w2193), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1856 (.Q(w2193), .D(w1165), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1857 (.Q(w316), .D(w2194), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1858 (.Q(w2194), .D(w1104), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1859 (.Q(w295), .D(w2195), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1860 (.Q(w2195), .D(w1106), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_NOT g_1861 (.A(w271), .nZ(w755) );
	ym3438_NOT g_1862 (.A(w214), .nZ(w2196) );
	ym3438_SR_BIT g_1863 (.Q(w737), .D(w2000), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SR_BIT g_1864 (.Q(w4447), .D(w1105), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SR_BIT g_1865 (.Q(w311), .D(w2167), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SR_BIT g_1866 (.Q(w2167), .D(w1107), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SR_BIT g_1867 (.Q(w739), .D(w2176), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_SR_BIT g_1868 (.Q(w2176), .D(w2177), .C1(w17), .C2(w18), .nC1(w248), .nC2(w545) );
	ym3438_NOT g_1869 (.A(w752), .nZ(w2168) );
	ym3438_NOR g_1870 (.Z(w756), .B(w753), .A(w738) );
	ym3438_AND g_1871 (.Z(w753), .B(w2168), .A(w2169) );
	ym3438_AOI21 g_1872 (.A1(w752), .Z(w2173), .B(w753), .A2(w739) );
	ym3438_COMP_STR g_1873 (.Z(w2174), .A(w2173) );
	ym3438_SR_BIT g_1874 (.Q(w2197), .D(w756), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_SR_BIT g_1875 (.Q(w757), .D(w2197), .nC1(w248), .nC2(w545), .C1(w17), .C2(w18) );
	ym3438_NOT g_1876 (.A(w214), .nZ(w262) );
	ym3438_AND g_1877 (.A(w27), .Z(w1173), .B(w26) );
	ym3438_AON22 g_1878 (.A1(w31), .Z(w27), .B2(w30), .A2(w28), .B1(w29) );
	ym3438_NOR g_1879 (.A(w2205), .Z(w2202), .B(w156) );
	ym3438_NOR g_1880 (.A(w4316), .Z(w4315), .B(w156) );
	ym3438_AOI22 g_1881 (.A1(w31), .Z(w2205), .B2(w338), .A2(w2203), .B1(w2204) );
	ym3438_AOI22 g_1882 (.A1(w30), .Z(w4316), .B2(w338), .A2(w327), .B1(w326) );
	ym3438_AND4 g_1883 (.A(w1104), .B(w1106), .Z(w1165), .C(w1105), .D(w1107) );
	ym3438_AON22 g_1884 (.A1(w2206), .Z(w26), .B2(w321), .A2(w28), .B1(w29) );
	ym3438_SDELAY12 g_1885 (.A(w2202), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w31) );
	ym3438_SDELAY12 g_1886 (.A(w4315), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w30) );
	ym3438_SDELAY12 g_1887 (.A(w2212), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w322) );
	ym3438_SDELAY12 g_1888 (.A(w4313), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w323) );
	ym3438_SDELAY12 g_1889 (.A(w4319), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w324) );
	ym3438_SDELAY12 g_1890 (.A(w2214), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w325) );
	ym3438_AON22 g_1891 (.A1(w322), .Z(w195), .B2(w323), .A2(w28), .B1(w29) );
	ym3438_NOR g_1892 (.A(w4314), .Z(w4313), .B(w156) );
	ym3438_NOR g_1893 (.A(w2213), .Z(w2212), .B(w156) );
	ym3438_AOI22 g_1894 (.A1(w322), .Z(w2213), .B2(w336), .A2(w2203), .B1(w2204) );
	ym3438_AOI22 g_1895 (.A1(w323), .Z(w4314), .B2(w336), .A2(w327), .B1(w326) );
	ym3438_AON22 g_1896 (.A1(w324), .Z(w334), .B2(w325), .A2(w28), .B1(w29) );
	ym3438_AND g_1897 (.A(w215), .Z(w2204), .B(w2215) );
	ym3438_AND g_1898 (.A(w2216), .Z(w326), .B(w2215) );
	ym3438_AOI22 g_1899 (.A1(w324), .Z(w4320), .B2(w332), .A2(w2203), .B1(w2204) );
	ym3438_NOR g_1900 (.A(w4320), .Z(w4319), .B(w156) );
	ym3438_NOR g_1901 (.A(w4321), .Z(w2214), .B(w156) );
	ym3438_AOI22 g_1902 (.A1(w325), .Z(w4321), .B2(w332), .A2(w327), .B1(w326) );
	ym3438_NOT g_1903 (.A(w2204), .nZ(w2203) );
	ym3438_NOT g_1904 (.A(w326), .nZ(w327) );
	ym3438_NOT g_1913 (.nZ(w121), .A(w2246) );
	ym3438_SR_BIT g_1914 (.D(w1081), .C1(w213), .C2(w216), .nC1(w212), .nC2(w217), .Q(w1087) );
	ym3438_SLATCH g_1915 (.nQ(w1108), .C(w1085), .nC(w1088), .D(w1067) );
	ym3438_SR_BIT g_1916 (.D(w1084), .C1(w213), .C2(w216), .nC1(w212), .nC2(w217), .Q(w2252) );
	ym3438_NOT g_1917 (.nZ(w1103), .A(w4080) );
	ym3438_TRI g_1918 (.Z(w1156), .A(w1108), .E(w1089) );
	ym3438_TRI g_1919 (.Z(w1155), .A(w1109), .E(w1089) );
	ym3438_NOR g_1920 (.Z(w1079), .A(w1108), .B(w1109) );
	ym3438_SLATCH g_1921 (.nQ(w1109), .C(w1085), .nC(w1088), .D(w1161) );
	ym3438_NOT g_1922 (.nZ(w1085), .A(w1088) );
	ym3438_NOT g_1923 (.nZ(w2261), .A(w1172) );
	ym3438_NOT g_1924 (.nZ(w2263), .A(w2262) );
	ym3438_AND g_1925 (.Z(w1089), .B(w2261), .A(w1088) );
	ym3438_AOI21 g_1926 (.Z(w2264), .B(w121), .A1(w2263), .A2(w1110) );
	ym3438_SR_BIT g_1927 (.D(w2264), .C1(w213), .C2(w216), .nC1(w212), .nC2(w217), .Q(w2265) );
	ym3438_NOT g_1928 (.nZ(w1110), .A(w2265) );
	ym3438_TRI g_1929 (.Z(w1078), .A(w1110), .E(w1089) );
	ym3438_NOT g_1930 (.nZ(w1088), .A(w4081) );
	ym3438_NOT g_1931 (.nZ(w1101), .A(w214) );
	ym3438_NOT g_1932 (.nZ(w214), .A(w1095) );
	ym3438_CNT_BIT g_1933 (.CI(w1110), .C1(w213), .C2(w216), .nC1(w212), .nC2(w217), .RES(w1101), .CO(w2266) );
	ym3438_CNT_BIT g_1934 (.CI(w2266), .C1(w213), .C2(w216), .nC1(w212), .nC2(w217), .RES(w1101), .CO(w2267) );
	ym3438_CNT_BIT g_1935 (.CI(w2267), .C1(w213), .C2(w216), .nC1(w212), .nC2(w217), .RES(w1101), .CO(w2284) );
	ym3438_CNT_BIT g_1936 (.CI(w2284), .C1(w213), .C2(w216), .nC1(w212), .nC2(w217), .RES(w1101), .CO(w2285) );
	ym3438_CNT_BIT g_1937 (.CI(w2285), .C1(w213), .C2(w216), .nC1(w212), .nC2(w217), .RES(w1101), .CO(w2286) );
	ym3438_OR g_1938 (.Z(w2262), .B(w2286), .A(w1101) );
	ym3438_TRI g_1939 (.Z(w112), .A(w1100), .E(w1096) );
	ym3438_TRI g_1940 (.Z(w108), .A(w2271), .E(w1096) );
	ym3438_TRI g_1941 (.Z(w958), .A(w2272), .E(w1096) );
	ym3438_TRI g_1942 (.Z(w959), .A(w2273), .E(w1096) );
	ym3438_TRI g_1943 (.Z(w960), .A(w2287), .E(w1096) );
	ym3438_TRI g_1944 (.Z(w132), .A(w1099), .E(w1096) );
	ym3438_TRI g_1945 (.Z(w961), .A(w1098), .E(w1096) );
	ym3438_TRI g_1946 (.Z(w123), .A(w2270), .E(w1096) );
	ym3438_NOT g_1947 (.nZ(w120), .A(w2268) );
	ym3438_NOT g_1948 (.nZ(w2268), .A(w2269) );
	ym3438_SLATCH g_1949 (.Q(w2270), .C(w1093), .nC(w1097), .D(w1314) );
	ym3438_SLATCH g_1950 (.Q(w2269), .C(w1093), .nC(w1097), .D(w2260) );
	ym3438_SLATCH g_1951 (.Q(w1098), .C(w1093), .nC(w1097), .D(w1313) );
	ym3438_SLATCH g_1952 (.Q(w1099), .C(w1093), .nC(w1097), .D(w1077) );
	ym3438_SLATCH g_1953 (.Q(w2287), .C(w1093), .nC(w1097), .D(w1075) );
	ym3438_SLATCH g_1954 (.Q(w2273), .C(w1093), .nC(w1097), .D(w1317) );
	ym3438_SLATCH g_1955 (.Q(w2272), .C(w1093), .nC(w1097), .D(w1312) );
	ym3438_SLATCH g_1956 (.Q(w2271), .C(w1093), .nC(w1097), .D(w1311) );
	ym3438_SLATCH g_1957 (.Q(w1100), .C(w1093), .nC(w1097), .D(w1074) );
	ym3438_NAND3 g_1958 (.Z(w2276), .B(w1091), .A(w1092), .C(w2258) );
	ym3438_NOT g_1959 (.nZ(w1093), .A(w2274) );
	ym3438_NOT g_1960 (.nZ(w1097), .A(w1093) );
	ym3438_NAND g_1961 (.Z(w2275), .B(w2276), .A(w1091) );
	ym3438_NAND g_1962 (.Z(w2274), .B(w2259), .A(w2258) );
	ym3438_NOT g_1963 (.nZ(w1096), .A(w2275) );
	ym3438_NOT g_1964 (.nZ(w1076), .A(w2277) );
	ym3438_NOT g_1965 (.nZ(w2277), .A(w2276) );
	ym3438_NOT g_1966 (.nZ(w2246), .A(w2247) );
	ym3438_NOT g_1967 (.nZ(w2248), .A(w1087) );
	ym3438_NOT g_1968 (.nZ(w1086), .A(w216) );
	ym3438_AND g_1969 (.Z(w2247), .A(w2248), .B(w1081) );
	ym3438_SLATCH g_1970 (.Q(w1081), .C(w216), .nC(w1086), .D(w2249) );
	ym3438_SRFF g_1971 (.Q(w1080), .nQ(w2250), .S(w1083), .R(w1081) );
	ym3438_SYNC_SRFF g_1972 (.Q(w2249), .C(w213), .S(w1080), .R(w2250) );
	ym3438_SYNC_SRFF g_1973 (.Q(w2254), .C(w213), .S(w2255), .R(w2256) );
	ym3438_SRFF g_1974 (.Q(w2255), .nQ(w2256), .S(w2257), .R(w1084) );
	ym3438_SLATCH g_1975 (.Q(w1084), .C(w216), .nC(w2253), .D(w2254) );
	ym3438_NOT g_1976 (.nZ(w2253), .A(w216) );
	ym3438_NOT g_1977 (.nZ(w1082), .A(w2252) );
	ym3438_NOT g_1978 (.nZ(w4080), .A(w2251) );
	ym3438_AND g_1979 (.Z(w2251), .A(w1082), .B(w1084) );
	ym3438_AND4 g_1980 (.D(w1090), .Z(w1083), .B(w2259), .A(w2258), .C(w1091) );
	ym3438_AND3 g_1981 (.Z(w1094), .B(w2259), .A(w2258), .C(w1304) );
	ym3438_NAND5 g_1982 (.D(w1304), .Z(w4081), .B(w2258), .A(w1091), .C(w1092), .E(w2260) );
	ym3438_NOT g_1983 (.nZ(w2260), .A(w1318) );
	ym3438_NOT g_1984 (.nZ(w1095), .A(w1315) );
	ym3438_NOT g_1985 (.A(w1095), .nZ(w1091) );
	ym3438_NOT g_1986 (.nZ(w1092), .A(w1154) );
	ym3438_NOT g_1987 (.nZ(w1304), .A(w1090) );
	ym3438_NOT g_1988 (.nZ(w2259), .A(w1316) );
	ym3438_NOT g_1989 (.nZ(w2258), .A(w1152) );
	ym3438_OR g_1990 (.Z(w2257), .B(w1095), .A(w1094) );
	ym3438_AOI22 g_1991 (.A1(w2378), .Z(w2375), .B2(w332), .A2(w2379), .B1(w2369) );
	ym3438_NOR g_1992 (.A(w2375), .Z(w2376), .B(w156) );
	ym3438_SDELAY12 g_1993 (.A(w2376), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2378) );
	ym3438_AOI22 g_1994 (.A1(w2377), .Z(w4213), .B2(w336), .A2(w2379), .B1(w2369) );
	ym3438_NOR g_1995 (.A(w4213), .Z(w4214), .B(w156) );
	ym3438_SDELAY12 g_1996 (.A(w4214), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2377) );
	ym3438_AOI22 g_1997 (.A1(w2374), .Z(w2371), .B2(w337), .A2(w2379), .B1(w2369) );
	ym3438_NOR g_1998 (.A(w2371), .Z(w2372), .B(w156) );
	ym3438_SDELAY12 g_1999 (.A(w2372), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2374) );
	ym3438_AOI22 g_2000 (.A1(w2373), .Z(w2370), .B2(w338), .A2(w2379), .B1(w2369) );
	ym3438_NOR g_2001 (.A(w2370), .Z(w4212), .B(w156) );
	ym3438_SDELAY12 g_2002 (.A(w4212), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2373) );
	ym3438_AOI22 g_2003 (.A1(w2368), .Z(w2365), .B2(w331), .A2(w2379), .B1(w2369) );
	ym3438_NOR g_2004 (.A(w2365), .Z(w2366), .B(w156) );
	ym3438_SDELAY12 g_2005 (.A(w2366), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2368) );
	ym3438_AOI22 g_2006 (.A1(w2367), .Z(w2364), .B2(w330), .A2(w2379), .B1(w2369) );
	ym3438_NOR g_2007 (.A(w2364), .Z(w4215), .B(w156) );
	ym3438_SDELAY12 g_2008 (.A(w4215), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2367) );
	ym3438_AOI22 g_2009 (.A1(w2382), .Z(w4216), .B2(w329), .A2(w2379), .B1(w2369) );
	ym3438_NOR g_2010 (.A(w4216), .Z(w4217), .B(w156) );
	ym3438_SDELAY12 g_2011 (.A(w4217), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2382) );
	ym3438_AOI22 g_2012 (.A1(w2381), .Z(w2380), .B2(w331), .A2(w2210), .B1(w2211) );
	ym3438_NOR g_2013 (.A(w2380), .Z(w4211), .B(w156) );
	ym3438_SDELAY12 g_2014 (.A(w4211), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2381) );
	ym3438_AOI22 g_2015 (.A1(w2363), .Z(w2360), .B2(w338), .A2(w2210), .B1(w2211) );
	ym3438_NOR g_2016 (.A(w2360), .Z(w2361), .B(w156) );
	ym3438_SDELAY12 g_2017 (.A(w2361), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2363) );
	ym3438_AOI22 g_2018 (.A1(w2362), .Z(w2359), .B2(w337), .A2(w2210), .B1(w2211) );
	ym3438_NOR g_2019 (.A(w2359), .Z(w4210), .B(w156) );
	ym3438_SDELAY12 g_2020 (.A(w4210), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2362) );
	ym3438_AOI22 g_2021 (.A1(w2358), .Z(w2355), .B2(w336), .A2(w2210), .B1(w2211) );
	ym3438_NOR g_2022 (.A(w2355), .Z(w2356), .B(w156) );
	ym3438_SDELAY12 g_2023 (.A(w2356), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2358) );
	ym3438_AOI22 g_2024 (.A1(w2357), .Z(w2354), .B2(w332), .A2(w2210), .B1(w2211) );
	ym3438_NOR g_2025 (.A(w2354), .Z(w4209), .B(w156) );
	ym3438_SDELAY12 g_2026 (.A(w4209), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2357) );
	ym3438_AOI22 g_2027 (.A1(w226), .Z(w2221), .B2(w340), .A2(w2218), .B1(w2217) );
	ym3438_NOR g_2028 (.A(w2221), .Z(w2222), .B(w156) );
	ym3438_SDELAY12 g_2029 (.A(w2222), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w226) );
	ym3438_AOI22 g_2030 (.A1(w2220), .Z(w2223), .B2(w329), .A2(w2218), .B1(w2217) );
	ym3438_NOR g_2031 (.A(w2223), .Z(w4139), .B(w156) );
	ym3438_SDELAY12 g_2032 (.A(w4139), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2220) );
	ym3438_AOI22 g_2033 (.A1(w2219), .Z(w2224), .B2(w331), .A2(w2218), .B1(w2217) );
	ym3438_NOR g_2034 (.A(w2224), .Z(w2225), .B(w156) );
	ym3438_SDELAY12 g_2035 (.A(w2225), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2219) );
	ym3438_AOI22 g_2036 (.A1(w225), .Z(w2226), .B2(w338), .A2(w2218), .B1(w2217) );
	ym3438_NOR g_2037 (.A(w2226), .Z(w4140), .B(w156) );
	ym3438_SDELAY12 g_2038 (.A(w4140), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w225) );
	ym3438_AOI22 g_2039 (.A1(w224), .Z(w2227), .B2(w337), .A2(w2218), .B1(w2217) );
	ym3438_NOR g_2040 (.A(w2227), .Z(w2228), .B(w156) );
	ym3438_SDELAY12 g_2041 (.A(w2228), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w224) );
	ym3438_AOI22 g_2042 (.A1(w2232), .Z(w2229), .B2(w336), .A2(w2218), .B1(w2217) );
	ym3438_NOR g_2043 (.A(w2229), .Z(w4141), .B(w156) );
	ym3438_SDELAY12 g_2044 (.A(w4141), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2232) );
	ym3438_AOI22 g_2045 (.A1(w2233), .Z(w2230), .B2(w332), .A2(w2218), .B1(w2217) );
	ym3438_NOR g_2046 (.A(w2230), .Z(w2231), .B(w156) );
	ym3438_SDELAY12 g_2047 (.A(w2231), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2233) );
	ym3438_AOI22 g_2048 (.A1(w133), .Z(w2386), .B2(w340), .A2(w144), .B1(w2389) );
	ym3438_NOR g_2049 (.A(w2386), .Z(w4170), .B(w156) );
	ym3438_SDELAY12 g_2050 (.A(w4170), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w133) );
	ym3438_AOI22 g_2051 (.A1(w134), .Z(w2387), .B2(w329), .A2(w144), .B1(w2389) );
	ym3438_NOR g_2052 (.A(w2387), .Z(w2388), .B(w156) );
	ym3438_SDELAY12 g_2053 (.A(w2388), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w134) );
	ym3438_AOI22 g_2054 (.A1(w137), .Z(w2390), .B2(w330), .A2(w144), .B1(w2389) );
	ym3438_NOR g_2055 (.A(w2390), .Z(w4171), .B(w156) );
	ym3438_SDELAY12 g_2056 (.A(w4171), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w137) );
	ym3438_AOI22 g_2057 (.A1(w136), .Z(w2391), .B2(w331), .A2(w144), .B1(w2389) );
	ym3438_NOR g_2058 (.A(w2391), .Z(w2392), .B(w156) );
	ym3438_SDELAY12 g_2059 (.A(w2392), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w136) );
	ym3438_AOI22 g_2060 (.A1(w138), .Z(w2393), .B2(w338), .A2(w144), .B1(w2389) );
	ym3438_NOR g_2061 (.A(w2393), .Z(w4172), .B(w156) );
	ym3438_SDELAY12 g_2062 (.A(w4172), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w138) );
	ym3438_AOI22 g_2063 (.A1(w139), .Z(w2394), .B2(w337), .A2(w144), .B1(w2389) );
	ym3438_NOR g_2064 (.A(w2394), .Z(w2395), .B(w156) );
	ym3438_SDELAY12 g_2065 (.A(w2395), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w139) );
	ym3438_AOI22 g_2066 (.A1(w142), .Z(w2396), .B2(w336), .A2(w144), .B1(w2389) );
	ym3438_NOR g_2067 (.A(w2396), .Z(w4173), .B(w156) );
	ym3438_SDELAY12 g_2068 (.A(w4173), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w142) );
	ym3438_AOI22 g_2069 (.A1(w141), .Z(w2397), .B2(w332), .A2(w144), .B1(w2389) );
	ym3438_NOR g_2070 (.A(w2397), .Z(w2398), .B(w156) );
	ym3438_SDELAY12 g_2071 (.A(w2398), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w141) );
	ym3438_AOI22 g_2072 (.A1(w179), .B2(w332), .A2(w2401), .B1(w2400), .Z(w4242) );
	ym3438_NOR g_2073 (.A(w4242), .Z(w4244), .B(w156) );
	ym3438_SDELAY12 g_2074 (.A(w4244), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w179) );
	ym3438_AOI22 g_2075 (.A1(w178), .B2(w336), .A2(w2401), .B1(w2400), .Z(w4243) );
	ym3438_NOR g_2076 (.A(w4243), .Z(w2399), .B(w156) );
	ym3438_SDELAY12 g_2077 (.A(w2399), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w178) );
	ym3438_AOI22 g_2078 (.A1(w177), .B2(w337), .A2(w2401), .B1(w2400), .Z(w4246) );
	ym3438_NOR g_2079 (.A(w4246), .Z(w4245), .B(w156) );
	ym3438_SDELAY12 g_2080 (.A(w4245), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w177) );
	ym3438_AOI22 g_2081 (.A1(w176), .B2(w338), .A2(w2401), .B1(w2400), .Z(w4247) );
	ym3438_NOR g_2082 (.A(w4247), .Z(w2402), .B(w156) );
	ym3438_SDELAY12 g_2083 (.A(w2402), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w176) );
	ym3438_AOI22 g_2084 (.A1(w175), .B2(w331), .A2(w2401), .B1(w2400), .Z(w4250) );
	ym3438_NOR g_2085 (.A(w4250), .Z(w4249), .B(w156) );
	ym3438_SDELAY12 g_2086 (.A(w4249), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w175) );
	ym3438_AOI22 g_2087 (.A1(w174), .B2(w340), .A2(w2401), .B1(w2400), .Z(w4251) );
	ym3438_NOR g_2088 (.A(w4251), .Z(w4248), .B(w156) );
	ym3438_SDELAY12 g_2089 (.A(w4248), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w174) );
	ym3438_AOI22 g_2090 (.A1(w173), .B2(w329), .A2(w2404), .B1(w2403), .Z(w4256) );
	ym3438_NOR g_2091 (.A(w4256), .Z(w4257), .B(w156) );
	ym3438_SDELAY12 g_2092 (.A(w4257), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w173) );
	ym3438_AOI22 g_2093 (.A1(w172), .B2(w330), .A2(w2404), .B1(w2403), .Z(w4254) );
	ym3438_NOR g_2094 (.A(w4254), .Z(w4253), .B(w156) );
	ym3438_SDELAY12 g_2095 (.A(w4253), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w172) );
	ym3438_AOI22 g_2096 (.A1(w171), .B2(w331), .A2(w2404), .B1(w2403), .Z(w4255) );
	ym3438_NOR g_2097 (.A(w4255), .Z(w4252), .B(w156) );
	ym3438_SDELAY12 g_2098 (.A(w4252), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w171) );
	ym3438_AOI22 g_2099 (.A1(w170), .B2(w338), .A2(w2404), .B1(w2403), .Z(w4260) );
	ym3438_NOR g_2100 (.A(w4260), .Z(w4259), .B(w156) );
	ym3438_SDELAY12 g_2101 (.A(w4259), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w170) );
	ym3438_AOI22 g_2102 (.A1(w169), .B2(w337), .A2(w2404), .B1(w2403), .Z(w4261) );
	ym3438_NOR g_2103 (.A(w4261), .Z(w4258), .B(w156) );
	ym3438_SDELAY12 g_2104 (.A(w4258), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w169) );
	ym3438_AOI22 g_2105 (.A1(w168), .B2(w336), .A2(w2404), .B1(w2403), .Z(w4264) );
	ym3438_NOR g_2106 (.A(w4264), .Z(w4263), .B(w156) );
	ym3438_SDELAY12 g_2107 (.A(w4263), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w168) );
	ym3438_AOI22 g_2108 (.A1(w2405), .B2(w332), .A2(w2404), .B1(w2403), .Z(w4265) );
	ym3438_NOR g_2109 (.A(w4265), .Z(w4262), .B(w156) );
	ym3438_SDELAY12 g_2110 (.A(w4262), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2405) );
	ym3438_SDELAY12 g_2111 (.A(w2322), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2324) );
	ym3438_NOR g_2112 (.A(w2323), .Z(w2322), .B(w156) );
	ym3438_AOI22 g_2113 (.A1(w2324), .Z(w2323), .B2(w340), .A2(w149), .B1(w148) );
	ym3438_SDELAY12 g_2114 (.A(w4182), .Q(w2325), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .nC9(w25), .nC10(w24), .C3(w23), .C4(w22) );
	ym3438_NOR g_2115 (.A(w4188), .Z(w4182), .B(w156) );
	ym3438_AOI22 g_2116 (.A1(w2325), .Z(w4188), .B2(w329), .A2(w149), .B1(w148) );
	ym3438_SDELAY12 g_2117 (.A(w2326), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w135) );
	ym3438_NOR g_2118 (.A(w2327), .Z(w2326), .B(w156) );
	ym3438_AOI22 g_2119 (.A1(w135), .Z(w2327), .B2(w330), .A2(w149), .B1(w148) );
	ym3438_SDELAY12 g_2120 (.A(w4183), .Q(w2328), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .nC9(w25), .nC10(w24), .C3(w23), .C4(w22) );
	ym3438_NOR g_2121 (.A(w4187), .Z(w4183), .B(w156) );
	ym3438_AOI22 g_2122 (.A1(w2328), .Z(w4187), .B2(w331), .A2(w149), .B1(w148) );
	ym3438_SDELAY12 g_2123 (.A(w2329), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w151) );
	ym3438_NOR g_2124 (.A(w2331), .Z(w2329), .B(w156) );
	ym3438_AOI22 g_2125 (.A1(w151), .Z(w2331), .B2(w338), .A2(w149), .B1(w148) );
	ym3438_SDELAY12 g_2126 (.A(w4184), .Q(w150), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .nC9(w25), .nC10(w24), .C3(w23), .C4(w22) );
	ym3438_NOR g_2127 (.A(w2330), .Z(w4184), .B(w156) );
	ym3438_AOI22 g_2128 (.A1(w150), .Z(w2330), .B2(w337), .A2(w149), .B1(w148) );
	ym3438_SDELAY12 g_2129 (.A(w2332), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2334) );
	ym3438_NOR g_2130 (.A(w2333), .Z(w2332), .B(w156) );
	ym3438_AOI22 g_2131 (.A1(w2334), .Z(w2333), .B2(w336), .A2(w149), .B1(w148) );
	ym3438_SDELAY12 g_2132 (.A(w4185), .Q(w140), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .nC9(w25), .nC10(w24), .C3(w23), .C4(w22) );
	ym3438_NOR g_2133 (.A(w4186), .Z(w4185), .B(w156) );
	ym3438_AOI22 g_2134 (.A1(w140), .Z(w4186), .B2(w332), .A2(w149), .B1(w148) );
	ym3438_SDELAY12 g_2135 (.A(w2335), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2337) );
	ym3438_NOR g_2136 (.A(w2336), .Z(w2335), .B(w156) );
	ym3438_AOI22 g_2137 (.A1(w2337), .Z(w2336), .B2(w332), .A2(w2339), .B1(w2340) );
	ym3438_SDELAY12 g_2138 (.A(w4292), .Q(w2338), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .nC9(w25), .nC10(w24), .C3(w23), .C4(w22) );
	ym3438_NOR g_2139 (.A(w4293), .Z(w4292), .B(w156) );
	ym3438_AOI22 g_2140 (.A1(w2338), .Z(w4293), .B2(w336), .A2(w2339), .B1(w2340) );
	ym3438_SDELAY12 g_2141 (.A(w2341), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w157) );
	ym3438_NOR g_2142 (.A(w2342), .Z(w2341), .B(w156) );
	ym3438_AOI22 g_2143 (.A1(w157), .Z(w2342), .B2(w337), .A2(w2339), .B1(w2340) );
	ym3438_SDELAY12 g_2144 (.A(w4294), .Q(w158), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .nC9(w25), .nC10(w24), .C3(w23), .C4(w22) );
	ym3438_NOR g_2145 (.A(w4295), .Z(w4294), .B(w156) );
	ym3438_AOI22 g_2146 (.A1(w158), .Z(w4295), .B2(w338), .A2(w2339), .B1(w2340) );
	ym3438_SDELAY12 g_2147 (.A(w2343), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w159) );
	ym3438_NOR g_2148 (.A(w2344), .Z(w2343), .B(w156) );
	ym3438_AOI22 g_2149 (.A1(w159), .Z(w2344), .B2(w331), .A2(w2339), .B1(w2340) );
	ym3438_SDELAY12 g_2150 (.A(w4296), .Q(w160), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .nC9(w25), .nC10(w24), .C3(w23), .C4(w22) );
	ym3438_NOR g_2151 (.A(w4297), .Z(w4296), .B(w156) );
	ym3438_AOI22 g_2152 (.A1(w160), .Z(w4297), .B2(w340), .A2(w2339), .B1(w2340) );
	ym3438_SDELAY12 g_2153 (.A(w4298), .Q(w161), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .nC9(w25), .nC10(w24), .C3(w23), .C4(w22) );
	ym3438_NOR g_2154 (.A(w4299), .Z(w4298), .B(w156) );
	ym3438_AOI22 g_2155 (.A1(w161), .Z(w4299), .B2(w329), .A2(w2347), .B1(w2348) );
	ym3438_SDELAY12 g_2156 (.A(w2345), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w162) );
	ym3438_NOR g_2157 (.A(w2346), .Z(w2345), .B(w156) );
	ym3438_AOI22 g_2158 (.A1(w162), .Z(w2346), .B2(w330), .A2(w2347), .B1(w2348) );
	ym3438_SDELAY12 g_2159 (.A(w4304), .Q(w166), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .nC9(w25), .nC10(w24), .C3(w23), .C4(w22) );
	ym3438_NOR g_2160 (.A(w4305), .Z(w4304), .B(w156) );
	ym3438_AOI22 g_2161 (.A1(w166), .Z(w4305), .B2(w332), .A2(w2347), .B1(w2348) );
	ym3438_SDELAY12 g_2162 (.A(w2351), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2353) );
	ym3438_NOR g_2163 (.A(w2352), .Z(w2351), .B(w156) );
	ym3438_AOI22 g_2164 (.A1(w2353), .Z(w2352), .B2(w336), .A2(w2347), .B1(w2348) );
	ym3438_SDELAY12 g_2165 (.A(w4302), .Q(w165), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .nC9(w25), .nC10(w24), .C3(w23), .C4(w22) );
	ym3438_NOR g_2166 (.A(w4303), .Z(w4302), .B(w156) );
	ym3438_AOI22 g_2167 (.A1(w165), .Z(w4303), .B2(w337), .A2(w2347), .B1(w2348) );
	ym3438_SDELAY12 g_2168 (.A(w2349), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w164) );
	ym3438_NOR g_2169 (.A(w2350), .Z(w2349), .B(w156) );
	ym3438_AOI22 g_2170 (.A1(w164), .Z(w2350), .B2(w338), .A2(w2347), .B1(w2348) );
	ym3438_SDELAY12 g_2171 (.A(w4300), .Q(w163), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .nC9(w25), .nC10(w24), .C3(w23), .C4(w22) );
	ym3438_NOR g_2172 (.A(w4301), .Z(w4300), .B(w156) );
	ym3438_AOI22 g_2173 (.A1(w163), .Z(w4301), .B2(w331), .A2(w2347), .B1(w2348) );
	ym3438_SDELAY12 g_2174 (.A(w2283), .Q(w227), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .nC9(w25), .nC10(w24) );
	ym3438_NOR g_2175 (.A(w2288), .Z(w2283), .B(w156) );
	ym3438_AOI22 g_2176 (.A1(w227), .Z(w2288), .B2(w340), .A2(w2289), .B1(w218) );
	ym3438_SDELAY12 g_2177 (.A(w2290), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w230) );
	ym3438_NOR g_2178 (.A(w2292), .Z(w2290), .B(w156) );
	ym3438_AOI22 g_2179 (.A1(w230), .Z(w2292), .B2(w329), .A2(w2289), .B1(w218) );
	ym3438_SDELAY12 g_2180 (.A(w4158), .Q(w229), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .nC9(w25), .nC10(w24) );
	ym3438_NOR g_2181 (.A(w2291), .Z(w4158), .B(w156) );
	ym3438_AOI22 g_2182 (.A1(w229), .Z(w2291), .B2(w331), .A2(w2289), .B1(w218) );
	ym3438_AON22 g_2183 (.A1(w2219), .Z(w201), .B2(w229), .A2(w28), .B1(w29) );
	ym3438_SDELAY12 g_2184 (.A(w2293), .Q(w2296), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24) );
	ym3438_NOR g_2185 (.A(w2295), .Z(w2293), .B(w156) );
	ym3438_AOI22 g_2186 (.A1(w2296), .Z(w2295), .B2(w338), .A2(w2289), .B1(w218) );
	ym3438_AON22 g_2187 (.A1(w225), .Z(w221), .B2(w2296), .A2(w28), .B1(w29) );
	ym3438_SDELAY12 g_2188 (.A(w4159), .Q(w228), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .nC9(w25), .nC10(w24) );
	ym3438_NOR g_2189 (.A(w2294), .Z(w4159), .B(w156) );
	ym3438_AOI22 g_2190 (.A1(w228), .Z(w2294), .B2(w337), .A2(w2289), .B1(w218) );
	ym3438_AON22 g_2191 (.A1(w224), .Z(w220), .B2(w228), .A2(w28), .B1(w29) );
	ym3438_SDELAY12 g_2192 (.A(w2297), .Q(w223), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24) );
	ym3438_NOR g_2193 (.A(w2299), .Z(w2297), .B(w156) );
	ym3438_AOI22 g_2194 (.A1(w223), .Z(w2299), .B2(w336), .A2(w2289), .B1(w218) );
	ym3438_AON22 g_2195 (.A1(w2232), .Z(w202), .B2(w223), .A2(w28), .B1(w29) );
	ym3438_SDELAY12 g_2196 (.A(w4160), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w222) );
	ym3438_NOR g_2197 (.A(w2298), .Z(w4160), .B(w156) );
	ym3438_AOI22 g_2198 (.A1(w222), .Z(w2298), .B2(w332), .A2(w2289), .B1(w218) );
	ym3438_AON22 g_2199 (.A1(w2233), .Z(w219), .B2(w222), .A2(w28), .B1(w29) );
	ym3438_SDELAY12 g_2200 (.A(w2300), .Q(w2303), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24) );
	ym3438_NOR g_2201 (.A(w2302), .Z(w2300), .B(w156) );
	ym3438_AOI22 g_2202 (.A1(w2303), .Z(w2302), .B2(w332), .A2(w2281), .B1(w2282) );
	ym3438_AON22 g_2203 (.A1(w2357), .Z(w4196), .B2(w2303), .A2(w28), .B1(w29) );
	ym3438_SDELAY12 g_2204 (.A(w4220), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2304) );
	ym3438_NOR g_2205 (.A(w2301), .Z(w4220), .B(w156) );
	ym3438_AOI22 g_2206 (.A1(w2304), .B2(w336), .A2(w2281), .B1(w2282), .Z(w2301) );
	ym3438_AON22 g_2207 (.A1(w2358), .Z(w2383), .B2(w2304), .A2(w28), .B1(w29) );
	ym3438_SDELAY12 g_2208 (.A(w2305), .Q(w189), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24) );
	ym3438_NOR g_2209 (.A(w2306), .Z(w2305), .B(w156) );
	ym3438_AOI22 g_2210 (.A1(w189), .B2(w337), .A2(w2281), .B1(w2282), .Z(w2306) );
	ym3438_AON22 g_2211 (.A1(w2362), .Z(w2241), .B2(w189), .A2(w28), .B1(w29) );
	ym3438_SDELAY12 g_2212 (.A(w4218), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2307) );
	ym3438_NOR g_2213 (.A(w4219), .Z(w4218), .B(w156) );
	ym3438_AOI22 g_2214 (.A1(w2307), .B2(w338), .A2(w2281), .B1(w2282), .Z(w4219) );
	ym3438_AON22 g_2215 (.A1(w2363), .Z(w2240), .B2(w2307), .A2(w28), .B1(w29) );
	ym3438_SDELAY12 g_2216 (.A(w2308), .Q(w2311), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24) );
	ym3438_NOR g_2217 (.A(w2310), .Z(w2308), .B(w156) );
	ym3438_AOI22 g_2218 (.A1(w2311), .B2(w331), .A2(w2281), .B1(w2282), .Z(w2310) );
	ym3438_AON22 g_2219 (.A1(w2381), .Z(w193), .B2(w2311), .A2(w28), .B1(w29) );
	ym3438_SDELAY12 g_2220 (.A(w4221), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2312) );
	ym3438_NOR g_2221 (.A(w2309), .Z(w4221), .B(w156) );
	ym3438_AOI22 g_2222 (.A1(w2312), .B2(w329), .A2(w2316), .B1(w2317), .Z(w2309) );
	ym3438_AON22 g_2223 (.A1(w2382), .Z(w333), .B2(w2312), .A2(w28), .B1(w29) );
	ym3438_SDELAY12 g_2224 (.A(w2313), .Q(w188), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24) );
	ym3438_NOR g_2225 (.A(w2314), .Z(w2313), .B(w156) );
	ym3438_AOI22 g_2226 (.A1(w188), .B2(w330), .A2(w2316), .B1(w2317), .Z(w2314) );
	ym3438_AON22 g_2227 (.A1(w2367), .Z(w335), .B2(w188), .A2(w28), .B1(w29) );
	ym3438_SDELAY12 g_2228 (.A(w4222), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2315) );
	ym3438_NOR g_2229 (.A(w4223), .Z(w4222), .B(w156) );
	ym3438_AOI22 g_2230 (.A1(w2315), .B2(w331), .A2(w2316), .B1(w2317), .Z(w4223) );
	ym3438_AON22 g_2231 (.A1(w2368), .Z(w232), .B2(w2315), .A2(w28), .B1(w29) );
	ym3438_SDELAY12 g_2232 (.A(w4226), .Q(w2319), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24) );
	ym3438_NOR g_2233 (.A(w2318), .Z(w4226), .B(w156) );
	ym3438_AOI22 g_2234 (.A1(w2319), .B2(w338), .A2(w2316), .B1(w2317), .Z(w2318) );
	ym3438_AON22 g_2235 (.A1(w2373), .Z(w4013), .B2(w2319), .A2(w28), .B1(w29) );
	ym3438_SDELAY12 g_2236 (.A(w4224), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2320) );
	ym3438_NOR g_2237 (.A(w4225), .Z(w4224), .B(w156) );
	ym3438_AOI22 g_2238 (.A1(w2320), .B2(w337), .A2(w2316), .B1(w2317), .Z(w4225) );
	ym3438_AON22 g_2239 (.A1(w2374), .Z(w2384), .B2(w2320), .A2(w28), .B1(w29) );
	ym3438_SDELAY12 g_2240 (.A(w4227), .Q(w186), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24) );
	ym3438_NOR g_2241 (.A(w2321), .Z(w4227), .B(w156) );
	ym3438_AOI22 g_2242 (.A1(w186), .B2(w336), .A2(w2316), .B1(w2317), .Z(w2321) );
	ym3438_AON22 g_2243 (.A1(w2377), .Z(w185), .B2(w186), .A2(w28), .B1(w29) );
	ym3438_SDELAY12 g_2244 (.A(w4228), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w187) );
	ym3438_NOR g_2245 (.A(w4229), .Z(w4228), .B(w156) );
	ym3438_AOI22 g_2246 (.A1(w187), .B2(w332), .A2(w2316), .B1(w2317), .Z(w4229) );
	ym3438_AON22 g_2247 (.A1(w2378), .Z(w2385), .B2(w187), .A2(w28), .B1(w29) );
	ym3438_AON22 g_2248 (.A1(w2220), .Z(w200), .B2(w230), .A2(w28), .B1(w29) );
	ym3438_AON22 g_2249 (.A1(w226), .Z(w784), .B2(w227), .A2(w28), .B1(w29) );
	ym3438_AON22 g_2250 (.A1(w2324), .Z(w1104), .B2(w133), .A2(w28), .B1(w29) );
	ym3438_AON22 g_2251 (.A1(w2325), .Z(w1106), .B2(w134), .A2(w28), .B1(w29) );
	ym3438_AON22 g_2252 (.A1(w135), .Z(w1105), .B2(w137), .A2(w28), .B1(w29) );
	ym3438_AON22 g_2253 (.A1(w2328), .Z(w1107), .B2(w136), .A2(w28), .B1(w29) );
	ym3438_AON22 g_2254 (.A1(w151), .Z(w2406), .B2(w138), .A2(w28), .B1(w29) );
	ym3438_AON22 g_2255 (.A1(w150), .Z(w339), .B2(w139), .A2(w28), .B1(w29) );
	ym3438_AON22 g_2256 (.A1(w2334), .Z(w154), .B2(w142), .A2(w28), .B1(w29) );
	ym3438_AON22 g_2257 (.A1(w140), .Z(w2407), .B2(w141), .A2(w28), .B1(w29) );
	ym3438_AON22 g_2258 (.A1(w2337), .B2(w179), .A2(w28), .B1(w29), .Z(w2408) );
	ym3438_AON22 g_2259 (.A1(w2338), .B2(w178), .A2(w28), .B1(w29), .Z(w344) );
	ym3438_AON22 g_2260 (.A1(w157), .B2(w177), .A2(w28), .B1(w29), .Z(w343) );
	ym3438_AON22 g_2261 (.A1(w158), .B2(w176), .A2(w28), .B1(w29), .Z(w2409) );
	ym3438_AON22 g_2262 (.A1(w159), .B2(w175), .A2(w28), .B1(w29), .Z(w342) );
	ym3438_AON22 g_2263 (.A1(w160), .B2(w174), .A2(w28), .B1(w29), .Z(w180) );
	ym3438_AON22 g_2264 (.A1(w161), .B2(w173), .A2(w28), .B1(w29), .Z(w345) );
	ym3438_AON22 g_2265 (.A1(w162), .B2(w172), .A2(w28), .B1(w29), .Z(w346) );
	ym3438_AON22 g_2266 (.A1(w163), .B2(w171), .A2(w28), .B1(w29), .Z(w347) );
	ym3438_AON22 g_2267 (.A1(w164), .B2(w170), .A2(w28), .B1(w29), .Z(w348) );
	ym3438_AON22 g_2268 (.A1(w165), .B2(w169), .A2(w28), .B1(w29), .Z(w349) );
	ym3438_AON22 g_2269 (.A1(w2353), .B2(w168), .A2(w28), .B1(w29), .Z(w631) );
	ym3438_AON22 g_2270 (.A1(w166), .B2(w2405), .A2(w28), .B1(w29), .Z(w602) );
	ym3438_NOT g_2271 (.A(w214), .nZ(w156) );
	ym3438_NOT g_2272 (.A(w2234), .nZ(w24) );
	ym3438_NOT g_2273 (.A(w2235), .nZ(w22) );
	ym3438_NOT g_2274 (.A(w2236), .nZ(w23) );
	ym3438_NOT g_2275 (.A(w2237), .nZ(w25) );
	ym3438_NOT g_2276 (.A(w341), .nZ(w28) );
	ym3438_NOT g_2277 (.A(w2280), .nZ(w29) );
	ym3438_NOT g_2278 (.A(w2340), .nZ(w2339) );
	ym3438_NOT g_2279 (.A(w148), .nZ(w149) );
	ym3438_NOT g_2280 (.A(w2389), .nZ(w144) );
	ym3438_NOT g_2281 (.A(w2400), .nZ(w2401) );
	ym3438_NOT g_2282 (.A(w218), .nZ(w2289) );
	ym3438_NOT g_2283 (.A(w341), .nZ(w2280) );
	ym3438_NOT g_2284 (.A(w2282), .nZ(w2281) );
	ym3438_NOT g_2285 (.A(w328), .nZ(w191) );
	ym3438_NOT g_2286 (.A(w192), .nZ(w190) );
	ym3438_NOT g_2287 (.A(w212), .nZ(w2237) );
	ym3438_NOT g_2288 (.A(w2217), .nZ(w2218) );
	ym3438_NOT g_2289 (.A(w217), .nZ(w2234) );
	ym3438_NOT g_2290 (.A(w213), .nZ(w2236) );
	ym3438_NOT g_2291 (.A(w2211), .nZ(w2210) );
	ym3438_AND g_2292 (.A(w215), .Z(w2217), .B(w203) );
	ym3438_AND g_2293 (.A(w215), .Z(w2211), .B(w211) );
	ym3438_NOT g_2294 (.A(w216), .nZ(w2235) );
	ym3438_OR4 g_2295 (.A(w2242), .Z(w209), .B(w146), .C(w181), .D(w2238) );
	ym3438_AND g_2296 (.A(w199), .Z(w2242), .B(w201) );
	ym3438_OR4 g_2297 (.A(w2243), .Z(w210), .B(w147), .C(w184), .D(w2239) );
	ym3438_AND g_2298 (.A(w199), .Z(w2243), .B(w221) );
	ym3438_OR4 g_2299 (.A(w2245), .Z(w208), .B(w197), .C(w183), .D(w2244) );
	ym3438_AND g_2300 (.A(w199), .Z(w2245), .B(w220) );
	ym3438_OR4 g_2301 (.A(w2278), .Z(w207), .B(w198), .C(w182), .D(w205) );
	ym3438_AND g_2302 (.A(w199), .Z(w2278), .B(w202) );
	ym3438_OR4 g_2303 (.A(w2279), .Z(w206), .B(w155), .C(w153), .D(w204) );
	ym3438_AND g_2304 (.A(w199), .Z(w2279), .B(w219) );
	ym3438_AND g_2305 (.A(w2216), .Z(w218), .B(w203) );
	ym3438_AND g_2306 (.A(w211), .Z(w2282), .B(w2216) );
	ym3438_AND g_2307 (.A(w191), .Z(w199), .B(w190) );
	ym3438_AND g_2308 (.A(w193), .Z(w2238), .B(w196) );
	ym3438_AND g_2309 (.A(w2240), .Z(w2239), .B(w196) );
	ym3438_AND g_2310 (.A(w2241), .Z(w2244), .B(w196) );
	ym3438_AND g_2311 (.A(w2383), .Z(w205), .B(w196) );
	ym3438_AND g_2312 (.A(w4196), .Z(w204), .B(w196) );
	ym3438_AND g_2313 (.A(w192), .Z(w153), .B(w328) );
	ym3438_AND g_2314 (.A(w190), .Z(w196), .B(w328) );
	ym3438_AND g_2315 (.A(w192), .Z(w152), .B(w191) );
	ym3438_FA g_2316 (.S(w730), .A(w1305), .B(1'b1), .CI(w2070) );
	ym3438_SDELAY12 g_2317 (.A(w4312), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w2206) );
	ym3438_SDELAY12 g_2318 (.A(w2207), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24), .C3(w23), .C4(w22), .C5(w23), .C6(w22), .C7(w23), .C8(w22), .C9(w23), .C10(w22), .C11(w23), .C12(w22), .C13(w23), .C14(w22), .C15(w23), .C16(w22), .C17(w23), .C18(w22), .C19(w23), .C20(w22), .C21(w23), .C22(w22), .C23(w23), .C24(w22), .nC3(w25), .nC4(w24), .nC5(w25), .nC6(w24), .nC7(w25), .nC8(w24), .nC9(w25), .nC10(w24), .nC11(w25), .nC12(w24), .nC13(w25), .nC14(w24), .nC15(w25), .nC16(w24), .nC17(w25), .nC18(w24), .nC19(w25), .nC20(w24), .nC21(w25), .nC22(w24), .nC23(w25), .nC24(w24), .Q(w321) );
	ym3438_NOR g_2319 (.A(w2208), .Z(w4312), .B(w156) );
	ym3438_AOI22 g_2320 (.A1(w2206), .Z(w2208), .B2(w337), .A2(w2203), .B1(w2204) );
	ym3438_NOR g_2321 (.A(w2209), .Z(w2207), .B(w156) );
	ym3438_AOI22 g_2322 (.A1(w321), .Z(w2209), .B2(w337), .A2(w327), .B1(w326) );
	ym3438_AND g_2323 (.A(w215), .Z(w2340), .B(w145) );
	ym3438_AND g_2324 (.A(w215), .Z(w148), .B(w143) );
	ym3438_AND g_2325 (.A(w153), .Z(w181), .B(w2406) );
	ym3438_AND g_2326 (.A(w153), .Z(w184), .B(w339) );
	ym3438_AND g_2327 (.A(w153), .Z(w182), .B(w2407) );
	ym3438_AND g_2328 (.A(w153), .Z(w183), .B(w154) );
	ym3438_AND g_2329 (.A(w152), .Z(w155), .B(w2408) );
	ym3438_AND g_2330 (.A(w152), .Z(w198), .B(w344) );
	ym3438_AND g_2331 (.A(w152), .Z(w197), .B(w343) );
	ym3438_AND g_2332 (.A(w152), .Z(w147), .B(w2409) );
	ym3438_AND g_2333 (.A(w152), .Z(w146), .B(w342) );
	ym3438_AND g_2334 (.A(w2216), .Z(w2389), .B(w143) );
	ym3438_AND g_2335 (.A(w2216), .Z(w2400), .B(w145) );
	ym3438_CNT_BIT g_40 (.CI(w831), .Q(w1349), .C1(w57), .C2(w56), .nC1(w834), .nC2(w833), .RES(w827), .CO(w845) );
	ym3438_NOT g_2336 (.A(w1485), .nZ(w924) );
	ym3438_DLATCH_INV g_2337 (.nQ(w3883), .D(w3191), .C(w2545), .nC(w1150) );
	ym3438_SR_BIT g_2338 (.Q(w3191), .D(w1145), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_COMP_STR g_2339 (.A(w3884), .Z(w2552) );
	ym3438_AND g_2340 (.Z(w3884), .B(w2540), .A(w2542) );
	ym3438_AND g_2341 (.Z(w4150), .B(w2540), .A(w2543) );
	ym3438_AND g_2342 (.Z(w3885), .B(w2542), .A(w2541) );
	ym3438_COMP_STR g_2343 (.A(w4150), .Z(w2553) );
	ym3438_COMP_STR g_2344 (.A(w3885), .Z(w2741) );
	ym3438_COMP_STR g_2345 (.A(w3886), .Z(w2572) );
	ym3438_AND g_2346 (.Z(w3886), .B(w2543), .A(w2541) );
	ym3438_COMP_WE g_2347 (.A(w4366), .nZ(w2541), .Z(w2540) );
	ym3438_COMP_WE g_2348 (.A(w3887), .nZ(w2543), .Z(w2542) );
	ym3438_NOT g_2349 (.A(w3888), .nZ(w3887) );
	ym3438_DLATCH_INV g_2350 (.nQ(w3888), .D(w2544), .C(w2545), .nC(w1150) );
	ym3438_SR_BIT g_2351 (.Q(w2544), .D(w808), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_COMP_WE g_2352 (.A(w2571), .nZ(w2558), .Z(w2557) );
	ym3438_COMP_WE g_2353 (.A(w2570), .nZ(w2563), .Z(w2555) );
	ym3438_COMP_WE g_2354 (.A(w2569), .nZ(w2562), .Z(w2556) );
	ym3438_COMP_WE g_2355 (.A(w2568), .nZ(w2565), .Z(w2554) );
	ym3438_NOT g_2356 (.A(w3890), .nZ(w3889) );
	ym3438_NAND5 g_2357 (.Z(w3890), .B(w2565), .A(w2561), .C(w2556), .D(w2563), .E(w2557) );
	ym3438_NAND5 g_2358 (.Z(w3896), .B(w2565), .A(w2561), .C(w2555), .D(w2558), .E(w2556) );
	ym3438_NOT g_2359 (.A(w3896), .nZ(w2567) );
	ym3438_NOT g_2360 (.A(w3895), .nZ(w2566) );
	ym3438_NOT g_2361 (.A(w3894), .nZ(w3893) );
	ym3438_NOT g_2362 (.A(w3892), .nZ(w3891) );
	ym3438_NAND5 g_2363 (.Z(w3892), .B(w2563), .A(w2557), .C(w2562), .D(w2561), .E(w2554) );
	ym3438_NAND5 g_2364 (.Z(w3894), .B(w2563), .A(w2558), .C(w2562), .D(w2561), .E(w2554) );
	ym3438_NAND5 g_2365 (.Z(w3895), .B(w2565), .A(w2561), .C(w2556), .D(w2555), .E(w2557) );
	ym3438_NOT g_2366 (.A(w3897), .nZ(w2581) );
	ym3438_DLATCH_INV g_2367 (.nQ(w3897), .D(w2576), .C(w2545), .nC(w1150) );
	ym3438_FA g_2368 (.S(w2576), .CI(w2601), .A(w2602), .B(w2575) );
	ym3438_DLATCH_INV g_2369 (.nQ(w2575), .D(w2577), .C(w2546), .nC(w1149) );
	ym3438_AOI22 g_2370 (.A2(w2548), .A1(w2574), .Z(w2577), .B2(w2547), .B1(1'b0) );
	ym3438_NOT g_2371 (.A(w3913), .nZ(w2643) );
	ym3438_DLATCH_INV g_2372 (.nQ(w3913), .D(w2641), .C(w2545), .nC(w1150) );
	ym3438_FA g_2373 (.CO(w2601), .S(w2641), .CI(w2642), .A(w2602), .B(w2638) );
	ym3438_DLATCH_INV g_2374 (.nQ(w2638), .D(w2637), .C(w2546), .nC(w1149) );
	ym3438_AOI22 g_2375 (.A2(w2548), .A1(w2636), .Z(w2637), .B2(w2547), .B1(1'b0) );
	ym3438_NOT g_2376 (.A(w3898), .nZ(w2662) );
	ym3438_DLATCH_INV g_2377 (.nQ(w3898), .D(w2640), .C(w2545), .nC(w1150) );
	ym3438_FA g_2378 (.CO(w2642), .S(w2640), .CI(w2661), .A(w2602), .B(w2639) );
	ym3438_DLATCH_INV g_2379 (.nQ(w2639), .D(w3914), .C(w2546), .nC(w1149) );
	ym3438_AOI22 g_2380 (.A2(w2548), .A1(w2634), .Z(w3914), .B2(w2547), .B1(1'b0) );
	ym3438_AON2222 g_2381 (.A2(1'b0), .Z(w2634), .B2(w2812), .C2(w2553), .B1(w2741), .D1(w1142), .D2(w2552), .A1(w2572), .C1(w1143) );
	ym3438_NOT g_2382 (.A(w3912), .nZ(w2694) );
	ym3438_DLATCH_INV g_2383 (.nQ(w3912), .D(w2693), .C(w2545), .nC(w1150) );
	ym3438_FA g_2384 (.CO(w2661), .S(w2693), .CI(w2692), .A(w2602), .B(w2691) );
	ym3438_DLATCH_INV g_2385 (.nQ(w2691), .D(w2688), .C(w2546), .nC(w1149) );
	ym3438_AOI22 g_2386 (.A2(w2548), .A1(w2686), .Z(w2688), .B2(w2547), .B1(1'b0) );
	ym3438_AON2222 g_2387 (.A2(w2812), .Z(w2686), .B2(w1143), .C2(w2553), .B1(w2741), .D1(w3970), .D2(w2552), .A1(w2572), .C1(w1142) );
	ym3438_NOT g_2388 (.A(w3899), .nZ(w2725) );
	ym3438_DLATCH_INV g_2389 (.nQ(w3899), .D(w2690), .C(w2545), .nC(w1150) );
	ym3438_FA g_2390 (.CO(w2692), .S(w2690), .CI(w2724), .A(w2602), .B(w2689) );
	ym3438_DLATCH_INV g_2391 (.nQ(w2689), .D(w2687), .C(w2546), .nC(w1149) );
	ym3438_AOI22 g_2392 (.A2(w2548), .A1(w2685), .Z(w2687), .B2(w2547), .B1(w2574) );
	ym3438_AON2222 g_2393 (.A2(w1143), .Z(w2685), .B2(w1142), .C2(w2553), .B1(w2741), .D1(w2684), .D2(w2552), .A1(w2572), .C1(w3970) );
	ym3438_NOT g_2394 (.A(w3911), .nZ(w2764) );
	ym3438_DLATCH_INV g_2395 (.nQ(w3911), .D(w2762), .C(w2545), .nC(w1150) );
	ym3438_FA g_2396 (.CO(w2724), .S(w2762), .CI(w2761), .A(w2602), .B(w2760) );
	ym3438_DLATCH_INV g_2397 (.nQ(w2760), .D(w2758), .C(w2546), .nC(w1149) );
	ym3438_AOI22 g_2398 (.A2(w2548), .A1(w2750), .Z(w2758), .B2(w2547), .B1(w2636) );
	ym3438_AON2222 g_2399 (.A2(w1142), .Z(w2750), .B2(w3970), .C2(w2553), .B1(w2741), .D1(w2749), .D2(w2552), .A1(w2572), .C1(w2684) );
	ym3438_NOT g_2400 (.A(w3905), .nZ(w2840) );
	ym3438_DLATCH_INV g_2401 (.nQ(w3905), .D(w2763), .C(w2545), .nC(w1150) );
	ym3438_FA g_2402 (.CO(w2761), .S(w2763), .CI(w2796), .A(w2602), .B(w2759) );
	ym3438_DLATCH_INV g_2403 (.nQ(w2759), .D(w2757), .C(w2546), .nC(w1149) );
	ym3438_AOI22 g_2404 (.A2(w2548), .A1(w2751), .Z(w2757), .B2(w2547), .B1(w2634) );
	ym3438_AON2222 g_2405 (.A2(w3970), .Z(w2751), .B2(w2684), .C2(w2553), .B1(w2741), .D1(w2756), .D2(w2552), .A1(w2572), .C1(w2749) );
	ym3438_NOT g_2406 (.A(w3910), .nZ(w2834) );
	ym3438_DLATCH_INV g_2407 (.nQ(w3910), .D(w2833), .C(w2545), .nC(w1150) );
	ym3438_FA g_2408 (.CO(w2796), .S(w2833), .CI(w2832), .A(w2602), .B(w2831) );
	ym3438_DLATCH_INV g_2409 (.nQ(w2831), .D(w2828), .C(w2546), .nC(w1149) );
	ym3438_AOI22 g_2410 (.A2(w2548), .A1(w2826), .Z(w2828), .B2(w2547), .B1(w2686) );
	ym3438_AON2222 g_2411 (.A2(w2684), .Z(w2826), .B2(w2749), .C2(w2553), .B1(w2741), .D1(w2823), .D2(w2552), .A1(w2572), .C1(w2756) );
	ym3438_NOT g_2412 (.A(w3904), .nZ(w2905) );
	ym3438_DLATCH_INV g_2413 (.nQ(w3904), .D(w2830), .C(w2545), .nC(w1150) );
	ym3438_FA g_2414 (.CO(w2832), .S(w2830), .CI(w2863), .A(w2602), .B(w2829) );
	ym3438_DLATCH_INV g_2415 (.nQ(w2829), .D(w2827), .C(w2546), .nC(w1149) );
	ym3438_AOI22 g_2416 (.A2(w2548), .A1(w2825), .Z(w2827), .B2(w2547), .B1(w2685) );
	ym3438_AON2222 g_2417 (.A2(w2749), .Z(w2825), .B2(w2756), .C2(w2553), .B1(w2741), .D1(w2824), .D2(w2552), .A1(w2572), .C1(w2823) );
	ym3438_NOT g_2418 (.A(w3909), .nZ(w2899) );
	ym3438_DLATCH_INV g_2419 (.nQ(w3909), .D(w2897), .C(w2545), .nC(w1150) );
	ym3438_FA g_2420 (.CO(w2863), .S(w2897), .CI(w2898), .A(w2602), .B(w2896) );
	ym3438_DLATCH_INV g_2421 (.nQ(w2896), .D(w2893), .C(w2546), .nC(w1149) );
	ym3438_AOI22 g_2422 (.A2(w2548), .A1(w2891), .Z(w2893), .B2(w2547), .B1(w2750) );
	ym3438_AON2222 g_2423 (.A2(w2756), .Z(w2891), .B2(w2823), .C2(w2553), .B1(w2741), .D1(w2889), .D2(w2552), .A1(w2572), .C1(w2824) );
	ym3438_NOT g_2424 (.A(w3903), .nZ(w2964) );
	ym3438_DLATCH_INV g_2425 (.nQ(w3903), .D(w2895), .C(w2545), .nC(w1150) );
	ym3438_FA g_2426 (.CO(w2898), .S(w2895), .CI(w2930), .A(w2602), .B(w2894) );
	ym3438_DLATCH_INV g_2427 (.nQ(w2894), .D(w2892), .C(w2546), .nC(w1149) );
	ym3438_AOI22 g_2428 (.A2(w2548), .A1(w2890), .Z(w2892), .B2(w2547), .B1(w2751) );
	ym3438_AON2222 g_2429 (.A2(w2823), .Z(w2890), .B2(w2824), .C2(w2553), .B1(w2741), .D1(w2888), .D2(w2552), .A1(w2572), .C1(w2889) );
	ym3438_NOT g_2430 (.A(w3908), .nZ(w2958) );
	ym3438_DLATCH_INV g_2431 (.nQ(w3908), .D(w2956), .C(w2545), .nC(w1150) );
	ym3438_FA g_2432 (.CO(w2930), .S(w2956), .CI(w2957), .A(w2602), .B(w2953) );
	ym3438_DLATCH_INV g_2433 (.nQ(w2953), .D(w2952), .C(w2546), .nC(w1149) );
	ym3438_AOI22 g_2434 (.A2(w2548), .A1(w2950), .Z(w2952), .B2(w2547), .B1(w2826) );
	ym3438_AON2222 g_2435 (.A2(w2824), .Z(w2950), .B2(w2889), .C2(w2553), .B1(w2741), .D1(w2929), .D2(w2552), .C1(w2888), .A1(w2572) );
	ym3438_NOT g_2436 (.A(w3902), .nZ(w3112) );
	ym3438_DLATCH_INV g_2437 (.nQ(w3902), .D(w2955), .C(w2545), .nC(w1150) );
	ym3438_FA g_2438 (.CO(w2957), .S(w2955), .CI(w3092), .A(w3091), .B(w2954) );
	ym3438_DLATCH_INV g_2439 (.nQ(w2954), .D(w2951), .C(w2546), .nC(w1149) );
	ym3438_AOI22 g_2440 (.A2(w2548), .A1(w2949), .Z(w2951), .B2(w2547), .B1(w2825) );
	ym3438_AON2222 g_2441 (.A2(w2889), .Z(w2949), .B2(w2888), .C2(w2553), .B1(w2741), .D1(1'b0), .D2(w2552), .A1(w2572), .C1(w2929) );
	ym3438_NOT g_2442 (.A(w3907), .nZ(w3106) );
	ym3438_DLATCH_INV g_2443 (.nQ(w3907), .D(w2995), .C(w2545), .nC(w1150) );
	ym3438_FA g_2444 (.CO(w3092), .S(w2995), .CI(w2994), .A(w3090), .B(w2993) );
	ym3438_DLATCH_INV g_2445 (.nQ(w2993), .D(w2990), .C(w2546), .nC(w1149) );
	ym3438_AOI22 g_2446 (.A2(w2548), .A1(w2988), .Z(w2990), .B2(w2547), .B1(w2891) );
	ym3438_AON22 g_2447 (.A2(w2553), .A1(w2812), .Z(w2636), .B2(w2552), .B1(w1143) );
	ym3438_AON22 g_2448 (.A2(w2553), .A1(1'b0), .Z(w2574), .B2(w2552), .B1(w2812) );
	ym3438_SR_BIT g_2449 (.Q(w3192), .D(w806), .nC1(w1150), .nC2(w1149), .C1(w2545), .C2(w2546) );
	ym3438_DLATCH_INV g_2450 (.nQ(w3969), .D(w3192), .C(w2545), .nC(w1150) );
	ym3438_AON222222 g_2451 (.A2(1'b0), .B1(w2615), .A1(1'b0), .Z(w3150), .C1(w2614), .C2(w3893), .D1(w2617), .D2(w2566), .E1(w3889), .E2(w3889), .F1(w2618), .F2(w2567) );
	ym3438_AON2222 g_2452 (.A2(w2567), .A1(w2567), .Z(w3123), .B2(w2618), .C1(w3893), .C2(w2617), .B1(w2566), .D1(w3891), .D2(w2614) );
	ym3438_AON222 g_2453 (.A2(w3891), .A1(w2617), .Z(w2560), .B2(w3893), .C1(w2566), .C2(w2566), .B1(w2618) );
	ym3438_AND g_2454 (.Z(w2604), .B(w3891), .A(w3891) );
	ym3438_NOT g_2455 (.A(w3967), .nZ(w2561) );
	ym3438_NOT g_2456 (.A(w2605), .nZ(w3967) );
	ym3438_SR_BIT g_2457 (.Q(w2613), .D(w232), .nC1(w1150), .nC2(w1149), .C1(w2545), .C2(w2546) );
	ym3438_SR_BIT g_2458 (.Q(w2564), .D(w335), .nC1(w1150), .nC2(w1149), .C1(w2545), .C2(w2546) );
	ym3438_AND g_2459 (.A(w215), .Z(w2369), .B(w3198) );
	ym3438_AND g_2460 (.A(w334), .Z(w1185), .B(w195) );
	ym3438_AON33 g_2461 (.A1(w334), .Z(w1184), .B2(w195), .A2(w194), .B1(w334), .A3(w26), .B3(w3199) );
	ym3438_AND g_2462 (.A(w1178), .Z(w1179), .B(w195) );
	ym3438_AND g_2463 (.A(w1178), .Z(w727), .B(w194) );
	ym3438_AND5 g_2464 (.A(w3204), .Z(w3198), .B(w3205), .C(w3210), .D(w3206), .E(w3207) );
	ym3438_AND5 g_2465 (.A(w3209), .Z(w2410), .B(w3208), .C(w4308), .D(w3206), .E(w3207) );
	ym3438_AND g_2466 (.A(w2216), .Z(w2317), .B(w3198) );
	ym3438_NOT g_2467 (.A(w2317), .nZ(w2316) );
	ym3438_SR_BIT g_2468 (.Q(w3203), .D(w2385), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24) );
	ym3438_SR_BIT g_2469 (.Q(w1183), .D(w3203), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24) );
	ym3438_SR_BIT g_2470 (.Q(w3202), .D(w185), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24) );
	ym3438_SR_BIT g_2471 (.Q(w1182), .D(w3202), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24) );
	ym3438_SR_BIT g_2472 (.Q(w3200), .D(w4013), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24) );
	ym3438_SR_BIT g_2473 (.Q(w1180), .D(w3200), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24) );
	ym3438_SR_BIT g_2474 (.Q(w3201), .D(w2384), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24) );
	ym3438_SR_BIT g_2475 (.Q(w1181), .D(w3201), .C1(w23), .C2(w22), .nC1(w25), .nC2(w24) );
	ym3438_NOT g_2476 (.A(w2369), .nZ(w2379) );
	ym3438_NOT g_2477 (.A(w26), .nZ(w3199) );
	ym3438_NOT g_2478 (.A(w195), .nZ(w194) );
	ym3438_NOT g_2479 (.A(w334), .nZ(w1178) );
	ym3438_COMP_STR g_2480 (.A(w2424), .Z(w2216), .nZ(w215) );
	ym3438_NOT g_2481 (.A(w2439), .nZ(w3215) );
	ym3438_AOI22 g_2482 (.A2(w2439), .B1(w2414), .A1(w3216), .Z(w3217), .B2(w3215) );
	ym3438_NOR g_2483 (.Z(w3218), .B(w1111), .A(w3217) );
	ym3438_SR_BIT g_2484 (.Q(w2414), .D(w3218), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_2485 (.A(w2439), .nZ(w3219) );
	ym3438_AOI22 g_2486 (.A2(w2439), .B1(w2423), .A1(w123), .Z(w3220), .B2(w3219) );
	ym3438_NOR g_2487 (.Z(w3221), .B(w1111), .A(w3220) );
	ym3438_SR_BIT g_2488 (.Q(w2423), .D(w3221), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_2489 (.A(w2439), .nZ(w3222) );
	ym3438_AOI22 g_2490 (.A2(w2439), .B1(w2422), .A1(w961), .Z(w3223), .B2(w3222) );
	ym3438_NOR g_2491 (.Z(w3224), .B(w1111), .A(w3223) );
	ym3438_SR_BIT g_2492 (.Q(w2422), .D(w3224), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_2493 (.A(w2439), .nZ(w3225) );
	ym3438_AOI22 g_2494 (.A2(w2439), .B1(w2421), .A1(w132), .Z(w3226), .B2(w3225) );
	ym3438_SR_BIT g_2496 (.Q(w2421), .D(w3227), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_2497 (.A(w2439), .nZ(w3228) );
	ym3438_AOI22 g_2498 (.A2(w2439), .B1(w2420), .A1(w960), .Z(w3229), .B2(w3228) );
	ym3438_NOR g_2499 (.Z(w3230), .B(w1111), .A(w3229) );
	ym3438_SR_BIT g_2500 (.Q(w2420), .D(w3230), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_2501 (.A(w2439), .nZ(w3231) );
	ym3438_AOI22 g_2502 (.A2(w2439), .B1(w2424), .A1(w959), .Z(w3232), .B2(w3231) );
	ym3438_SR_BIT g_2504 (.Q(w2424), .D(w3233), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_2505 (.A(w2439), .nZ(w3234) );
	ym3438_AOI22 g_2506 (.A2(w2439), .B1(w2413), .A1(w958), .Z(w3235), .B2(w3234) );
	ym3438_NOR g_2507 (.Z(w3236), .B(w1111), .A(w3235) );
	ym3438_SR_BIT g_2508 (.Q(w2413), .D(w3236), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_2509 (.A(w2439), .nZ(w3237) );
	ym3438_AOI22 g_2510 (.A2(w2439), .B1(w2412), .A1(w108), .Z(w3238), .B2(w3237) );
	ym3438_NOR g_2511 (.Z(w3239), .B(w1111), .A(w3238) );
	ym3438_SR_BIT g_2512 (.Q(w2412), .D(w3239), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_2513 (.A(w2439), .nZ(w3240) );
	ym3438_AOI22 g_2514 (.A2(w2439), .B1(w2411), .A1(w112), .Z(w3241), .B2(w3240) );
	ym3438_NOR g_2515 (.Z(w3242), .B(w1111), .A(w3241) );
	ym3438_SR_BIT g_2516 (.Q(w2411), .D(w3242), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_2517 (.A(w3250), .nZ(w340) );
	ym3438_NOT g_2518 (.A(w2447), .nZ(w3250) );
	ym3438_SR_BIT g_2519 (.Q(w2447), .D(w3251), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOR g_2520 (.Z(w3251), .B(w1111), .A(w3252) );
	ym3438_AOI22 g_2521 (.A2(w2437), .B1(w2447), .A1(w123), .Z(w3252), .B2(w3253) );
	ym3438_NOT g_2522 (.A(w2437), .nZ(w3253) );
	ym3438_NOT g_2523 (.A(w3254), .nZ(w329) );
	ym3438_NOT g_2524 (.A(w2446), .nZ(w3254) );
	ym3438_SR_BIT g_2525 (.Q(w2446), .D(w3255), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOR g_2526 (.Z(w3255), .B(w1111), .A(w3256) );
	ym3438_AOI22 g_2527 (.A2(w2437), .B1(w2446), .A1(w961), .Z(w3256), .B2(w3257) );
	ym3438_NOT g_2528 (.A(w2437), .nZ(w3257) );
	ym3438_NOT g_2529 (.A(w3258), .nZ(w330) );
	ym3438_NOT g_2530 (.A(w2445), .nZ(w3258) );
	ym3438_SR_BIT g_2531 (.Q(w2445), .D(w3259), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOR g_2532 (.Z(w3259), .B(w1111), .A(w3260) );
	ym3438_AOI22 g_2533 (.A2(w2437), .B1(w2445), .A1(w132), .Z(w3260), .B2(w3261) );
	ym3438_NOT g_2534 (.A(w2437), .nZ(w3261) );
	ym3438_NOT g_2535 (.A(w3262), .nZ(w331) );
	ym3438_NOT g_2536 (.A(w2444), .nZ(w3262) );
	ym3438_SR_BIT g_2537 (.Q(w2444), .D(w3263), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOR g_2538 (.Z(w3263), .B(w1111), .A(w3264) );
	ym3438_AOI22 g_2539 (.A2(w2437), .B1(w2444), .A1(w960), .Z(w3264), .B2(w3265) );
	ym3438_NOT g_2540 (.A(w2437), .nZ(w3265) );
	ym3438_NOT g_2541 (.A(w3266), .nZ(w338) );
	ym3438_NOT g_2542 (.A(w2443), .nZ(w3266) );
	ym3438_SR_BIT g_2543 (.Q(w2443), .D(w3267), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOR g_2544 (.Z(w3267), .B(w1111), .A(w3268) );
	ym3438_AOI22 g_2545 (.A2(w2437), .B1(w2443), .A1(w959), .Z(w3268), .B2(w3269) );
	ym3438_NOT g_2546 (.A(w2437), .nZ(w3269) );
	ym3438_NOT g_2547 (.A(w3270), .nZ(w337) );
	ym3438_SR_BIT g_2549 (.Q(w2442), .D(w3271), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOR g_2550 (.Z(w3271), .B(w1111), .A(w3272) );
	ym3438_AOI22 g_2551 (.A2(w2437), .B1(w2442), .A1(w958), .Z(w3272), .B2(w3273) );
	ym3438_NOT g_2552 (.A(w2437), .nZ(w3273) );
	ym3438_NOT g_2553 (.A(w3274), .nZ(w336) );
	ym3438_NOT g_2554 (.A(w2441), .nZ(w3274) );
	ym3438_SR_BIT g_2555 (.Q(w2441), .D(w3275), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOR g_2556 (.Z(w3275), .B(w1111), .A(w3276) );
	ym3438_AOI22 g_2557 (.A2(w2437), .B1(w2441), .A1(w108), .Z(w3276), .B2(w3277) );
	ym3438_NOT g_2558 (.A(w2437), .nZ(w3277) );
	ym3438_NOT g_2559 (.A(w3278), .nZ(w332) );
	ym3438_SR_BIT g_2561 (.Q(w2440), .D(w3279), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOR g_2562 (.Z(w3279), .B(w1111), .A(w3280) );
	ym3438_AOI22 g_2563 (.A2(w2437), .B1(w2440), .A1(w112), .Z(w3280), .B2(w3281) );
	ym3438_NOT g_2564 (.A(w2437), .nZ(w3281) );
	ym3438_NOT g_2565 (.A(w3282), .nZ(w2438) );
	ym3438_SR_BIT g_2566 (.Q(w3282), .D(w3283), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI21 g_2567 (.A1(w3284), .Z(w3283), .B(w2439), .A2(w2438) );
	ym3438_NOT g_2568 (.A(w1103), .nZ(w3284) );
	ym3438_NOT g_2569 (.A(w3285), .nZ(w2415) );
	ym3438_SR_BIT g_2570 (.Q(w3285), .D(w3286), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI21 g_2571 (.A1(w3287), .Z(w3286), .A2(w2415), .B(w2437) );
	ym3438_NOT g_2572 (.A(w1103), .nZ(w3287) );
	ym3438_AND g_2573 (.A(w2216), .Z(w2403), .B(w2410) );
	ym3438_AND5 g_2574 (.A(w3204), .Z(w203), .B(w3208), .C(w4308), .D(w3206), .E(w3207) );
	ym3438_AND5 g_2575 (.A(w3209), .Z(w145), .B(w3205), .C(w4308), .D(w3206), .E(w3207) );
	ym3438_AND5 g_2576 (.A(w3204), .Z(w211), .B(w3205), .C(w4308), .D(w3206), .E(w3207) );
	ym3438_AND5 g_2577 (.A(w3209), .Z(w143), .B(w3208), .C(w3210), .D(w167), .E(w3207) );
	ym3438_AND5 g_2578 (.A(w3204), .Z(w2215), .B(w3208), .C(w3210), .D(w167), .E(w3207) );
	ym3438_COMP_WE g_2579 (.A(w2423), .nZ(w3206), .Z(w167) );
	ym3438_COMP_WE g_2580 (.A(w2422), .nZ(w3210), .Z(w4308) );
	ym3438_COMP_WE g_2581 (.A(w2421), .nZ(w3208), .Z(w3205) );
	ym3438_COMP_WE g_2582 (.A(w2420), .nZ(w3209), .Z(w3204) );
	ym3438_AND g_2583 (.A(w2415), .Z(w3207), .B(w3211) );
	ym3438_XOR g_2584 (.A(w1176), .Z(w3212), .B(w2414) );
	ym3438_NOR4 g_2585 (.A(w3212), .Z(w3211), .B(w3213), .C(w3214), .D(w4309) );
	ym3438_XOR g_2586 (.A(w2413), .Z(w4309), .B(w1177) );
	ym3438_XOR g_2587 (.A(w2412), .Z(w3213), .B(w1007) );
	ym3438_XOR g_2588 (.A(w2411), .Z(w3214), .B(w988) );
	ym3438_AND g_2589 (.A(w2410), .Z(w2348), .B(w215) );
	ym3438_NOT g_2590 (.A(w2348), .nZ(w2347) );
	ym3438_NOT g_2591 (.A(w2403), .nZ(w2404) );
	ym3438_NOT g_2592 (.A(w120), .nZ(w3216) );
	ym3438_OR4 g_2593 (.A(w960), .Z(w3243), .B(w961), .D(w123), .C(w132) );
	ym3438_NAND g_2594 (.A(w3243), .Z(w3244), .B(w1103) );
	ym3438_NOT g_2595 (.A(w3244), .nZ(w2439) );
	ym3438_NAND g_2596 (.A(w2438), .Z(w3245), .B(w121) );
	ym3438_NOT g_2597 (.A(w3245), .nZ(w2437) );
	ym3438_XOR g_2598 (.A(w2414), .Z(w2419), .B(w1176) );
	ym3438_XOR g_2599 (.A(w2412), .Z(w3246), .B(w1007) );
	ym3438_XOR g_2600 (.A(w2411), .Z(w3247), .B(w988) );
	ym3438_NOR3 g_2601 (.C(w3247), .A(w2419), .Z(w3248), .B(w3246) );
	ym3438_AND g_2602 (.A(w3248), .Z(w3249), .B(w2415) );
	ym3438_COMP_WE g_2603 (.A(w2413), .nZ(w2435), .Z(w2434) );
	ym3438_COMP_WE g_2604 (.A(w2424), .nZ(w2433), .Z(w2436) );
	ym3438_COMP_WE g_2605 (.A(w2420), .nZ(w2432), .Z(w2431) );
	ym3438_NOT g_2606 (.A(w2422), .nZ(w2418) );
	ym3438_NAND7 g_2607 (.A(w3249), .Z(w1114), .B(w2423), .G(w2435), .D(w2421), .F(w2433), .C(w2418), .E(w2432) );
	ym3438_NAND7 g_2608 (.A(w3249), .Z(w2430), .B(w2423), .G(w2434), .D(w2421), .F(w2433), .C(w2418), .E(w2432) );
	ym3438_NAND7 g_2609 (.A(w3249), .Z(w1113), .B(w2423), .G(w2435), .D(w2421), .F(w2432), .C(w2418), .E(w2436) );
	ym3438_NAND7 g_2610 (.A(w3249), .Z(w2429), .B(w2423), .G(w2434), .D(w2421), .F(w2436), .C(w2418), .E(w2432) );
	ym3438_NAND7 g_2611 (.A(w3249), .Z(w2428), .B(w2423), .G(w2435), .D(w2421), .F(w2433), .C(w2418), .E(w2431) );
	ym3438_NAND7 g_2612 (.A(w3249), .Z(w2427), .B(w2423), .G(w2434), .D(w2421), .F(w2433), .C(w2418), .E(w2431) );
	ym3438_NOR g_2613 (.Z(w3314), .B(w1111), .A(w3289) );
	ym3438_SR_BIT g_2614 (.Q(w3315), .D(w3314), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2615 (.Q(w3316), .D(w3315), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2616 (.Q(w3317), .D(w3316), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2617 (.Q(w3318), .D(w3317), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2618 (.Q(w2463), .D(w3318), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2619 (.Q(w2462), .D(w2463), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2620 (.A2(w2462), .B1(w340), .A1(w3288), .Z(w3289), .B2(w1112) );
	ym3438_NOR g_2621 (.Z(w3327), .B(w1111), .A(w3324) );
	ym3438_SR_BIT g_2622 (.Q(w4331), .D(w3327), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2623 (.Q(w3329), .D(w4331), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2624 (.Q(w3331), .D(w3329), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2625 (.Q(w3334), .D(w3331), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2626 (.Q(w2461), .D(w3334), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2627 (.Q(w2459), .D(w2461), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2628 (.A2(w2459), .B1(w329), .A1(w3288), .Z(w3324), .B2(w1112) );
	ym3438_NOR g_2629 (.Z(w3339), .B(w1111), .A(w3338) );
	ym3438_SR_BIT g_2630 (.Q(w3342), .D(w3339), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2631 (.Q(w3343), .D(w3342), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2632 (.Q(w3345), .D(w3343), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2633 (.Q(w3347), .D(w3345), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2634 (.Q(w2460), .D(w3347), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2635 (.Q(w2458), .D(w2460), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2636 (.A2(w2458), .B1(w330), .A1(w3288), .Z(w3338), .B2(w1112) );
	ym3438_NOR g_2637 (.Z(w3350), .B(w1111), .A(w3349) );
	ym3438_SR_BIT g_2638 (.Q(w3353), .D(w3350), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2639 (.Q(w3355), .D(w3353), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2640 (.Q(w3357), .D(w3355), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2641 (.Q(w3359), .D(w3357), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2642 (.Q(w2457), .D(w3359), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2643 (.Q(w2456), .D(w2457), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2644 (.A2(w2456), .B1(w331), .A1(w3288), .Z(w3349), .B2(w1112) );
	ym3438_NOR g_2645 (.Z(w3364), .B(w1111), .A(w3362) );
	ym3438_SR_BIT g_2646 (.Q(w3366), .D(w3364), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2647 (.Q(w3368), .D(w3366), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2648 (.Q(w3370), .D(w3368), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2649 (.Q(w3372), .D(w3370), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2650 (.Q(w2455), .D(w3372), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2651 (.Q(w2454), .D(w2455), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2652 (.A2(w2454), .B1(w338), .A1(w3288), .Z(w3362), .B2(w1112) );
	ym3438_NOR g_2653 (.Z(w3377), .B(w1111), .A(w3376) );
	ym3438_SR_BIT g_2654 (.Q(w3379), .D(w3377), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2655 (.Q(w3380), .D(w3379), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2656 (.Q(w3383), .D(w3380), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2657 (.Q(w3385), .D(w3383), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2658 (.Q(w2453), .D(w3385), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2659 (.Q(w2452), .D(w2453), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2660 (.A2(w2452), .B1(w337), .A1(w3288), .Z(w3376), .B2(w1112) );
	ym3438_NOR g_2661 (.Z(w3312), .B(w1111), .A(w3388) );
	ym3438_SR_BIT g_2662 (.Q(w3310), .D(w3312), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2663 (.Q(w3308), .D(w3310), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2664 (.Q(w3306), .D(w3308), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2665 (.Q(w3304), .D(w3306), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2666 (.Q(w2451), .D(w3304), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2667 (.Q(w2449), .D(w2451), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2668 (.A2(w2449), .B1(w336), .A1(w3288), .Z(w3388), .B2(w1112) );
	ym3438_NOR g_2669 (.Z(w3301), .B(w1111), .A(w3390) );
	ym3438_SR_BIT g_2670 (.Q(w3300), .D(w3301), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2671 (.Q(w3299), .D(w3300), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2672 (.Q(w3293), .D(w3299), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2673 (.Q(w3292), .D(w3293), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2674 (.Q(w2450), .D(w3292), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2675 (.Q(w2448), .D(w2450), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2676 (.A2(w2448), .B1(w332), .A1(w3288), .Z(w3390), .B2(w1112) );
	ym3438_NOR g_2677 (.Z(w3319), .B(w1111), .A(w3291) );
	ym3438_SR_BIT g_2678 (.Q(w3320), .D(w3319), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2679 (.Q(w3321), .D(w3320), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2680 (.Q(w3322), .D(w3321), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2681 (.Q(w3323), .D(w3322), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2682 (.Q(w2472), .D(w3323), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2683 (.Q(w2470), .D(w2472), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2684 (.A2(w2470), .B1(w340), .A1(w3290), .Z(w3291), .B2(w1115) );
	ym3438_NOR g_2685 (.Z(w3326), .B(w1111), .A(w3325) );
	ym3438_SR_BIT g_2686 (.Q(w3328), .D(w3326), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2687 (.Q(w3330), .D(w3328), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2688 (.Q(w3332), .D(w3330), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2689 (.Q(w3333), .D(w3332), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2690 (.Q(w3335), .D(w3333), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2691 (.Q(w2471), .D(w3335), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2692 (.A2(w2471), .B1(w329), .A1(w3290), .Z(w3325), .B2(w1115) );
	ym3438_NOR g_2693 (.Z(w3341), .B(w1111), .A(w3340) );
	ym3438_SR_BIT g_2694 (.Q(w3337), .D(w3341), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2695 (.Q(w3344), .D(w3337), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2696 (.Q(w3346), .D(w3344), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2697 (.Q(w3348), .D(w3346), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2698 (.Q(w3336), .D(w3348), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2699 (.Q(w2469), .D(w3336), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2700 (.A2(w2469), .B1(w330), .A1(w3290), .Z(w3340), .B2(w1115) );
	ym3438_NOR g_2701 (.Z(w3417), .B(w1111), .A(w3416) );
	ym3438_SR_BIT g_2702 (.Q(w2503), .D(w3417), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2703 (.Q(w3420), .D(w2503), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2704 (.Q(w3423), .D(w3420), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2705 (.Q(w3424), .D(w3423), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2706 (.Q(w3398), .D(w3424), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2707 (.Q(w2502), .D(w3398), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2708 (.A2(w2502), .B1(w2524), .A1(w3415), .Z(w3416), .B2(w1115) );
	ym3438_NOR g_2709 (.Z(w3418), .B(w1111), .A(w3471) );
	ym3438_SR_BIT g_2710 (.Q(w3419), .D(w3418), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2711 (.Q(w3421), .D(w3419), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2712 (.Q(w3422), .D(w3421), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2713 (.Q(w3425), .D(w3422), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2714 (.Q(w2504), .D(w3425), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2715 (.Q(w2510), .D(w2504), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2716 (.A2(w2510), .B1(w2523), .A1(w3470), .Z(w3471), .B2(w1112) );
	ym3438_NOR g_2717 (.Z(w3426), .B(w1111), .A(w3472) );
	ym3438_SR_BIT g_2718 (.Q(w2500), .D(w3426), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2719 (.Q(w3429), .D(w2500), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2720 (.Q(w3431), .D(w3429), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2721 (.Q(w3433), .D(w3431), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2722 (.Q(w3400), .D(w3433), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2723 (.Q(w2499), .D(w3400), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2724 (.A2(w2499), .B1(w2522), .A1(w3415), .Z(w3472), .B2(w1115) );
	ym3438_NOR g_2725 (.Z(w3435), .B(w1111), .A(w3473) );
	ym3438_SR_BIT g_2726 (.Q(w2497), .D(w3435), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2727 (.Q(w3438), .D(w2497), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2728 (.Q(w3440), .D(w3438), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2729 (.Q(w3442), .D(w3440), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2730 (.Q(w3401), .D(w3442), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2731 (.Q(w2496), .D(w3401), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2732 (.A2(w2496), .B1(w2520), .A1(w3415), .Z(w3473), .B2(w1115) );
	ym3438_NOR g_2733 (.Z(w3444), .B(w1111), .A(w3475) );
	ym3438_SR_BIT g_2734 (.Q(w2494), .D(w3444), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2735 (.Q(w3447), .D(w2494), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2736 (.Q(w3449), .D(w3447), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2737 (.Q(w3451), .D(w3449), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2738 (.Q(w3402), .D(w3451), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2739 (.Q(w2493), .D(w3402), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2740 (.A2(w2493), .B1(w2518), .A1(w3415), .Z(w3475), .B2(w1115) );
	ym3438_NOR g_2741 (.Z(w3453), .B(w1111), .A(w3478) );
	ym3438_SR_BIT g_2742 (.Q(w2491), .D(w3453), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2743 (.Q(w3456), .D(w2491), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2744 (.Q(w3458), .D(w3456), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2745 (.Q(w3460), .D(w3458), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2746 (.Q(w3408), .D(w3460), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2747 (.Q(w2490), .D(w3408), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2748 (.A2(w2490), .B1(w2516), .A1(w3415), .Z(w3478), .B2(w1115) );
	ym3438_NOR g_2749 (.Z(w4336), .B(w1111), .A(w3479) );
	ym3438_SR_BIT g_2750 (.Q(w3410), .D(w4336), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2751 (.Q(w3464), .D(w3410), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2752 (.Q(w3466), .D(w3464), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2753 (.Q(w3468), .D(w3466), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2754 (.Q(w3409), .D(w3468), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2755 (.Q(w2487), .D(w3409), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2756 (.A2(w2487), .B1(w2514), .A1(w3415), .Z(w3479), .B2(w1115) );
	ym3438_NOR g_2757 (.Z(w3427), .B(w1111), .A(w4337) );
	ym3438_SR_BIT g_2758 (.Q(w3428), .D(w3427), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2759 (.Q(w3430), .D(w3428), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2760 (.Q(w3432), .D(w3430), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2761 (.Q(w3434), .D(w3432), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2762 (.Q(w2501), .D(w3434), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2763 (.Q(w2509), .D(w2501), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2764 (.A2(w2509), .B1(w2521), .A1(w3470), .Z(w4337), .B2(w1112) );
	ym3438_NOR g_2765 (.Z(w3436), .B(w1111), .A(w3474) );
	ym3438_SR_BIT g_2766 (.Q(w3437), .D(w3436), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2767 (.Q(w3439), .D(w3437), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2768 (.Q(w3441), .D(w3439), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2769 (.Q(w3443), .D(w3441), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2770 (.Q(w2498), .D(w3443), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2771 (.Q(w2508), .D(w2498), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2772 (.A2(w2508), .B1(w2519), .A1(w3470), .Z(w3474), .B2(w1112) );
	ym3438_NOR g_2773 (.Z(w3445), .B(w1111), .A(w3476) );
	ym3438_SR_BIT g_2774 (.Q(w3446), .D(w3445), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2775 (.Q(w3448), .D(w3446), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2776 (.Q(w3450), .D(w3448), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2777 (.Q(w3452), .D(w3450), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2778 (.Q(w2495), .D(w3452), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2779 (.Q(w2507), .D(w2495), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2780 (.A2(w2507), .B1(w2517), .A1(w3470), .Z(w3476), .B2(w1112) );
	ym3438_NOR g_2781 (.Z(w3454), .B(w1111), .A(w3477) );
	ym3438_SR_BIT g_2782 (.Q(w3455), .D(w3454), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2783 (.Q(w3457), .D(w3455), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2784 (.Q(w3459), .D(w3457), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2785 (.Q(w3461), .D(w3459), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2786 (.Q(w2492), .D(w3461), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2787 (.Q(w2506), .D(w2492), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2788 (.A2(w2506), .B1(w2515), .A1(w3470), .Z(w3477), .B2(w1112) );
	ym3438_NOR g_2789 (.Z(w3462), .B(w1111), .A(w3480) );
	ym3438_SR_BIT g_2790 (.Q(w3463), .D(w3462), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2791 (.Q(w3465), .D(w3463), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2792 (.Q(w3467), .D(w3465), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2793 (.Q(w3469), .D(w3467), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2794 (.Q(w2488), .D(w3469), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2795 (.Q(w2505), .D(w2488), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2796 (.A2(w2505), .B1(w2513), .A1(w3470), .Z(w3480), .B2(w1112) );
	ym3438_NOR g_2797 (.Z(w3352), .B(w1111), .A(w3351) );
	ym3438_SR_BIT g_2798 (.Q(w3354), .D(w3352), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2799 (.Q(w3356), .D(w3354), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2800 (.Q(w3358), .D(w3356), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2801 (.Q(w3360), .D(w3358), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2802 (.Q(w3361), .D(w3360), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2803 (.Q(w2468), .D(w3361), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2804 (.A2(w2468), .B1(w331), .A1(w3290), .Z(w3351), .B2(w1115) );
	ym3438_NOR g_2805 (.Z(w3365), .B(w1111), .A(w3363) );
	ym3438_SR_BIT g_2806 (.Q(w3367), .D(w3365), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2807 (.Q(w3369), .D(w3367), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2808 (.Q(w3371), .D(w3369), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2809 (.Q(w3373), .D(w3371), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2810 (.Q(w3374), .D(w3373), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2811 (.Q(w2467), .D(w3374), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2812 (.A2(w2467), .B1(w338), .A1(w3290), .Z(w3363), .B2(w1115) );
	ym3438_NOR g_2813 (.Z(w3378), .B(w1111), .A(w3375) );
	ym3438_SR_BIT g_2814 (.Q(w3381), .D(w3378), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2815 (.Q(w3382), .D(w3381), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2816 (.Q(w3384), .D(w3382), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2817 (.Q(w3386), .D(w3384), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2818 (.Q(w3387), .D(w3386), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2819 (.Q(w2466), .D(w3387), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2820 (.A2(w2466), .B1(w337), .A1(w3290), .Z(w3375), .B2(w1115) );
	ym3438_NOR g_2821 (.Z(w3313), .B(w1111), .A(w3389) );
	ym3438_SR_BIT g_2822 (.Q(w3311), .D(w3313), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2823 (.Q(w3309), .D(w3311), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2824 (.Q(w3307), .D(w3309), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2825 (.Q(w3305), .D(w3307), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2826 (.Q(w3303), .D(w3305), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2827 (.Q(w2465), .D(w3303), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2828 (.A2(w2465), .B1(w336), .A1(w3290), .Z(w3389), .B2(w1115) );
	ym3438_NOR g_2829 (.Z(w3302), .B(w1111), .A(w3391) );
	ym3438_SR_BIT g_2830 (.Q(w3297), .D(w3302), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2831 (.Q(w3296), .D(w3297), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2832 (.Q(w3295), .D(w3296), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2833 (.Q(w3294), .D(w3295), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2834 (.Q(w3298), .D(w3294), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2835 (.Q(w2464), .D(w3298), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2836 (.A2(w2464), .B1(w332), .A1(w3290), .Z(w3391), .B2(w1115) );
	ym3438_NOR g_2837 (.Z(w3587), .B(w1111), .A(w3588) );
	ym3438_SR_BIT g_2838 (.Q(w3530), .D(w3587), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2839 (.Q(w3586), .D(w3530), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2840 (.Q(w3585), .D(w3586), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2841 (.Q(w3584), .D(w3585), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2842 (.Q(w3583), .D(w3584), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2843 (.Q(w2530), .D(w3583), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2844 (.A2(w2530), .B1(w330), .A1(w3536), .Z(w3588), .B2(w1116) );
	ym3438_NOR g_2845 (.Z(w3593), .B(w1111), .A(w3589) );
	ym3438_SR_BIT g_2846 (.Q(w3594), .D(w3593), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2847 (.Q(w3595), .D(w3594), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2848 (.Q(w3596), .D(w3595), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2849 (.Q(w3597), .D(w3596), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2850 (.Q(w3529), .D(w3597), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2851 (.Q(w3590), .D(w3529), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2852 (.A2(w3590), .B1(w3591), .A1(w3537), .Z(w3589), .B2(w1117) );
	ym3438_NOR g_2853 (.Z(w3580), .B(w1111), .A(w3581) );
	ym3438_SR_BIT g_2854 (.Q(w3531), .D(w3580), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2855 (.Q(w3579), .D(w3531), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2856 (.Q(w3578), .D(w3579), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2857 (.Q(w3577), .D(w3578), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2858 (.Q(w3576), .D(w3577), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2859 (.Q(w2532), .D(w3576), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2860 (.A2(w2532), .B1(w331), .A1(w3536), .Z(w3581), .B2(w1116) );
	ym3438_NOR g_2861 (.Z(w3598), .B(w1111), .A(w3582) );
	ym3438_SR_BIT g_2862 (.Q(w3599), .D(w3598), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2863 (.Q(w3600), .D(w3599), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2864 (.Q(w3601), .D(w3600), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2865 (.Q(w3602), .D(w3601), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2866 (.Q(w3592), .D(w3602), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2867 (.Q(w3575), .D(w3592), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2868 (.A2(w3575), .B1(w2531), .A1(w3537), .Z(w3582), .B2(w1117) );
	ym3438_NOR g_2869 (.Z(w3572), .B(w1111), .A(w3573) );
	ym3438_SR_BIT g_2870 (.Q(w3532), .D(w3572), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2871 (.Q(w3571), .D(w3532), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2872 (.Q(w3570), .D(w3571), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2873 (.Q(w4340), .D(w3570), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2874 (.Q(w3569), .D(w4340), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2875 (.Q(w2533), .D(w3569), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2876 (.A2(w2533), .B1(w338), .A1(w3536), .Z(w3573), .B2(w1116) );
	ym3438_NOR g_2877 (.Z(w3603), .B(w1111), .A(w3574) );
	ym3438_SR_BIT g_2878 (.Q(w3604), .D(w3603), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2879 (.Q(w3605), .D(w3604), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2880 (.Q(w3606), .D(w3605), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2881 (.Q(w3607), .D(w3606), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2882 (.Q(w3608), .D(w3607), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2883 (.Q(w3543), .D(w3608), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2884 (.A2(w3543), .B1(w330), .A1(w3537), .Z(w3574), .B2(w1117) );
	ym3438_NOR g_2885 (.Z(w3566), .B(w1111), .A(w3567) );
	ym3438_SR_BIT g_2886 (.Q(w3565), .D(w3566), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2887 (.Q(w3564), .D(w3565), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2888 (.Q(w3563), .D(w3564), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2889 (.Q(w3562), .D(w3563), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2890 (.Q(w3561), .D(w3562), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2891 (.Q(w3533), .D(w3561), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2892 (.A2(w3533), .B1(w337), .A1(w3536), .Z(w3567), .B2(w1116) );
	ym3438_NOR g_2893 (.Z(w3609), .B(w1111), .A(w3568) );
	ym3438_SR_BIT g_2894 (.Q(w3610), .D(w3609), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2895 (.Q(w3611), .D(w3610), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2896 (.Q(w3612), .D(w3611), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2897 (.Q(w3613), .D(w3612), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2898 (.Q(w3614), .D(w3613), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2899 (.Q(w2999), .D(w3614), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2900 (.A2(w2999), .B1(w331), .A1(w3537), .Z(w3568), .B2(w1117) );
	ym3438_NOR g_2901 (.Z(w3558), .B(w1111), .A(w4341) );
	ym3438_SR_BIT g_2902 (.Q(w3557), .D(w3558), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2903 (.Q(w3556), .D(w3557), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2904 (.Q(w3555), .D(w3556), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2905 (.Q(w3554), .D(w3555), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2906 (.Q(w3553), .D(w3554), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2907 (.Q(w3534), .D(w3553), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2908 (.A2(w3534), .B1(w336), .A1(w3536), .Z(w4341), .B2(w1116) );
	ym3438_NOR g_2909 (.Z(w3560), .B(w1111), .A(w3559) );
	ym3438_SR_BIT g_2910 (.Q(w3615), .D(w3560), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2911 (.Q(w3616), .D(w3615), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2912 (.Q(w3617), .D(w3616), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2913 (.Q(w3618), .D(w3617), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2914 (.Q(w3619), .D(w3618), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2915 (.Q(w2998), .D(w3619), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2916 (.A2(w2998), .B1(w337), .A1(w3537), .Z(w3559), .B2(w1117) );
	ym3438_NOR g_2917 (.Z(w3550), .B(w1111), .A(w3551) );
	ym3438_SR_BIT g_2918 (.Q(w3549), .D(w3550), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2919 (.Q(w3547), .D(w3549), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2920 (.Q(w3548), .D(w3547), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2921 (.Q(w3546), .D(w3548), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2922 (.Q(w3545), .D(w3546), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2923 (.Q(w3535), .D(w3545), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2924 (.A2(w3535), .B1(w332), .A1(w3536), .Z(w3551), .B2(w1116) );
	ym3438_NOR g_2925 (.Z(w3620), .B(w1111), .A(w3552) );
	ym3438_SR_BIT g_2926 (.Q(w3621), .D(w3620), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2927 (.Q(w3622), .D(w3621), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2928 (.Q(w3623), .D(w3622), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2929 (.Q(w3624), .D(w3623), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2930 (.Q(w3625), .D(w3624), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_2931 (.Q(w2997), .D(w3625), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AOI22 g_2932 (.A2(w2997), .B1(w336), .A1(w3537), .Z(w3552), .B2(w1117) );
	ym3438_AON2222 g_2933 (.A2(w2470), .B1(w3320), .A1(w3396), .Z(w3394), .B2(w3395), .C2(w2472), .D1(w2463), .C1(w3393), .D2(w3392) );
	ym3438_AON2222 g_2934 (.A2(w2502), .B1(w2503), .A1(w3396), .Z(w1133), .B2(w3395), .C2(w3398), .D1(w2504), .C1(w3393), .D2(w3392) );
	ym3438_AON2222 g_2935 (.A2(w2471), .B1(w3328), .A1(w3396), .Z(w2473), .B2(w3395), .C2(w3335), .D1(w2461), .C1(w3393), .D2(w3392) );
	ym3438_SR_BIT g_2936 (.Q(w3397), .D(w3394), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_COMP_STR g_2937 (.A(w3397), .Z(w1121) );
	ym3438_SR_BIT g_2938 (.Q(w3399), .D(w2473), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_COMP_STR g_2939 (.A(w3399), .Z(w1122) );
	ym3438_AON2222 g_2940 (.A2(w2499), .B1(w2500), .A1(w3396), .Z(w1132), .B2(w3395), .D1(w2501), .C1(w3393), .D2(w3392), .C2(w3400) );
	ym3438_COMP_STR g_2941 (.A(w2474), .Z(w1123) );
	ym3438_SR_BIT g_2942 (.Q(w2474), .D(w2475), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AON2222 g_2943 (.A2(w2469), .B1(w3337), .A1(w3396), .Z(w2475), .B2(w3395), .C2(w3336), .D1(w2460), .C1(w3393), .D2(w3392) );
	ym3438_AON2222 g_2944 (.A2(w2496), .B1(w2497), .A1(w3396), .Z(w1131), .B2(w3395), .D1(w2498), .C1(w3393), .D2(w3392), .C2(w3401) );
	ym3438_COMP_STR g_2945 (.A(w2476), .Z(w1124) );
	ym3438_SR_BIT g_2946 (.Q(w2476), .D(w2477), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AON2222 g_2947 (.A2(w2457), .B1(w3361), .A1(w3392), .Z(w2477), .B2(w3393), .C2(w3354), .D1(w2468), .C1(w3395), .D2(w3396) );
	ym3438_AOI2222 g_2948 (.A2(w2493), .B1(w2494), .A1(w3396), .Z(w3403), .B2(w3395), .C2(w3402), .D1(w2495), .C1(w3393), .D2(w3392) );
	ym3438_NOT g_2949 (.A(w3403), .nZ(w1130) );
	ym3438_SR_BIT g_2950 (.Q(w3404), .D(w1130), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_COMP_STR g_2951 (.A(w3404), .Z(w1118) );
	ym3438_COMP_STR g_2952 (.A(w2478), .Z(w1125) );
	ym3438_SR_BIT g_2953 (.Q(w2478), .D(w2479), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AON2222 g_2954 (.A2(w2467), .B1(w3367), .A1(w3396), .Z(w2479), .B2(w3395), .C2(w3374), .D1(w2455), .C1(w3393), .D2(w3392) );
	ym3438_COMP_STR g_2955 (.A(w2480), .Z(w1119) );
	ym3438_SR_BIT g_2956 (.Q(w2480), .D(w2485), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AON2222 g_2957 (.A2(w2490), .B1(w2491), .A1(w3396), .Z(w2485), .B2(w3395), .D1(w2492), .C1(w3393), .D2(w3392), .C2(w3408) );
	ym3438_COMP_STR g_2958 (.A(w3405), .Z(w1126) );
	ym3438_SR_BIT g_2959 (.Q(w3405), .D(w2489), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_AON2222 g_2960 (.A2(w2466), .B1(w3381), .A1(w3396), .Z(w2489), .B2(w3395), .C2(w3387), .D1(w2453), .C1(w3393), .D2(w3392) );
	ym3438_AON2222 g_2961 (.A2(w2487), .B1(w3410), .A1(w3396), .Z(w2484), .B2(w3395), .D1(w2488), .C1(w3393), .D2(w3392), .C2(w3409) );
	ym3438_SR_BIT g_2962 (.Q(w3406), .D(w2484), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_COMP_STR g_2963 (.A(w3406), .Z(w1120) );
	ym3438_AON2222 g_2964 (.A2(w2465), .B1(w3311), .A1(w3396), .Z(w2486), .B2(w3395), .C2(w3303), .D1(w2451), .C1(w3393), .D2(w3392) );
	ym3438_SR_BIT g_2965 (.Q(w3407), .D(w2486), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_COMP_STR g_2966 (.A(w3407), .Z(w1127) );
	ym3438_OR3 g_2967 (.Z(w3411), .B(w2485), .A(w2484), .C(w3394) );
	ym3438_AND g_2968 (.Z(w3412), .B(w1130), .A(w3411) );
	ym3438_OR g_2969 (.Z(w1129), .B(w3413), .A(w3412) );
	ym3438_AND4 g_2970 (.Z(w3413), .B(w2485), .A(w3394), .C(w2484), .D(w3414) );
	ym3438_NOT g_2971 (.A(w1130), .nZ(w3414) );
	ym3438_AON2222 g_2972 (.A2(w2464), .B1(w3297), .A1(w3396), .Z(w2482), .B2(w3395), .C2(w3298), .D1(w2450), .C1(w3393), .D2(w3392) );
	ym3438_SR_BIT g_2973 (.Q(w2481), .D(w2482), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_COMP_STR g_2974 (.A(w2481), .Z(w1128) );
	ym3438_NOT g_2975 (.A(w214), .nZ(w1111) );
	ym3438_NOT g_2976 (.A(w1115), .nZ(w3415) );
	ym3438_NAND3 g_2977 (.Z(w3484), .B(w4194), .A(w1162), .C(w2483) );
	ym3438_NAND3 g_2978 (.Z(w3483), .B(w1162), .A(w4193), .C(w2483) );
	ym3438_NAND3 g_2979 (.Z(w3482), .B(w2483), .A(w3481), .C(w1162) );
	ym3438_AND g_2980 (.Z(w2483), .B(w3486), .A(w988) );
	ym3438_NOR g_2981 (.Z(w3486), .B(w1176), .A(w1007) );
	ym3438_NOT g_2982 (.A(w3485), .nZ(w3392) );
	ym3438_NOT g_2983 (.A(w3482), .nZ(w3396) );
	ym3438_NOT g_2984 (.A(w3483), .nZ(w3395) );
	ym3438_NOT g_2985 (.A(w3484), .nZ(w3393) );
	ym3438_AND g_2986 (.Z(w4194), .B(w2512), .A(w341) );
	ym3438_AND g_2987 (.Z(w4193), .B(w1177), .A(w2511) );
	ym3438_AND g_2988 (.Z(w3481), .B(w2512), .A(w2511) );
	ym3438_NAND3 g_2989 (.Z(w3485), .B(w3483), .A(w3484), .C(w3482) );
	ym3438_NOT g_2990 (.A(w1177), .nZ(w2512) );
	ym3438_NOT g_2991 (.A(w341), .nZ(w2511) );
	ym3438_NOT g_2992 (.A(w1112), .nZ(w3470) );
	ym3438_NOT g_2993 (.A(w217), .nZ(w3487) );
	ym3438_NOT g_2994 (.A(w212), .nZ(w3488) );
	ym3438_NOT g_2995 (.A(w216), .nZ(w3489) );
	ym3438_NOT g_2996 (.A(w1114), .nZ(w1112) );
	ym3438_NOT g_2997 (.A(w1113), .nZ(w1115) );
	ym3438_NOT g_2998 (.A(w213), .nZ(w3490) );
	ym3438_NOT g_2999 (.A(w3487), .nZ(w2416) );
	ym3438_NOT g_3000 (.A(w3488), .nZ(w2417) );
	ym3438_NOT g_3001 (.A(w3489), .nZ(w2426) );
	ym3438_NOT g_3002 (.A(w3490), .nZ(w2425) );
	ym3438_NOT g_3003 (.A(w2429), .nZ(w3491) );
	ym3438_NOT g_3004 (.A(w2430), .nZ(w3496) );
	ym3438_NOT g_3005 (.A(w2428), .nZ(w1116) );
	ym3438_NOT g_3006 (.A(w2427), .nZ(w1117) );
	ym3438_NOT g_3007 (.A(w3491), .nZ(w3492) );
	ym3438_AOI22 g_3008 (.A2(w3491), .B1(w2524), .A1(w330), .Z(w3493), .B2(w3492) );
	ym3438_NOR g_3009 (.Z(w3494), .B(w1111), .A(w3493) );
	ym3438_SR_BIT g_3010 (.Q(w2524), .D(w3494), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_3011 (.A(w3496), .nZ(w3495) );
	ym3438_AOI22 g_3012 (.A2(w3496), .B1(w2523), .A1(w330), .Z(w3497), .B2(w3495) );
	ym3438_NOR g_3013 (.Z(w3498), .B(w1111), .A(w3497) );
	ym3438_SR_BIT g_3014 (.Q(w2523), .D(w3498), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_3015 (.A(w3491), .nZ(w3499) );
	ym3438_AOI22 g_3016 (.A2(w3491), .B1(w2522), .A1(w331), .Z(w3500), .B2(w3499) );
	ym3438_NOR g_3017 (.Z(w3501), .B(w1111), .A(w3500) );
	ym3438_SR_BIT g_3018 (.Q(w2522), .D(w3501), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_3019 (.A(w3496), .nZ(w3502) );
	ym3438_AOI22 g_3020 (.A2(w3496), .B1(w2521), .A1(w331), .Z(w3503), .B2(w3502) );
	ym3438_NOR g_3021 (.Z(w3504), .B(w1111), .A(w3503) );
	ym3438_SR_BIT g_3022 (.Q(w2521), .D(w3504), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_3023 (.A(w3491), .nZ(w3505) );
	ym3438_AOI22 g_3024 (.A2(w3491), .B1(w2520), .A1(w338), .Z(w3506), .B2(w3505) );
	ym3438_NOR g_3025 (.Z(w3507), .B(w1111), .A(w3506) );
	ym3438_SR_BIT g_3026 (.Q(w2520), .D(w3507), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_3027 (.A(w3496), .nZ(w3508) );
	ym3438_AOI22 g_3028 (.A2(w3496), .B1(w2519), .A1(w338), .Z(w3509), .B2(w3508) );
	ym3438_NOR g_3029 (.Z(w3510), .B(w1111), .A(w3509) );
	ym3438_SR_BIT g_3030 (.Q(w2519), .D(w3510), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_3031 (.A(w3491), .nZ(w3511) );
	ym3438_AOI22 g_3032 (.A2(w3491), .B1(w2518), .A1(w337), .Z(w3512), .B2(w3511) );
	ym3438_NOR g_3033 (.Z(w3513), .B(w1111), .A(w3512) );
	ym3438_SR_BIT g_3034 (.Q(w2518), .D(w3513), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_3035 (.A(w3496), .nZ(w3514) );
	ym3438_AOI22 g_3036 (.A2(w3496), .B1(w2517), .A1(w337), .Z(w3515), .B2(w3514) );
	ym3438_NOR g_3037 (.Z(w3516), .B(w1111), .A(w3515) );
	ym3438_SR_BIT g_3038 (.Q(w2517), .D(w3516), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_3039 (.A(w3491), .nZ(w3517) );
	ym3438_AOI22 g_3040 (.A2(w3491), .B1(w2516), .A1(w336), .Z(w3518), .B2(w3517) );
	ym3438_NOR g_3041 (.Z(w3519), .B(w1111), .A(w3518) );
	ym3438_SR_BIT g_3042 (.Q(w2516), .D(w3519), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_3043 (.A(w3496), .nZ(w3520) );
	ym3438_AOI22 g_3044 (.A2(w3496), .B1(w2515), .A1(w336), .Z(w3521), .B2(w3520) );
	ym3438_NOR g_3045 (.Z(w3522), .B(w1111), .A(w3521) );
	ym3438_SR_BIT g_3046 (.Q(w2515), .D(w3522), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_3047 (.A(w3491), .nZ(w3523) );
	ym3438_AOI22 g_3048 (.A2(w3491), .B1(w2514), .A1(w332), .Z(w3524), .B2(w3523) );
	ym3438_NOR g_3049 (.Z(w3525), .B(w1111), .A(w3524) );
	ym3438_SR_BIT g_3050 (.Q(w2514), .D(w3525), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_3051 (.A(w3496), .nZ(w3526) );
	ym3438_AOI22 g_3052 (.A2(w3496), .B1(w2513), .A1(w332), .Z(w3527), .B2(w3526) );
	ym3438_NOR g_3053 (.Z(w3528), .B(w1111), .A(w3527) );
	ym3438_SR_BIT g_3054 (.Q(w2513), .D(w3528), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_3055 (.Q(w3542), .D(w2534), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_3056 (.Q(w3541), .D(w3542), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_3057 (.Q(w3540), .D(w3541), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_3058 (.Q(w3539), .D(w3540), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_3059 (.Q(w3538), .D(w3539), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_SR_BIT g_3060 (.Q(w2535), .D(w3538), .C1(w2425), .C2(w2426), .nC1(w2417), .nC2(w2416) );
	ym3438_NOT g_3061 (.A(w1116), .nZ(w3536) );
	ym3438_NOT g_3062 (.A(w1117), .nZ(w3537) );
	ym3438_AOI22 g_3063 (.A2(w2535), .B1(w332), .A1(w3537), .Z(w3544), .B2(w1117) );
	ym3438_NOR g_3064 (.Z(w2534), .B(w1111), .A(w3544) );
	ym3438_AND g_3065 (.Z(w584), .B(w180), .A(w3543) );
	ym3438_AND g_3066 (.Z(w553), .B(w180), .A(w2999) );
	ym3438_COMP_STR g_3067 (.A(w2998), .Z(w1146) );
	ym3438_COMP_STR g_3068 (.A(w2997), .Z(w1147) );
	ym3438_COMP_STR g_3069 (.A(w2535), .Z(w1148) );
	ym3438_NOT g_3070 (.A(w329), .nZ(w2531) );
	ym3438_NOT g_3071 (.A(w1166), .nZ(w2525) );
	ym3438_NOT g_3072 (.A(w2525), .nZ(w2526) );
	ym3438_AON22 g_3073 (.A2(w4077), .B1(w4076), .A1(w2525), .Z(w2528), .B2(w2526) );
	ym3438_AON22 g_3074 (.A2(w4079), .B1(w4078), .A1(w2525), .Z(w2527), .B2(w2526) );
	ym3438_COMP_WE g_3075 (.A(w3530), .Z(w1187) );
	ym3438_COMP_WE g_3076 (.A(w3531), .Z(w389) );
	ym3438_COMP_WE g_3077 (.A(w3532), .Z(w388) );
	ym3438_COMP_WE g_3078 (.A(w3533), .Z(w33) );
	ym3438_COMP_WE g_3079 (.A(w3534), .Z(w1168) );
	ym3438_COMP_WE g_3080 (.A(w3535), .Z(w1171) );
	ym3438_NOT g_3081 (.A(w3575), .nZ(w4076) );
	ym3438_NOT g_3082 (.A(w3592), .nZ(w4077) );
	ym3438_NOT g_3083 (.A(w3590), .nZ(w4078) );
	ym3438_NOT g_3084 (.A(w3529), .nZ(w4079) );
	ym3438_EDGE_DET g_3085 (.Q(w3000), .D(w1167), .C1(w2425), .nC1(w2417) );
	ym3438_NOT g_3086 (.A(w3000), .nZ(w2529) );
	ym3438_SLATCH g_3087 (.Q(w1470), .D(w2528), .C(w3000), .nC(w2529) );
	ym3438_SLATCH g_3088 (.Q(w1174), .D(w2527), .C(w3000), .nC(w2529) );
	ym3438_NOT g_3089 (.A(w340), .nZ(w3591) );
	ym3438_COMP_STR g_3090 (.A(w3626), .Z(w976) );
	ym3438_NOT g_3091 (.A(w3627), .nZ(w1195) );
	ym3438_NOT g_3092 (.A(w726), .nZ(w3627) );
	ym3438_NOT g_3093 (.A(w3628), .nZ(w1194) );
	ym3438_NAND g_3094 (.Z(w3628), .B(w3630), .A(w3629) );
	ym3438_NOT g_3095 (.A(w918), .nZ(w3630) );
	ym3438_SR_BIT g_3096 (.Q(w3629), .D(w1193), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_NOT g_3097 (.A(w3631), .nZ(w2586) );
	ym3438_NAND g_3098 (.Z(w3631), .B(w1193), .A(w3026) );
	ym3438_NOT g_3099 (.A(w3632), .nZ(w1193) );
	ym3438_NOT g_3100 (.A(w757), .nZ(w3632) );
	ym3438_SR_BIT g_3101 (.Q(w3026), .D(w3633), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3102 (.nQ(w3634), .D(w3635), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3103 (.A(w3634), .nZ(w3633) );
	ym3438_NOT g_3104 (.A(w3637), .nZ(w2677) );
	ym3438_DLATCH_INV g_3105 (.nQ(w3637), .D(w3009), .C(w2545), .nC(w1150) );
	ym3438_OR g_3106 (.Z(w3009), .B(w3638), .A(w3638) );
	ym3438_OR g_3107 (.Z(w3008), .B(w3639), .A(w3639) );
	ym3438_NOT g_3108 (.A(w3636), .nZ(w2536) );
	ym3438_DLATCH_INV g_3109 (.nQ(w3636), .D(w3008), .C(w2545), .nC(w1150) );
	ym3438_DLATCH_INV g_3110 (.nQ(w2877), .D(1'b1), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3111 (.A(w3640), .nZ(w2629) );
	ym3438_DLATCH_INV g_3112 (.nQ(w3640), .D(w3006), .C(w2545), .nC(w1150) );
	ym3438_OR6 g_3113 (.Z(w3006), .B(w3642), .A(w3641), .C(w3643), .D(w3644), .E(w3645), .F(w3646) );
	ym3438_NOT g_3114 (.A(w3647), .nZ(w2539) );
	ym3438_DLATCH_INV g_3115 (.nQ(w3647), .D(w3005), .C(w2545), .nC(w1150) );
	ym3438_OR g_3116 (.Z(w3005), .B(w3648), .A(w3648) );
	ym3438_NOT g_3117 (.A(w3649), .nZ(w2538) );
	ym3438_DLATCH_INV g_3118 (.nQ(w3649), .D(w3004), .C(w2545), .nC(w1150) );
	ym3438_OR g_3119 (.Z(w3004), .B(w3651), .A(w3650) );
	ym3438_NOT g_3120 (.A(w3652), .nZ(w3635) );
	ym3438_DLATCH_INV g_3121 (.nQ(w3652), .D(w3003), .C(w2545), .nC(w1150) );
	ym3438_OR7 g_3122 (.Z(w3003), .B(w3642), .A(w3020), .C(w3653), .D(w3644), .E(w3654), .F(w3646), .G(w3650) );
	ym3438_NOR g_3123 (.Z(w3655), .B(w2536), .A(w2539) );
	ym3438_DLATCH_INV g_3124 (.nQ(w3656), .D(w3655), .C(w2546), .nC(w1149) );
	ym3438_COMP_WE g_3125 (.A(w1183), .Z(w3658), .nZ(w3657) );
	ym3438_COMP_WE g_3126 (.A(w1182), .Z(w3660), .nZ(w3659) );
	ym3438_COMP_WE g_3127 (.A(w1181), .Z(w3662), .nZ(w3661) );
	ym3438_COMP_WE g_3128 (.A(w1180), .Z(w3018), .nZ(w3002) );
	ym3438_NAND4 g_3129 (.Z(w3663), .B(w3661), .A(w3002), .C(w3659), .D(w3657) );
	ym3438_NOT g_3130 (.A(w3663), .nZ(w3638) );
	ym3438_NAND4 g_3131 (.Z(w3664), .B(w3661), .A(w3002), .C(w3659), .D(w3658) );
	ym3438_NAND4 g_3132 (.Z(w3665), .B(w3661), .A(w3002), .C(w3660), .D(w3657) );
	ym3438_NOT g_3133 (.A(w3664), .nZ(w3020) );
	ym3438_NOT g_3134 (.A(w3665), .nZ(w3641) );
	ym3438_NOT g_3135 (.A(w3667), .nZ(w3668) );
	ym3438_NOT g_3136 (.A(w3669), .nZ(w3653) );
	ym3438_NAND4 g_3137 (.Z(w3666), .B(w3661), .A(w3002), .C(w3660), .D(w3658) );
	ym3438_NAND4 g_3138 (.Z(w3667), .B(w3002), .A(w3662), .C(w3659), .D(w3657) );
	ym3438_NAND4 g_3139 (.Z(w3669), .B(w3002), .A(w3662), .C(w3659), .D(w3658) );
	ym3438_NAND4 g_3140 (.Z(w3670), .B(w3002), .A(w3662), .C(w3660), .D(w3657) );
	ym3438_NAND4 g_3141 (.Z(w3671), .B(w3002), .A(w3662), .C(w3660), .D(w3658) );
	ym3438_NAND4 g_3142 (.Z(w3672), .B(w3018), .A(w3661), .C(w3659), .D(w3657) );
	ym3438_NAND4 g_3143 (.Z(w3673), .B(w3018), .A(w3661), .C(w3659), .D(w3658) );
	ym3438_NAND4 g_3144 (.Z(w3674), .B(w3018), .A(w3661), .C(w3660), .D(w3657) );
	ym3438_NAND4 g_3145 (.Z(w3675), .B(w3661), .A(w3018), .C(w3660), .D(w3658) );
	ym3438_NAND4 g_3146 (.Z(w3676), .B(w3662), .A(w3018), .C(w3659), .D(w3657) );
	ym3438_NAND4 g_3147 (.Z(w3677), .B(w3662), .A(w3018), .C(w3659), .D(w3658) );
	ym3438_NAND4 g_3148 (.Z(w3678), .B(w3662), .A(w3018), .C(w3660), .D(w3657) );
	ym3438_NAND4 g_3149 (.Z(w3679), .B(w3018), .A(w3658), .C(w3662), .D(w3660) );
	ym3438_OR4 g_3150 (.Z(w3017), .B(w3643), .A(w3653), .C(w3668), .D(w3644) );
	ym3438_OR6 g_3151 (.Z(w3016), .B(w3654), .A(w3001), .C(w3645), .D(w3646), .E(w3651), .F(w3650) );
	ym3438_OR g_3152 (.Z(w3015), .B(w3639), .A(w3648) );
	ym3438_DLATCH_INV g_3153 (.nQ(w3681), .D(w3016), .C(w2545), .nC(w1150) );
	ym3438_DLATCH_INV g_3154 (.nQ(w3682), .D(w3015), .C(w2545), .nC(w1150) );
	ym3438_NOT g_3155 (.A(w3681), .nZ(w2550) );
	ym3438_NOT g_3156 (.A(w3682), .nZ(w2549) );
	ym3438_NOT g_3157 (.A(w3680), .nZ(w2551) );
	ym3438_NOT g_3158 (.A(w3679), .nZ(w3639) );
	ym3438_NOT g_3159 (.A(w3678), .nZ(w3648) );
	ym3438_NOT g_3160 (.A(w3677), .nZ(w3650) );
	ym3438_NOT g_3161 (.A(w3676), .nZ(w3651) );
	ym3438_NOT g_3162 (.A(w3675), .nZ(w3646) );
	ym3438_NOT g_3163 (.A(w3674), .nZ(w3645) );
	ym3438_NOT g_3164 (.A(w3670), .nZ(w3643) );
	ym3438_NOT g_3165 (.A(w3671), .nZ(w3644) );
	ym3438_NOT g_3166 (.A(w3672), .nZ(w3001) );
	ym3438_NOT g_3167 (.A(w3673), .nZ(w3654) );
	ym3438_DLATCH_INV g_3168 (.nQ(w3680), .D(w3017), .C(w2545), .nC(w1150) );
	ym3438_NOT g_3169 (.A(w3666), .nZ(w3642) );
	ym3438_AON21SR g_3170 (.Q(w3626), .C2(w2546), .nC2(w1149), .C1(w2545), .nC1(w1150), .B(w3066), .A1(w3700), .A2(w1195) );
	ym3438_SDELAY24 g_3171 (.A(w3025), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .Q(w3700), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .C36(w2546), .nC36(w1149), .C35(w2545), .nC35(w1150), .C34(w2546), .nC34(w1149), .C33(w2545), .nC33(w1150), .C32(w2546), .nC32(w1149), .C31(w2545), .nC31(w1150), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150) );
	ym3438_AND g_3172 (.Z(w3064), .B(w1194), .A(w3700) );
	ym3438_FA g_3173 (.CO(w3703), .S(w3025), .CI(1'b0), .A(w3699), .B(w3064) );
	ym3438_NOT g_3174 (.A(w3698), .nZ(w3699) );
	ym3438_DLATCH_INV g_3175 (.nQ(w3698), .D(w3062), .C(w2546), .nC(w1149) );
	ym3438_FA g_3176 (.CO(w3063), .S(w3062), .CI(1'b0), .A(w3697), .B(w3061) );
	ym3438_DLATCH_INV g_3177 (.nQ(w3697), .D(w3024), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3178 (.Z(w3024), .B(w1193), .A(w3023) );
	ym3438_DLATCH_INV g_3179 (.nQ(w3061), .D(w3057), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3180 (.Z(w3057), .B(w3695), .A(w2586) );
	ym3438_SR_BIT g_3181 (.Q(w3695), .D(w3694), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3182 (.nQ(w3693), .D(w3056), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3183 (.A(w3693), .nZ(w3694) );
	ym3438_FA_SEQ g_3184 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .CO(w3055), .Q(w3023), .CI(w3656), .A(1'b0), .B(w3022) );
	ym3438_DLATCH_INV g_3185 (.nQ(w3022), .D(w3021), .C(w2546), .nC(w1149) );
	ym3438_AON21SR g_3186 (.Q(w3066), .C2(w2546), .nC2(w1149), .C1(w2545), .nC1(w1150), .B(w3701), .A1(w3065), .A2(w1195) );
	ym3438_SDELAY24 g_3187 (.A(w3084), .Q(w3065), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .nC36(w1149), .nC35(w1150), .nC34(w1149), .nC33(w1150), .nC32(w1149), .nC31(w1150), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .C36(w2546), .C35(w2545), .C34(w2546), .C33(w2545), .C32(w2546), .C31(w2545) );
	ym3438_AND g_3188 (.Z(w3702), .B(w3065), .A(w1194) );
	ym3438_FA g_3189 (.CO(w3085), .S(w3084), .CI(w3703), .A(w3704), .B(w3702) );
	ym3438_NOT g_3190 (.A(w3705), .nZ(w3704) );
	ym3438_DLATCH_INV g_3191 (.nQ(w3705), .D(w3060), .C(w2546), .nC(w1149) );
	ym3438_FA g_3192 (.CO(w3083), .S(w3060), .CI(w3063), .A(w3706), .B(w3059) );
	ym3438_DLATCH_INV g_3193 (.nQ(w3706), .D(w3081), .C(w2545), .nC(w1150) );
	ym3438_DLATCH_INV g_3194 (.nQ(w3059), .D(w3058), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3195 (.Z(w3081), .B(w3079), .A(w1193) );
	ym3438_NAND g_3196 (.Z(w3058), .B(w3696), .A(w2586) );
	ym3438_SR_BIT g_3197 (.Q(w3696), .D(w3707), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3198 (.nQ(w3708), .D(w3052), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3199 (.A(w3708), .nZ(w3707) );
	ym3438_FA_SEQ g_3200 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .CO(w3709), .Q(w3079), .CI(w3055), .A(1'b0), .B(w3076) );
	ym3438_AON21SR g_3201 (.Q(w3701), .C2(w2546), .nC2(w1149), .C1(w2545), .nC1(w1150), .B(w3189), .A1(w3722), .A2(w1195) );
	ym3438_SDELAY24 g_3202 (.A(w3086), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .Q(w3722), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .C36(w2546), .nC36(w1149), .C35(w2545), .nC35(w1150), .C34(w2546), .nC34(w1149), .C33(w2545), .nC33(w1150), .C32(w2546), .nC32(w1149), .C31(w2545), .nC31(w1150), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150) );
	ym3438_AND g_3203 (.Z(w3188), .B(w1194), .A(w3722) );
	ym3438_FA g_3204 (.CO(w3186), .S(w3086), .CI(w3085), .A(w3744), .B(w3188) );
	ym3438_NOT g_3205 (.A(w3745), .nZ(w3744) );
	ym3438_DLATCH_INV g_3206 (.nQ(w3745), .D(w3185), .C(w2546), .nC(w1149) );
	ym3438_FA g_3207 (.CO(w3183), .S(w3185), .CI(w3083), .A(w3783), .B(w3181) );
	ym3438_DLATCH_INV g_3208 (.nQ(w3783), .D(w3082), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3209 (.Z(w3082), .B(w1193), .A(w3080) );
	ym3438_DLATCH_INV g_3210 (.nQ(w3181), .D(w3179), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3211 (.Z(w3179), .B(w3785), .A(w2586) );
	ym3438_SR_BIT g_3212 (.Q(w3785), .D(w3782), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3213 (.nQ(w3837), .D(w3051), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3214 (.A(w3837), .nZ(w3782) );
	ym3438_FA_SEQ g_3215 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .CO(w3178), .Q(w3080), .CI(w3709), .A(w3176), .B(w3077) );
	ym3438_AON21SR g_3216 (.Q(w3189), .C2(w2546), .nC2(w1149), .C1(w2545), .nC1(w1150), .B(w3741), .A1(w3723), .A2(w1195) );
	ym3438_SDELAY24 g_3217 (.A(w3148), .Q(w3723), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .nC36(w1149), .nC35(w1150), .nC34(w1149), .nC33(w1150), .nC32(w1149), .nC31(w1150), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .C36(w2546), .C35(w2545), .C34(w2546), .C33(w2545), .C32(w2546), .C31(w2545) );
	ym3438_AND g_3218 (.Z(w3187), .B(w3723), .A(w1194) );
	ym3438_FA g_3219 (.CO(w3146), .S(w3148), .CI(w3186), .A(w3746), .B(w3187) );
	ym3438_NOT g_3220 (.A(w3747), .nZ(w3746) );
	ym3438_DLATCH_INV g_3221 (.nQ(w3747), .D(w3184), .C(w2546), .nC(w1149) );
	ym3438_FA g_3222 (.CO(w3145), .S(w3184), .CI(w3183), .A(w3784), .B(w3182) );
	ym3438_DLATCH_INV g_3223 (.nQ(w3784), .D(w3144), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3224 (.Z(w3144), .B(w3142), .A(w1193) );
	ym3438_DLATCH_INV g_3225 (.nQ(w3182), .D(w3180), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3226 (.Z(w3180), .B(w3786), .A(w2586) );
	ym3438_SR_BIT g_3227 (.Q(w3786), .D(w3820), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3228 (.nQ(w3838), .D(w3106), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3229 (.A(w3838), .nZ(w3820) );
	ym3438_FA_SEQ g_3230 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .CO(w3852), .Q(w3142), .CI(w3178), .A(w3177), .B(w3139) );
	ym3438_AON21SR g_3231 (.Q(w3741), .C2(w2546), .nC2(w1149), .C1(w2545), .nC1(w1150), .B(w3122), .A1(w3724), .A2(w1195) );
	ym3438_SDELAY24 g_3232 (.A(w3147), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .Q(w3724), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .C36(w2546), .nC36(w1149), .C35(w2545), .nC35(w1150), .C34(w2546), .nC34(w1149), .C33(w2545), .nC33(w1150), .C32(w2546), .nC32(w1149), .C31(w2545), .nC31(w1150), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150) );
	ym3438_AND g_3233 (.Z(w3121), .B(w1194), .A(w3724) );
	ym3438_FA g_3234 (.CO(w3119), .S(w3147), .CI(w3146), .A(w3748), .B(w3121) );
	ym3438_NOT g_3235 (.A(w3749), .nZ(w3748) );
	ym3438_DLATCH_INV g_3236 (.nQ(w3749), .D(w3118), .C(w2546), .nC(w1149) );
	ym3438_FA g_3237 (.CO(w3116), .S(w3118), .CI(w3145), .A(w3787), .B(w3115) );
	ym3438_NAND g_3238 (.Z(w3821), .B(w1193), .A(w3143) );
	ym3438_DLATCH_INV g_3239 (.nQ(w3787), .D(w3821), .C(w2545), .nC(w1150) );
	ym3438_DLATCH_INV g_3240 (.nQ(w3115), .D(w3789), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3241 (.Z(w3789), .B(w3790), .A(w2586) );
	ym3438_SR_BIT g_3242 (.Q(w3790), .D(w3822), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3243 (.nQ(w3839), .D(w3112), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3244 (.A(w3839), .nZ(w3822) );
	ym3438_FA_SEQ g_3245 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .CO(w3111), .Q(w3143), .CI(w3852), .A(w3108), .B(w3141) );
	ym3438_SDELAY24 g_3246 (.A(w3105), .Q(w3740), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .nC36(w1149), .nC35(w1150), .nC34(w1149), .nC33(w1150), .nC32(w1149), .nC31(w1150), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .C36(w2546), .C35(w2545), .C34(w2546), .C33(w2545), .C32(w2546), .C31(w2545) );
	ym3438_AON21SR g_3247 (.Q(w3122), .C2(w2546), .nC2(w1149), .C1(w2545), .nC1(w1150), .B(w3742), .A1(w3740), .A2(w1195) );
	ym3438_AND g_3248 (.Z(w3120), .B(w3740), .A(w1194) );
	ym3438_FA g_3249 (.CO(w3103), .S(w3105), .CI(w3119), .A(w3750), .B(w3120) );
	ym3438_NOT g_3250 (.A(w3751), .nZ(w3750) );
	ym3438_DLATCH_INV g_3251 (.nQ(w3751), .D(w3117), .C(w2546), .nC(w1149) );
	ym3438_FA g_3252 (.CO(w3102), .S(w3117), .CI(w3116), .A(w3788), .B(w3114) );
	ym3438_DLATCH_INV g_3253 (.nQ(w3788), .D(w3101), .C(w2545), .nC(w1150) );
	ym3438_DLATCH_INV g_3254 (.nQ(w3114), .D(w3113), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3255 (.Z(w3101), .B(w3099), .A(w1193) );
	ym3438_NAND g_3256 (.Z(w3113), .B(w3791), .A(w2586) );
	ym3438_SR_BIT g_3257 (.Q(w3791), .D(w3823), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3258 (.nQ(w3840), .D(w2958), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3259 (.A(w3840), .nZ(w3823) );
	ym3438_FA_SEQ g_3260 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .CO(w3853), .Q(w3099), .CI(w3111), .A(w3109), .B(w3095) );
	ym3438_AON21SR g_3261 (.Q(w3742), .C2(w2546), .nC2(w1149), .C1(w2545), .nC1(w1150), .B(w2975), .A1(w3725), .A2(w1195) );
	ym3438_SDELAY24 g_3262 (.A(w3104), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .Q(w3725), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .C36(w2546), .nC36(w1149), .C35(w2545), .nC35(w1150), .C34(w2546), .nC34(w1149), .C33(w2545), .nC33(w1150), .C32(w2546), .nC32(w1149), .C31(w2545), .nC31(w1150), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150) );
	ym3438_AND g_3263 (.Z(w2972), .B(w1194), .A(w3725) );
	ym3438_FA g_3264 (.CO(w2973), .S(w3104), .CI(w3103), .A(w3752), .B(w2972) );
	ym3438_NOT g_3265 (.A(w3753), .nZ(w3752) );
	ym3438_DLATCH_INV g_3266 (.nQ(w3753), .D(w2970), .C(w2546), .nC(w1149) );
	ym3438_FA g_3267 (.CO(w2971), .S(w2970), .CI(w3102), .A(w3792), .B(w2967) );
	ym3438_DLATCH_INV g_3268 (.nQ(w3792), .D(w3100), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3269 (.Z(w3100), .B(w1193), .A(w3098) );
	ym3438_DLATCH_INV g_3270 (.nQ(w2967), .D(w2965), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3271 (.Z(w2965), .B(w3794), .A(w2586) );
	ym3438_SR_BIT g_3272 (.Q(w3794), .D(w3824), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_NOT g_3273 (.A(w3841), .nZ(w3824) );
	ym3438_DLATCH_INV g_3274 (.nQ(w3841), .D(w2964), .C(w2546), .nC(w1149) );
	ym3438_FA_SEQ g_3275 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .CO(w2963), .Q(w3098), .CI(w3853), .A(w2962), .B(w3096) );
	ym3438_AON21SR g_3276 (.Q(w2975), .C2(w2546), .nC2(w1149), .C1(w2545), .nC1(w1150), .B(w2944), .A1(w3739), .A2(w1195) );
	ym3438_SDELAY24 g_3277 (.A(w2941), .Q(w3739), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .nC36(w1149), .nC35(w1150), .nC34(w1149), .nC33(w1150), .nC32(w1149), .nC31(w1150), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .C36(w2546), .C35(w2545), .C34(w2546), .C33(w2545), .C32(w2546), .C31(w2545) );
	ym3438_AND g_3278 (.Z(w2974), .B(w3739), .A(w1194) );
	ym3438_FA g_3279 (.CO(w2942), .S(w2941), .CI(w2973), .A(w3754), .B(w2974) );
	ym3438_NOT g_3280 (.A(w3755), .nZ(w3754) );
	ym3438_DLATCH_INV g_3281 (.nQ(w3755), .D(w2969), .C(w2546), .nC(w1149) );
	ym3438_FA g_3282 (.CO(w2940), .S(w2969), .CI(w2971), .A(w3793), .B(w2968) );
	ym3438_DLATCH_INV g_3283 (.nQ(w3793), .D(w2938), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3284 (.Z(w2938), .B(w2937), .A(w1193) );
	ym3438_DLATCH_INV g_3285 (.nQ(w2968), .D(w2966), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3286 (.Z(w2966), .B(w3795), .A(w2586) );
	ym3438_SR_BIT g_3287 (.Q(w3795), .D(w3825), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3288 (.nQ(w3842), .D(w2899), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3289 (.A(w3842), .nZ(w3825) );
	ym3438_FA_SEQ g_3290 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .CO(w3854), .Q(w2937), .CI(w2963), .A(w2961), .B(w2933) );
	ym3438_AON21SR g_3291 (.Q(w2944), .C2(w2546), .nC2(w1149), .C1(w2545), .nC1(w1150), .B(w2916), .A1(w3726), .A2(w1195) );
	ym3438_SDELAY24 g_3292 (.A(w2943), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .Q(w3726), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .C36(w2546), .nC36(w1149), .C35(w2545), .nC35(w1150), .C34(w2546), .nC34(w1149), .C33(w2545), .nC33(w1150), .C32(w2546), .nC32(w1149), .C31(w2545), .nC31(w1150), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150) );
	ym3438_AND g_3293 (.Z(w2915), .B(w1194), .A(w3726) );
	ym3438_FA g_3294 (.CO(w2913), .S(w2943), .CI(w2942), .A(w3756), .B(w2915) );
	ym3438_NOT g_3295 (.A(w3757), .nZ(w3756) );
	ym3438_DLATCH_INV g_3296 (.nQ(w3757), .D(w2909), .C(w2546), .nC(w1149) );
	ym3438_FA g_3297 (.CO(w2912), .S(w2909), .CI(w2940), .A(w3796), .B(w2908) );
	ym3438_DLATCH_INV g_3298 (.nQ(w3796), .D(w2939), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3299 (.Z(w2939), .B(w1193), .A(w2936) );
	ym3438_DLATCH_INV g_3300 (.nQ(w2908), .D(w2906), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3301 (.Z(w2906), .B(w3798), .A(w2586) );
	ym3438_SR_BIT g_3302 (.Q(w3798), .D(w3826), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3303 (.nQ(w3843), .D(w2905), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3304 (.A(w3843), .nZ(w3826) );
	ym3438_FA_SEQ g_3305 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .CO(w2904), .Q(w2936), .CI(w3854), .A(w2901), .B(w2935) );
	ym3438_AON21SR g_3306 (.Q(w2916), .C2(w2546), .nC2(w1149), .C1(w2545), .nC1(w1150), .B(w2877), .A1(w3738), .A2(w1195) );
	ym3438_SDELAY24 g_3307 (.A(w2876), .Q(w3738), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .nC36(w1149), .nC35(w1150), .nC34(w1149), .nC33(w1150), .nC32(w1149), .nC31(w1150), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .C36(w2546), .C35(w2545), .C34(w2546), .C33(w2545), .C32(w2546), .C31(w2545) );
	ym3438_AND g_3308 (.Z(w2914), .B(w3738), .A(w1194) );
	ym3438_FA g_3309 (.CO(w2874), .S(w2876), .CI(w2913), .A(w3758), .B(w2914) );
	ym3438_NOT g_3310 (.A(w3759), .nZ(w3758) );
	ym3438_DLATCH_INV g_3311 (.nQ(w3759), .D(w2911), .C(w2546), .nC(w1149) );
	ym3438_FA g_3312 (.CO(w2873), .S(w2911), .CI(w2912), .A(w3797), .B(w2910) );
	ym3438_DLATCH_INV g_3313 (.nQ(w3797), .D(w2872), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3314 (.Z(w2872), .B(w2869), .A(w1193) );
	ym3438_DLATCH_INV g_3315 (.nQ(w2910), .D(w2907), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3316 (.Z(w2907), .B(w3799), .A(w2586) );
	ym3438_SR_BIT g_3317 (.Q(w3799), .D(w3827), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3318 (.nQ(w3844), .D(w2834), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3319 (.A(w3844), .nZ(w3827) );
	ym3438_FA_SEQ g_3320 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .CO(w3855), .Q(w2869), .CI(w2904), .A(w2903), .B(w2866) );
	ym3438_SDELAY24 g_3321 (.A(w2875), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .Q(w3727), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .C36(w2546), .nC36(w1149), .C35(w2545), .nC35(w1150), .C34(w2546), .nC34(w1149), .C33(w2545), .nC33(w1150), .C32(w2546), .nC32(w1149), .C31(w2545), .nC31(w1150), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150), .Q40(w2878) );
	ym3438_AND g_3322 (.Z(w2848), .B(w1194), .A(w3727) );
	ym3438_FA g_3323 (.CO(w2849), .S(w2875), .CI(w2874), .A(w3760), .B(w2848) );
	ym3438_NOT g_3324 (.A(w3761), .nZ(w3760) );
	ym3438_DLATCH_INV g_3325 (.nQ(w3761), .D(w2844), .C(w2546), .nC(w1149) );
	ym3438_FA g_3326 (.CO(w2846), .S(w2844), .CI(w2873), .A(w3800), .B(w2843) );
	ym3438_DLATCH_INV g_3327 (.nQ(w3800), .D(w2871), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3328 (.Z(w2871), .B(w1193), .A(w2870) );
	ym3438_DLATCH_INV g_3329 (.nQ(w2843), .D(w2842), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3330 (.Z(w2842), .B(w3802), .A(w2586) );
	ym3438_SR_BIT g_3331 (.Q(w3802), .D(w3828), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3332 (.nQ(w3845), .D(w2840), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3333 (.A(w3845), .nZ(w3828) );
	ym3438_FA_SEQ g_3334 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .CO(w2839), .Q(w2870), .CI(w3855), .A(w2836), .B(w2868) );
	ym3438_SDELAY24 g_3335 (.A(w2809), .Q(w3736), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .nC36(w1149), .nC35(w1150), .nC34(w1149), .nC33(w1150), .nC32(w1149), .nC31(w1150), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .C36(w2546), .C35(w2545), .C34(w2546), .C33(w2545), .C32(w2546), .C31(w2545), .Q40(w2810) );
	ym3438_AND g_3336 (.Z(w3737), .B(w1194), .A(w3736) );
	ym3438_FA g_3337 (.S(w2809), .CI(w2849), .A(w3762), .B(w3737), .CO(w2807) );
	ym3438_NOT g_3338 (.A(w3763), .nZ(w3762) );
	ym3438_DLATCH_INV g_3339 (.nQ(w3763), .D(w2847), .C(w2546), .nC(w1149) );
	ym3438_FA g_3340 (.CO(w2806), .S(w2847), .CI(w2846), .A(w3801), .B(w2845) );
	ym3438_DLATCH_INV g_3341 (.nQ(w3801), .D(w2803), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3342 (.Z(w2803), .B(w2802), .A(w1193) );
	ym3438_DLATCH_INV g_3343 (.nQ(w2845), .D(w2841), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3344 (.Z(w2841), .B(w3803), .A(w2586) );
	ym3438_SR_BIT g_3345 (.Q(w3803), .D(w3829), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3346 (.nQ(w3846), .D(w2764), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3347 (.A(w3846), .nZ(w3829) );
	ym3438_FA_SEQ g_3348 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .CO(w3856), .Q(w2802), .CI(w2839), .A(w2838), .B(w2799) );
	ym3438_SDELAY24 g_3349 (.A(w2808), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .Q(w3728), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .C36(w2546), .nC36(w1149), .C35(w2545), .nC35(w1150), .C34(w2546), .nC34(w1149), .C33(w2545), .nC33(w1150), .C32(w2546), .nC32(w1149), .C31(w2545), .nC31(w1150), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150), .Q40(w2811) );
	ym3438_AND g_3350 (.Z(w2779), .B(w1194), .A(w3728) );
	ym3438_FA g_3351 (.CO(w2777), .S(w2808), .CI(w2807), .A(w3764), .B(w2779) );
	ym3438_NOT g_3352 (.A(w3765), .nZ(w3764) );
	ym3438_DLATCH_INV g_3353 (.nQ(w3765), .D(w2776), .C(w2546), .nC(w1149) );
	ym3438_FA g_3354 (.CO(w2774), .S(w2776), .CI(w2806), .A(w3804), .B(w2775) );
	ym3438_DLATCH_INV g_3355 (.nQ(w3804), .D(w2804), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3356 (.Z(w2804), .B(w1193), .A(w2805) );
	ym3438_DLATCH_INV g_3357 (.nQ(w2775), .D(w2771), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3358 (.Z(w2771), .B(w3806), .A(w2586) );
	ym3438_SR_BIT g_3359 (.Q(w3806), .D(w3830), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3360 (.nQ(w3847), .D(w2725), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3361 (.A(w3847), .nZ(w3830) );
	ym3438_FA_SEQ g_3362 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .CO(w2769), .Q(w2805), .CI(w3856), .A(w2766), .B(w2801) );
	ym3438_SDELAY24 g_3363 (.A(w2738), .Q(w3735), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .nC36(w1149), .nC35(w1150), .nC34(w1149), .nC33(w1150), .nC32(w1149), .nC31(w1150), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .C36(w2546), .C35(w2545), .C34(w2546), .C33(w2545), .C32(w2546), .C31(w2545), .Q40(w2739) );
	ym3438_AND g_3364 (.Z(w2778), .B(w1194), .A(w3735) );
	ym3438_FA g_3365 (.S(w2738), .CI(w2777), .A(w3766), .B(w2778), .CO(w2736) );
	ym3438_NOT g_3366 (.A(w3767), .nZ(w3766) );
	ym3438_DLATCH_INV g_3367 (.nQ(w3767), .D(w2773), .C(w2546), .nC(w1149) );
	ym3438_FA g_3368 (.CO(w2735), .S(w2773), .CI(w2774), .A(w3805), .B(w2772) );
	ym3438_DLATCH_INV g_3369 (.nQ(w3805), .D(w2733), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3370 (.Z(w2733), .B(w2732), .A(w1193) );
	ym3438_DLATCH_INV g_3371 (.nQ(w2772), .D(w2770), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3372 (.Z(w2770), .B(w3807), .A(w2586) );
	ym3438_SR_BIT g_3373 (.Q(w3807), .D(w4363), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3374 (.nQ(w3848), .D(w2694), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3375 (.A(w3848), .nZ(w4363) );
	ym3438_FA_SEQ g_3376 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .CO(w3857), .Q(w2732), .CI(w2769), .A(w2768), .B(w2729) );
	ym3438_SDELAY24 g_3377 (.A(w2737), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .Q(w3729), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .C36(w2546), .nC36(w1149), .C35(w2545), .nC35(w1150), .C34(w2546), .nC34(w1149), .C33(w2545), .nC33(w1150), .C32(w2546), .nC32(w1149), .C31(w2545), .nC31(w1150), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150), .Q40(w2740) );
	ym3438_AND g_3378 (.Z(w2707), .B(w1194), .A(w3729) );
	ym3438_FA g_3379 (.CO(w2708), .S(w2737), .CI(w2736), .A(w3768), .B(w2707) );
	ym3438_NOT g_3380 (.A(w3769), .nZ(w3768) );
	ym3438_DLATCH_INV g_3381 (.nQ(w3769), .D(w2704), .C(w2546), .nC(w1149) );
	ym3438_FA g_3382 (.CO(w2706), .S(w2704), .CI(w2735), .A(w3808), .B(w2703) );
	ym3438_DLATCH_INV g_3383 (.nQ(w3808), .D(w2734), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3384 (.Z(w2734), .B(w1193), .A(w2731) );
	ym3438_DLATCH_INV g_3385 (.nQ(w2703), .D(w2700), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3386 (.Z(w2700), .B(w3810), .A(w2586) );
	ym3438_SR_BIT g_3387 (.Q(w3810), .D(w3831), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3388 (.nQ(w3849), .D(w2662), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3389 (.A(w3849), .nZ(w3831) );
	ym3438_FA_SEQ g_3390 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .CO(w2699), .Q(w2731), .CI(w3857), .A(w2696), .B(w2730) );
	ym3438_COMP_STR g_3391 (.A(w2878), .Z(w1192) );
	ym3438_COMP_STR g_3392 (.A(w2810), .Z(w1191) );
	ym3438_COMP_STR g_3393 (.A(w2811), .Z(w1190) );
	ym3438_COMP_STR g_3394 (.A(w2739), .Z(w1189) );
	ym3438_COMP_STR g_3395 (.A(w2740), .Z(w1188) );
	ym3438_SDELAY24 g_3396 (.A(w2673), .Q(w3734), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .nC36(w1149), .nC35(w1150), .nC34(w1149), .nC33(w1150), .nC32(w1149), .nC31(w1150), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .C36(w2546), .C35(w2545), .C34(w2546), .C33(w2545), .C32(w2546), .C31(w2545), .Q40(w2676) );
	ym3438_AND g_3397 (.Z(w2709), .B(w1194), .A(w3734) );
	ym3438_FA g_3398 (.S(w2673), .CI(w2708), .A(w3770), .B(w2709), .CO(w2674) );
	ym3438_NOT g_3399 (.A(w3771), .nZ(w3770) );
	ym3438_DLATCH_INV g_3400 (.nQ(w3771), .D(w2705), .C(w2546), .nC(w1149) );
	ym3438_FA g_3401 (.CO(w2672), .S(w2705), .CI(w2706), .A(w3809), .B(w2702) );
	ym3438_DLATCH_INV g_3402 (.nQ(w3809), .D(w2671), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3403 (.Z(w2671), .B(w2668), .A(w1193) );
	ym3438_DLATCH_INV g_3404 (.nQ(w2702), .D(w2701), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3405 (.Z(w2701), .B(w3811), .A(w2586) );
	ym3438_SR_BIT g_3406 (.Q(w3811), .D(w3832), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3407 (.nQ(w3850), .D(w2643), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3408 (.A(w3850), .nZ(w3832) );
	ym3438_FA_SEQ g_3409 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .CO(w3858), .Q(w2668), .CI(w2699), .A(w2698), .B(w2666) );
	ym3438_COMP_STR g_3410 (.A(w2676), .Z(w1323) );
	ym3438_SDELAY24 g_3411 (.A(w2675), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .Q(w3730), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .C36(w2546), .nC36(w1149), .C35(w2545), .nC35(w1150), .C34(w2546), .nC34(w1149), .C33(w2545), .nC33(w1150), .C32(w2546), .nC32(w1149), .C31(w2545), .nC31(w1150), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150), .Q40(w3743) );
	ym3438_AND g_3412 (.Z(w2657), .B(w1194), .A(w3730) );
	ym3438_FA g_3413 (.CO(w2655), .S(w2675), .CI(w2674), .A(w3772), .B(w2657) );
	ym3438_NOT g_3414 (.A(w3773), .nZ(w3772) );
	ym3438_DLATCH_INV g_3415 (.nQ(w3773), .D(w2652), .C(w2546), .nC(w1149) );
	ym3438_FA g_3416 (.CO(w2654), .S(w2652), .CI(w2672), .A(w3812), .B(w2651) );
	ym3438_DLATCH_INV g_3417 (.nQ(w3812), .D(w2670), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3418 (.Z(w2670), .B(w1193), .A(w2669) );
	ym3438_DLATCH_INV g_3419 (.nQ(w2651), .D(w2650), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3420 (.Z(w2650), .B(w3814), .A(w2586) );
	ym3438_SR_BIT g_3421 (.Q(w3814), .D(w3833), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3422 (.nQ(w3851), .D(w2581), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3423 (.A(w3851), .nZ(w3833) );
	ym3438_FA_SEQ g_3424 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .CO(w2648), .Q(w2669), .CI(w3858), .A(w2645), .B(w2667) );
	ym3438_COMP_STR g_3425 (.A(w3743), .Z(w1270) );
	ym3438_SDELAY24 g_3426 (.A(w2627), .Q(w3733), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .nC36(w1149), .nC35(w1150), .nC34(w1149), .nC33(w1150), .nC32(w1149), .nC31(w1150), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .C36(w2546), .C35(w2545), .C34(w2546), .C33(w2545), .C32(w2546), .C31(w2545), .Q40(w2628) );
	ym3438_AND g_3427 (.Z(w2656), .B(w1194), .A(w3733) );
	ym3438_FA g_3428 (.S(w2627), .CI(w2655), .A(w3774), .B(w2656), .CO(w2598) );
	ym3438_NOT g_3429 (.A(w3775), .nZ(w3774) );
	ym3438_DLATCH_INV g_3430 (.nQ(w3775), .D(w2653), .C(w2546), .nC(w1149) );
	ym3438_FA g_3431 (.CO(w3780), .S(w2653), .CI(w2654), .A(w3813), .B(w3781) );
	ym3438_DLATCH_INV g_3432 (.nQ(w3813), .D(w2626), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3433 (.Z(w2626), .B(w2625), .A(w1193) );
	ym3438_DLATCH_INV g_3434 (.nQ(w3781), .D(w2649), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3435 (.Z(w2649), .B(w3815), .A(w2586) );
	ym3438_SR_BIT g_3436 (.Q(w3815), .D(1'b0), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_FA_SEQ g_3437 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .CO(w3859), .Q(w2625), .CI(w2648), .A(w2647), .B(w2621) );
	ym3438_COMP_STR g_3438 (.A(w2628), .Z(w1276) );
	ym3438_SDELAY24 g_3439 (.A(w2597), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .Q(w3731), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .C36(w2546), .nC36(w1149), .C35(w2545), .nC35(w1150), .C34(w2546), .nC34(w1149), .C33(w2545), .nC33(w1150), .C32(w2546), .nC32(w1149), .C31(w2545), .nC31(w1150), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150), .Q40(w2630) );
	ym3438_AND g_3440 (.Z(w2596), .B(w1194), .A(w3731) );
	ym3438_FA g_3441 (.CO(w2595), .S(w2597), .CI(w2598), .A(w3776), .B(w2596) );
	ym3438_NOT g_3442 (.A(w3777), .nZ(w3776) );
	ym3438_DLATCH_INV g_3443 (.nQ(w3777), .D(w2593), .C(w2546), .nC(w1149) );
	ym3438_FA g_3444 (.CO(w2591), .S(w2593), .CI(w3780), .A(w3816), .B(w2592) );
	ym3438_DLATCH_INV g_3445 (.nQ(w3816), .D(w2599), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3446 (.Z(w2599), .B(w1193), .A(w2600) );
	ym3438_DLATCH_INV g_3447 (.nQ(w2592), .D(w2588), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3448 (.Z(w2588), .B(w3818), .A(w2586) );
	ym3438_SR_BIT g_3449 (.Q(w3818), .D(1'b0), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_FA_SEQ g_3450 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .CO(w2585), .Q(w2600), .CI(w3859), .A(w2583), .B(w2624) );
	ym3438_COMP_STR g_3451 (.A(w2630), .Z(w1324) );
	ym3438_SDELAY24 g_3452 (.A(w3197), .Q(w3732), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .C3(w2545), .C4(w2546), .C5(w2545), .C6(w2546), .C7(w2545), .C8(w2546), .C9(w2545), .C10(w2546), .C11(w2545), .C12(w2546), .C13(w2545), .C14(w2546), .C15(w2545), .C16(w2546), .C17(w2545), .C18(w2546), .C19(w2545), .C20(w2546), .C21(w2545), .C22(w2546), .C23(w2545), .C24(w2546), .nC3(w1150), .nC4(w1149), .nC5(w1150), .nC6(w1149), .nC7(w1150), .nC8(w1149), .nC9(w1150), .nC10(w1149), .nC11(w1150), .nC12(w1149), .nC13(w1150), .nC14(w1149), .nC15(w1150), .nC16(w1149), .nC17(w1150), .nC18(w1149), .nC19(w1150), .nC20(w1149), .nC21(w1150), .nC22(w1149), .nC23(w1150), .nC24(w1149), .C42(w2546), .nC42(w1149), .C41(w2545), .nC41(w1150), .C40(w2546), .nC40(w1149), .C39(w2545), .nC39(w1150), .C38(w2546), .nC38(w1149), .C37(w2545), .nC37(w1150), .C44(w2546), .nC44(w1149), .C43(w2545), .nC43(w1150), .C46(w2546), .nC46(w1149), .C45(w2545), .nC45(w1150), .C48(w2546), .nC48(w1149), .C47(w2545), .nC47(w1150), .nC25(w1150), .nC26(w1149), .nC27(w1150), .nC28(w1149), .nC29(w1150), .nC30(w1149), .nC36(w1149), .nC35(w1150), .nC34(w1149), .nC33(w1150), .nC32(w1149), .nC31(w1150), .C25(w2545), .C26(w2546), .C27(w2545), .C28(w2546), .C29(w2545), .C30(w2546), .C36(w2546), .C35(w2545), .C34(w2546), .C33(w2545), .C32(w2546), .C31(w2545), .Q40(w2537) );
	ym3438_AND g_3453 (.Z(w2594), .B(w1194), .A(w3732) );
	ym3438_FA g_3454 (.S(w3197), .CI(w2595), .A(w3778), .B(w2594) );
	ym3438_NOT g_3455 (.A(w3779), .nZ(w3778) );
	ym3438_DLATCH_INV g_3456 (.nQ(w3779), .D(w2590), .C(w2546), .nC(w1149) );
	ym3438_FA g_3457 (.S(w2590), .CI(w2591), .A(w3817), .B(w2589) );
	ym3438_DLATCH_INV g_3458 (.nQ(w3817), .D(w3196), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3459 (.Z(w3196), .B(w3195), .A(w1193) );
	ym3438_DLATCH_INV g_3460 (.nQ(w2589), .D(w2587), .C(w2545), .nC(w1150) );
	ym3438_NAND g_3461 (.Z(w2587), .B(w3819), .A(w2586) );
	ym3438_SR_BIT g_3462 (.Q(w3819), .D(1'b0), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_FA_SEQ g_3463 (.C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .Q(w3195), .CI(w2585), .A(w2584), .B(w3194) );
	ym3438_COMP_STR g_3464 (.A(w2537), .Z(w1277) );
	ym3438_AOI222222 g_3465 (.A2(1'b0), .B1(w3052), .A1(1'b0), .Z(w3021), .B2(w2677), .C1(w3053), .C2(w2536), .D1(1'b0), .D2(w2629), .E1(1'b1), .E2(w2539), .F1(1'b0), .F2(w2538) );
	ym3438_SLATCH g_3466 (.Q(w3691), .D(w3047), .C(w3685), .nC(w3684) );
	ym3438_XOR g_3467 (.Z(w3690), .B(w3687), .A(w3691) );
	ym3438_XOR g_3468 (.Z(w3049), .B(w3687), .A(w3689) );
	ym3438_SLATCH g_3469 (.Q(w3689), .D(w3050), .C(w3685), .nC(w3684) );
	ym3438_SLATCH g_3470 (.Q(w3038), .D(w3046), .C(w3685), .nC(w3684) );
	ym3438_XOR g_3471 (.Z(w3048), .B(w3687), .A(w3038) );
	ym3438_SLATCH g_3472 (.Q(w3039), .D(w3044), .C(w3685), .nC(w3684) );
	ym3438_XOR g_3473 (.Z(w3045), .B(w3687), .A(w3039) );
	ym3438_SLATCH g_3474 (.Q(w3036), .D(w3042), .C(w3685), .nC(w3684) );
	ym3438_XOR g_3475 (.Z(w3043), .B(w3687), .A(w3036) );
	ym3438_SLATCH g_3476 (.Q(w3037), .D(w3041), .C(w3685), .nC(w3684) );
	ym3438_XOR g_3477 (.Z(w3688), .B(w3687), .A(w3037) );
	ym3438_SLATCH g_3478 (.Q(w3687), .D(w3040), .C(w3685), .nC(w3684) );
	ym3438_DLATCH_INV g_3479 (.nQ(w3686), .D(w3687), .C(w2545), .nC(w1150) );
	ym3438_NOT g_3480 (.A(w3686), .nZ(w2710) );
	ym3438_COMP_WE g_3481 (.A(w1140), .nZ(w3684), .Z(w3685) );
	ym3438_COMP_WE g_3482 (.A(w3035), .nZ(w3012), .Z(w3031) );
	ym3438_COMP_WE g_3483 (.A(w3034), .nZ(w3013), .Z(w3010) );
	ym3438_COMP_WE g_3484 (.A(w3033), .nZ(w3014), .Z(w3011) );
	ym3438_AND3 g_3485 (.B(w3014), .A(w3013), .C(w3012) );
	ym3438_AND3 g_3486 (.B(w3013), .A(w3014), .C(w3031) );
	ym3438_AND3 g_3487 (.Z(w3032), .B(w3010), .A(w3014), .C(w3012) );
	ym3438_AND3 g_3488 (.Z(w3683), .B(w3010), .A(w3014), .C(w3031) );
	ym3438_AND3 g_3489 (.Z(w3027), .B(w3013), .A(w3011), .C(w3012) );
	ym3438_AND3 g_3490 (.Z(w3028), .B(w3013), .A(w3031), .C(w3011) );
	ym3438_AND3 g_3491 (.Z(w3029), .B(w3010), .A(w3011), .C(w3012) );
	ym3438_AND3 g_3492 (.Z(w3030), .B(w3011), .A(w3031), .C(w3010) );
	ym3438_OR4 g_3493 (.Z(w3067), .B(w3029), .A(w3030), .C(w3028), .D(w3027) );
	ym3438_OR4 g_3494 (.Z(w3721), .B(w3028), .A(w3027), .C(w3029), .D(w3030) );
	ym3438_OR g_3495 (.Z(w3068), .B(w3030), .A(w3029) );
	ym3438_COMP_WE g_3496 (.A(w3030), .Z(w3926) );
	ym3438_OR4 g_3497 (.Z(w3720), .B(w3027), .A(w3683), .C(w3028), .D(w3029) );
	ym3438_OR g_3498 (.Z(w3719), .B(w3032), .A(w3683) );
	ym3438_OR4 g_3499 (.Z(w3718), .B(w3027), .A(w3028), .C(w3029), .D(w3030) );
	ym3438_OR3 g_3500 (.Z(w4142), .B(w3027), .A(w3683), .C(w3028) );
	ym3438_OR4 g_3501 (.Z(w4144), .B(w3683), .A(w3032), .C(w3029), .D(w3030) );
	ym3438_OR g_3502 (.Z(w4145), .B(w3029), .A(w3032) );
	ym3438_OR g_3503 (.Z(w4143), .B(w3683), .A(w3029) );
	ym3438_XOR g_3504 (.Z(w3033), .B(w3037), .A(w3036) );
	ym3438_XOR g_3505 (.Z(w3035), .B(w3037), .A(w3038) );
	ym3438_XOR g_3506 (.Z(w3034), .B(w3037), .A(w3039) );
	ym3438_AND g_3507 (.Z(w3717), .B(w1021), .A(w3069) );
	ym3438_AND g_3508 (.Z(w4343), .B(w1021), .A(w3071) );
	ym3438_AND g_3509 (.Z(w3716), .B(w1021), .A(w3070) );
	ym3438_AND g_3510 (.Z(w3711), .B(w1021), .A(w3072) );
	ym3438_AND g_3511 (.Z(w3712), .B(w1021), .A(w3074) );
	ym3438_AND g_3512 (.Z(w3713), .B(w1021), .A(w3073) );
	ym3438_AND g_3513 (.Z(w3715), .B(w1021), .A(w3714) );
	ym3438_SR_BIT g_3514 (.D(w3711), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .Q(w3047) );
	ym3438_SR_BIT g_3515 (.D(w3712), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .Q(w3050) );
	ym3438_SR_BIT g_3516 (.D(w3713), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .Q(w3046) );
	ym3438_SR_BIT g_3517 (.D(w3715), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .Q(w3044) );
	ym3438_SR_BIT g_3518 (.D(w3716), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .Q(w3042) );
	ym3438_SR_BIT g_3519 (.D(w4343), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .Q(w3041) );
	ym3438_SR_BIT g_3520 (.D(w3717), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .Q(w3040) );
	ym3438_NOT g_3521 (.A(w3690), .nZ(w1198) );
	ym3438_NOT g_3522 (.A(w3049), .nZ(w549) );
	ym3438_NOT g_3523 (.A(w3048), .nZ(w550) );
	ym3438_NOT g_3524 (.A(w3045), .nZ(w585) );
	ym3438_NOT g_3525 (.A(w3043), .nZ(w1197) );
	ym3438_NOT g_3526 (.A(w3688), .nZ(w1196) );
	ym3438_DLATCH_INV g_3527 (.nQ(w3076), .D(w3075), .C(w2546), .nC(w1149) );
	ym3438_AOI222222 g_3528 (.A2(1'b0), .B1(w3051), .A1(1'b0), .Z(w3075), .B2(w2677), .C1(w3710), .C2(w2536), .D1(w3056), .D2(w2629), .E2(w2539), .F1(1'b0), .F2(w2538), .E1(w3053) );
	ym3438_AOI222222 g_3529 (.A2(1'b0), .B1(w3106), .A1(1'b0), .Z(w3078), .B2(w2677), .C1(w3137), .C2(w2536), .D1(w3052), .D2(w2629), .E1(w3710), .E2(w2539), .F1(w3056), .F2(w2538) );
	ym3438_NOT g_3530 (.A(w3056), .nZ(w3053) );
	ym3438_NOT g_3531 (.A(w3052), .nZ(w3710) );
	ym3438_AOI222 g_3532 (.A2(w2551), .A1(w3056), .Z(w3175), .B2(w2550), .C1(1'b0), .C2(w2549), .B1(1'b0) );
	ym3438_DLATCH_INV g_3533 (.nQ(w3176), .D(w3175), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3534 (.nQ(w3077), .D(w3078), .C(w2546), .nC(w1149) );
	ym3438_AOI222222 g_3535 (.A2(1'b0), .B1(w3112), .A1(1'b0), .Z(w3138), .B2(w2677), .C1(w3862), .C2(w2536), .D1(w3051), .D2(w2629), .E2(w2539), .F1(w3052), .F2(w2538), .E1(w3137) );
	ym3438_NOT g_3536 (.A(w3051), .nZ(w3137) );
	ym3438_AOI222 g_3537 (.Z(w3174), .B2(w2550), .C1(1'b0), .C2(w2549), .B1(w3056), .A2(w2551), .A1(w3052) );
	ym3438_DLATCH_INV g_3538 (.nQ(w3177), .D(w3174), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3539 (.nQ(w3139), .D(w3138), .C(w2546), .nC(w1149) );
	ym3438_AOI222222 g_3540 (.A2(1'b0), .B1(w2958), .A1(1'b0), .Z(w3140), .B2(w2677), .C1(w3093), .C2(w2536), .D1(w3106), .D2(w2629), .E1(w3862), .E2(w2539), .F1(w3051), .F2(w2538) );
	ym3438_NOT g_3541 (.A(w3106), .nZ(w3862) );
	ym3438_AOI222 g_3542 (.A1(w3051), .Z(w3107), .C1(w3056), .C2(w2549), .B1(w3052), .B2(w2550), .A2(w2551) );
	ym3438_DLATCH_INV g_3543 (.nQ(w3108), .D(w3107), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3544 (.nQ(w3141), .D(w3140), .C(w2546), .nC(w1149) );
	ym3438_AOI222222 g_3545 (.A2(1'b0), .B1(w2964), .A1(1'b0), .Z(w3094), .B2(w2677), .C1(w3865), .C2(w2536), .D1(w3112), .D2(w2629), .E2(w2539), .F1(w3106), .F2(w2538), .E1(w3093) );
	ym3438_NOT g_3546 (.A(w3112), .nZ(w3093) );
	ym3438_AOI222 g_3547 (.Z(w3110), .B2(w2550), .C1(w3052), .C2(w2549), .B1(w3051), .A2(w2551), .A1(w3106) );
	ym3438_DLATCH_INV g_3548 (.nQ(w3109), .D(w3110), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3549 (.nQ(w3095), .D(w3094), .C(w2546), .nC(w1149) );
	ym3438_AOI222222 g_3550 (.A2(1'b0), .B1(w2899), .A1(1'b0), .Z(w3097), .B2(w2677), .C1(w2931), .C2(w2536), .D1(w2958), .D2(w2629), .E1(w3865), .E2(w2539), .F1(w3112), .F2(w2538) );
	ym3438_NOT g_3551 (.A(w2958), .nZ(w3865) );
	ym3438_AOI222 g_3552 (.A1(w3112), .Z(w2959), .C1(w3051), .C2(w2549), .B1(w3106), .B2(w2550), .A2(w2551) );
	ym3438_DLATCH_INV g_3553 (.nQ(w2962), .D(w2959), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3554 (.nQ(w3096), .D(w3097), .C(w2546), .nC(w1149) );
	ym3438_AOI222222 g_3555 (.A2(1'b0), .B1(w2905), .A1(1'b0), .Z(w2932), .B2(w2677), .C1(w3868), .C2(w2536), .D1(w2964), .D2(w2629), .E2(w2539), .F1(w2958), .F2(w2538), .E1(w2931) );
	ym3438_NOT g_3556 (.A(w2964), .nZ(w2931) );
	ym3438_AOI222 g_3557 (.Z(w2960), .B2(w2550), .C1(w3106), .C2(w2549), .B1(w3112), .A2(w2551), .A1(w2958) );
	ym3438_DLATCH_INV g_3558 (.nQ(w2961), .D(w2960), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3559 (.nQ(w2933), .D(w2932), .C(w2546), .nC(w1149) );
	ym3438_AOI222222 g_3560 (.A2(1'b0), .B1(w2834), .A1(1'b0), .Z(w2934), .B2(w2677), .C1(w2864), .C2(w2536), .D1(w2899), .D2(w2629), .E1(w3868), .E2(w2539), .F1(w2964), .F2(w2538) );
	ym3438_NOT g_3561 (.A(w2899), .nZ(w3868) );
	ym3438_AOI222 g_3562 (.A1(w2964), .Z(w2900), .C1(w3112), .C2(w2549), .B1(w2958), .B2(w2550), .A2(w2551) );
	ym3438_DLATCH_INV g_3563 (.nQ(w2901), .D(w2900), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3564 (.nQ(w2935), .D(w2934), .C(w2546), .nC(w1149) );
	ym3438_AOI222222 g_3565 (.A2(1'b0), .B1(w2840), .A1(1'b0), .Z(w2865), .B2(w2677), .C1(w3871), .C2(w2536), .D1(w2905), .D2(w2629), .E2(w2539), .F1(w2899), .F2(w2538), .E1(w2864) );
	ym3438_NOT g_3566 (.A(w2905), .nZ(w2864) );
	ym3438_AOI222 g_3567 (.Z(w2902), .B2(w2550), .C1(w2958), .C2(w2549), .B1(w2964), .A2(w2551), .A1(w2899) );
	ym3438_DLATCH_INV g_3568 (.nQ(w2903), .D(w2902), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3569 (.nQ(w2866), .D(w2865), .C(w2546), .nC(w1149) );
	ym3438_AOI222222 g_3570 (.A2(1'b0), .B1(w2764), .A1(1'b0), .Z(w2867), .B2(w2677), .C1(w2797), .C2(w2536), .D1(w2834), .D2(w2629), .E1(w3871), .E2(w2539), .F1(w2905), .F2(w2538) );
	ym3438_NOT g_3571 (.A(w2834), .nZ(w3871) );
	ym3438_AOI222 g_3572 (.A1(w2905), .Z(w2835), .C1(w2964), .C2(w2549), .B1(w2899), .B2(w2550), .A2(w2551) );
	ym3438_DLATCH_INV g_3573 (.nQ(w2836), .D(w2835), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3574 (.nQ(w2868), .D(w2867), .C(w2546), .nC(w1149) );
	ym3438_AOI222222 g_3575 (.A2(1'b0), .B1(w2725), .A1(1'b0), .Z(w2798), .B2(w2677), .C1(w3874), .C2(w2536), .D1(w2840), .D2(w2629), .E2(w2539), .F1(w2834), .F2(w2538), .E1(w2797) );
	ym3438_NOT g_3576 (.A(w2840), .nZ(w2797) );
	ym3438_AOI222 g_3577 (.Z(w2837), .B2(w2550), .C1(w2899), .C2(w2549), .B1(w2905), .A2(w2551), .A1(w2834) );
	ym3438_DLATCH_INV g_3578 (.nQ(w2838), .D(w2837), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3579 (.nQ(w2799), .D(w2798), .C(w2546), .nC(w1149) );
	ym3438_AOI222222 g_3580 (.A2(1'b0), .B1(w2694), .A1(1'b0), .Z(w2800), .B2(w2677), .C1(w2726), .C2(w2536), .D1(w2764), .D2(w2629), .E1(w3874), .E2(w2539), .F1(w2840), .F2(w2538) );
	ym3438_NOT g_3581 (.A(w2764), .nZ(w3874) );
	ym3438_AOI222 g_3582 (.A1(w2840), .Z(w2765), .C1(w2905), .C2(w2549), .B1(w2834), .B2(w2550), .A2(w2551) );
	ym3438_DLATCH_INV g_3583 (.nQ(w2766), .D(w2765), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3584 (.nQ(w2801), .D(w2800), .C(w2546), .nC(w1149) );
	ym3438_AOI222222 g_3585 (.A2(1'b0), .B1(w2662), .A1(1'b0), .Z(w2728), .B2(w2677), .C1(w3877), .C2(w2536), .D1(w2725), .D2(w2629), .E2(w2539), .F1(w2764), .F2(w2538), .E1(w2726) );
	ym3438_NOT g_3586 (.A(w2725), .nZ(w2726) );
	ym3438_AOI222 g_3587 (.Z(w2767), .B2(w2550), .C1(w2834), .C2(w2549), .B1(w2840), .A2(w2551), .A1(w2764) );
	ym3438_DLATCH_INV g_3588 (.nQ(w2768), .D(w2767), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3589 (.nQ(w2729), .D(w2728), .C(w2546), .nC(w1149) );
	ym3438_AOI222222 g_3590 (.A2(1'b0), .B1(w2643), .A1(1'b0), .Z(w2727), .B2(w2677), .C1(w2663), .C2(w2536), .D1(w2694), .D2(w2629), .E1(w3877), .E2(w2539), .F1(w2725), .F2(w2538) );
	ym3438_NOT g_3591 (.A(w2694), .nZ(w3877) );
	ym3438_AOI222 g_3592 (.A1(w2725), .Z(w2695), .C1(w2840), .C2(w2549), .B1(w2764), .B2(w2550), .A2(w2551) );
	ym3438_DLATCH_INV g_3593 (.nQ(w2696), .D(w2695), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3594 (.nQ(w2730), .D(w2727), .C(w2546), .nC(w1149) );
	ym3438_AOI222222 g_3595 (.A2(1'b0), .B1(w2581), .A1(1'b0), .Z(w2665), .B2(w2677), .C1(w3880), .C2(w2536), .D1(w2662), .D2(w2629), .E2(w2539), .F1(w2694), .F2(w2538), .E1(w2663) );
	ym3438_NOT g_3596 (.A(w2662), .nZ(w2663) );
	ym3438_AOI222 g_3597 (.Z(w2697), .B2(w2550), .C1(w2764), .C2(w2549), .B1(w2725), .A2(w2551), .A1(w2694) );
	ym3438_DLATCH_INV g_3598 (.nQ(w2698), .D(w2697), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3599 (.nQ(w2666), .D(w2665), .C(w2546), .nC(w1149) );
	ym3438_AOI222222 g_3600 (.A2(1'b0), .B1(1'b0), .A1(1'b0), .Z(w2664), .B2(w2677), .C1(w2619), .C2(w2536), .D1(w2643), .D2(w2629), .E1(w3880), .E2(w2539), .F1(w2662), .F2(w2538) );
	ym3438_NOT g_3601 (.A(w2643), .nZ(w3880) );
	ym3438_AOI222 g_3602 (.A1(w2662), .Z(w2644), .C1(w2725), .C2(w2549), .B1(w2694), .B2(w2550), .A2(w2551) );
	ym3438_DLATCH_INV g_3603 (.nQ(w2645), .D(w2644), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3604 (.nQ(w2667), .D(w2664), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3605 (.nQ(w2647), .D(w2646), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3606 (.nQ(w2621), .D(w2620), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3607 (.nQ(w2583), .D(w2582), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3608 (.nQ(w2624), .D(w2623), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3609 (.nQ(w2584), .D(w2579), .C(w2546), .nC(w1149) );
	ym3438_DLATCH_INV g_3610 (.nQ(w3194), .D(w3193), .C(w2546), .nC(w1149) );
	ym3438_AOI2222 g_3611 (.A2(w2536), .B1(w2581), .A1(1'b1), .Z(w2620), .B2(w2629), .C1(w2619), .C2(w2539), .D1(w2643), .D2(w2538) );
	ym3438_AOI222 g_3612 (.A2(w2536), .B1(1'b1), .A1(1'b1), .Z(w2623), .B2(w2539), .C1(w2581), .C2(w2538) );
	ym3438_AOI22 g_3613 (.A2(1'b1), .A1(w2539), .Z(w3193), .B2(1'b1), .B1(w2536) );
	ym3438_AOI222 g_3614 (.A2(w2551), .B1(w2581), .A1(1'b0), .Z(w2579), .B2(w2550), .C1(w2643), .C2(w2549) );
	ym3438_AOI222 g_3615 (.A2(w2551), .A1(w2581), .Z(w2582), .B2(w2550), .C1(w2662), .C2(w2549), .B1(w2643) );
	ym3438_AOI222 g_3616 (.Z(w2646), .B2(w2550), .C1(w2694), .C2(w2549), .B1(w2662), .A2(w2551), .A1(w2643) );
	ym3438_NOT g_3617 (.A(w2581), .nZ(w2619) );
	ym3438_NOT g_3618 (.A(w3190), .nZ(w2547) );
	ym3438_NOT g_3619 (.A(w3882), .nZ(w2548) );
	ym3438_NOT g_3620 (.A(w3190), .nZ(w3882) );
	ym3438_NOT g_3621 (.A(w3883), .nZ(w3190) );
	ym3438_AND g_3622 (.Z(w2631), .B(w2564), .A(w2613) );
	ym3438_OR g_3623 (.Z(w2605), .B(w2564), .A(w2613) );
	ym3438_NOT g_3624 (.A(w3969), .nZ(w4366) );
	ym3438_SR_BIT g_3625 (.Q(w4012), .D(w333), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_COMP_STR g_3626 (.A(w4012), .Z(w2603) );
	ym3438_COMP_STR g_3627 (.A(w4011), .Z(w2602) );
	ym3438_SR_BIT g_3628 (.Q(w4011), .D(w2603), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_AND3 g_3629 (.B(w4007), .A(w2606), .C(w4006) );
	ym3438_OR3 g_3630 (.Z(w2614), .B(w2609), .A(w2616), .C(w2607) );
	ym3438_AND3 g_3631 (.Z(w4010), .B(w4007), .A(w2606), .C(w2608) );
	ym3438_OR4 g_3632 (.Z(w2615), .B(w2607), .A(w4010), .C(w2616), .D(w2632) );
	ym3438_AND3 g_3633 (.Z(w2607), .B(w2610), .A(w2606), .C(w4006) );
	ym3438_AND3 g_3634 (.Z(w2632), .B(w2612), .A(w2610), .C(w2608) );
	ym3438_AND3 g_3635 (.Z(w2616), .B(w2610), .A(w2612), .C(w4006) );
	ym3438_AND3 g_3636 (.Z(w4008), .B(w4007), .A(w2608), .C(w2612) );
	ym3438_OR3 g_3637 (.Z(w2618), .B(w2616), .A(w4008), .C(w2632) );
	ym3438_AND3 g_3638 (.Z(w2609), .B(w4007), .A(w2612), .C(w4006) );
	ym3438_AND3 g_3639 (.Z(w4009), .B(w2606), .A(w2608), .C(w2610) );
	ym3438_OR3 g_3640 (.Z(w2617), .B(w2609), .A(w2632), .C(w4009) );
	ym3438_AND g_3641 (.Z(w2611), .B(w3982), .A(w2660) );
	ym3438_AND g_3642 (.Z(w3984), .B(w3983), .A(w2660) );
	ym3438_COMP_WE g_3643 (.A(w3984), .nZ(w4006), .Z(w2608) );
	ym3438_COMP_WE g_3644 (.A(w2611), .nZ(w4007), .Z(w2610) );
	ym3438_COMP_WE g_3645 (.A(w2633), .nZ(w2606), .Z(w2612) );
	ym3438_FA g_3646 (.CO(w2568), .S(w2569), .CI(w3985), .A(w2605), .B(1'b0) );
	ym3438_FA g_3647 (.CO(w3985), .S(w2570), .CI(w4003), .A(1'b0), .B(w2659) );
	ym3438_FA g_3648 (.CO(w4003), .S(w2571), .CI(w4004), .A(w2564), .B(w2680) );
	ym3438_FA g_3649 (.CO(w4004), .S(w2633), .CI(1'b1), .A(w2631), .B(w2658) );
	ym3438_NAND3 g_3650 (.Z(w2660), .B(w2658), .A(w2659), .C(w2680) );
	ym3438_SR_BIT g_3651 (.Q(w2680), .D(w806), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_SR_BIT g_3652 (.Q(w806), .D(w1132), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_SR_BIT g_3653 (.Q(w2659), .D(w1145), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_SR_BIT g_3654 (.Q(w1145), .D(w1133), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_SR_BIT g_3655 (.Q(w2658), .D(w808), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_SR_BIT g_3656 (.Q(w808), .D(w1131), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_SR_BIT g_3657 (.Q(w3983), .D(w1144), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_SR_BIT g_3658 (.Q(w1144), .D(w1129), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_SR_BIT g_3659 (.Q(w3982), .D(w783), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_SR_BIT g_3660 (.Q(w783), .D(w1130), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_FA g_3661 (.CO(w3999), .S(w2712), .CI(w2679), .A(w2678), .B(w2711) );
	ym3438_FA g_3662 (.CO(w3995), .S(w2743), .CI(w3999), .A(w2678), .B(w2742) );
	ym3438_NOT g_3663 (.A(w3980), .nZ(w2749) );
	ym3438_SR_BIT g_3664 (.Q(w3998), .D(w1123), .nC1(w1150), .nC2(w1149), .C1(w2545), .C2(w2546) );
	ym3438_DLATCH_INV g_3665 (.nQ(w2721), .D(w2720), .nC(w1149), .C(w2546) );
	ym3438_XNOR g_3666 (.Z(w2720), .B(w2710), .A(w2718) );
	ym3438_AON222 g_3667 (.A2(w1141), .A1(w2748), .Z(w2718), .B2(w1138), .C1(w1136), .C2(1'b0), .B1(w2716) );
	ym3438_FA g_3668 (.CO(w2716), .S(w2748), .CI(w3997), .A(w2745), .B(w2714) );
	ym3438_DLATCH_INV g_3669 (.nQ(w2714), .D(w2713), .nC(w1150), .C(w2545) );
	ym3438_DLATCH_INV g_3670 (.nQ(w2745), .D(w2744), .nC(w1150), .C(w2545) );
	ym3438_AOI22 g_3671 (.A2(w1118), .B1(1'b0), .A1(w1135), .Z(w2713), .B2(w2852) );
	ym3438_AOI22 g_3672 (.A2(1'b0), .B1(1'b0), .A1(w1134), .Z(w2744), .B2(w3151) );
	ym3438_NOT g_3673 (.A(w4000), .nZ(w1142) );
	ym3438_DLATCH_INV g_3674 (.nQ(w4000), .D(w2743), .nC(w1150), .C(w2545) );
	ym3438_SR_BIT g_3675 (.Q(w2742), .D(w1120), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_FA g_3676 (.CO(w3993), .S(w2783), .CI(w3995), .A(w2678), .B(w2782) );
	ym3438_NOT g_3677 (.A(w3979), .nZ(w2756) );
	ym3438_SR_BIT g_3678 (.Q(w2752), .D(w1124), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3679 (.nQ(w2791), .D(w2790), .C(w2546), .nC(w1149) );
	ym3438_XNOR g_3680 (.Z(w2790), .B(w2710), .A(w2789) );
	ym3438_AON222 g_3681 (.A2(w1141), .A1(w2788), .Z(w2789), .B2(w1138), .C1(w1136), .C2(w2716), .B1(w2748) );
	ym3438_FA g_3682 (.CO(w3997), .S(w2788), .CI(w3991), .A(w2747), .B(w2786) );
	ym3438_DLATCH_INV g_3683 (.nQ(w2786), .D(w2785), .C(w2545), .nC(w1150) );
	ym3438_DLATCH_INV g_3684 (.nQ(w2747), .D(w2746), .C(w2545), .nC(w1150) );
	ym3438_AOI22 g_3685 (.A2(w1119), .B1(w1118), .A1(w1135), .Z(w2785), .B2(w2852) );
	ym3438_AOI22 g_3686 (.A2(1'b0), .B1(w1118), .A1(w1134), .Z(w2746), .B2(w3151) );
	ym3438_NOT g_3687 (.A(w3994), .nZ(w1143) );
	ym3438_DLATCH_INV g_3688 (.nQ(w3994), .D(w2783), .C(w2545), .nC(w1150) );
	ym3438_SR_BIT g_3689 (.Q(w2782), .D(w1119), .nC1(w1150), .nC2(w1149), .C1(w2545), .C2(w2546) );
	ym3438_FA g_3690 (.S(w2781), .CI(w3993), .A(w2678), .B(w2780) );
	ym3438_NOT g_3691 (.A(w3977), .nZ(w2823) );
	ym3438_SR_BIT g_3692 (.Q(w2819), .D(w1125), .nC1(w1150), .nC2(w1149), .C1(w2545), .C2(w2546) );
	ym3438_DLATCH_INV g_3693 (.nQ(w2794), .D(w2793), .nC(w1149), .C(w2546) );
	ym3438_XNOR g_3694 (.Z(w2793), .B(w2710), .A(w2792) );
	ym3438_AON222 g_3695 (.A2(w1141), .A1(w2817), .Z(w2792), .B2(w1138), .C1(w1136), .C2(w2748), .B1(w2788) );
	ym3438_FA g_3696 (.CO(w3991), .S(w2817), .CI(w3990), .A(w2815), .B(w2787) );
	ym3438_DLATCH_INV g_3697 (.nQ(w2787), .D(w2784), .nC(w1150), .C(w2545) );
	ym3438_DLATCH_INV g_3698 (.nQ(w2815), .D(w2813), .nC(w1150), .C(w2545) );
	ym3438_AOI22 g_3699 (.A2(w1120), .B1(w1119), .A1(w1135), .Z(w2784), .B2(w2852) );
	ym3438_AOI22 g_3700 (.A1(w1134), .Z(w2813), .B2(w3151), .A2(w1118), .B1(w1119) );
	ym3438_NOT g_3701 (.A(w3992), .nZ(w2812) );
	ym3438_DLATCH_INV g_3702 (.nQ(w3992), .D(w2781), .nC(w1150), .C(w2545) );
	ym3438_SR_BIT g_3703 (.Q(w2780), .D(w1118), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3704 (.nQ(w3977), .D(w2821), .nC(w1150), .C(w2545) );
	ym3438_DLATCH_INV g_3705 (.nQ(w3979), .D(w2753), .C(w2545), .nC(w1150) );
	ym3438_DLATCH_INV g_3706 (.nQ(w3980), .D(w2755), .nC(w1150), .C(w2545) );
	ym3438_FA g_3707 (.CO(w2795), .S(w2821), .CI(w2820), .A(w2794), .B(w2819) );
	ym3438_FA g_3708 (.CO(w2754), .S(w2753), .CI(w2795), .A(w2791), .B(w2752) );
	ym3438_FA g_3709 (.CO(w2723), .S(w2755), .CI(w2754), .A(w2721), .B(w3998) );
	ym3438_FA g_3710 (.CO(w2679), .S(w2682), .CI(w2723), .A(w2722), .B(w2681) );
	ym3438_NOT g_3711 (.A(w3981), .nZ(w2684) );
	ym3438_DLATCH_INV g_3712 (.nQ(w3981), .D(w2682), .C(w2545), .nC(w1150) );
	ym3438_NOT g_3713 (.A(w3975), .nZ(w2824) );
	ym3438_SR_BIT g_3714 (.Q(w2818), .D(w1126), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3715 (.nQ(w2858), .D(w2857), .C(w2546), .nC(w1149) );
	ym3438_XNOR g_3716 (.Z(w2857), .B(w2710), .A(w2856) );
	ym3438_AON222 g_3717 (.A2(w1141), .A1(w2855), .Z(w2856), .B2(w1138), .C1(w1136), .C2(w2788), .B1(w2817) );
	ym3438_FA g_3718 (.CO(w3990), .S(w2855), .CI(w3989), .A(w2816), .B(w2851) );
	ym3438_DLATCH_INV g_3719 (.nQ(w2851), .D(w2850), .C(w2545), .nC(w1150) );
	ym3438_DLATCH_INV g_3720 (.nQ(w2816), .D(w2814), .C(w2545), .nC(w1150) );
	ym3438_AOI22 g_3721 (.A2(w1121), .B1(w1120), .A1(w1135), .Z(w2850), .B2(w2852) );
	ym3438_AOI22 g_3722 (.A2(w1119), .B1(w1120), .A1(w1134), .Z(w2814), .B2(w3151) );
	ym3438_DLATCH_INV g_3723 (.nQ(w3975), .D(w2822), .C(w2545), .nC(w1150) );
	ym3438_FA g_3724 (.CO(w2820), .S(w2822), .CI(w2859), .A(w2858), .B(w2818) );
	ym3438_NOT g_3725 (.A(w3974), .nZ(w2889) );
	ym3438_SR_BIT g_3726 (.Q(w3986), .D(w1127), .nC1(w1150), .nC2(w1149), .C1(w2545), .C2(w2546) );
	ym3438_DLATCH_INV g_3727 (.nQ(w2862), .D(w2861), .nC(w1149), .C(w2546) );
	ym3438_XNOR g_3728 (.Z(w2861), .B(w2710), .A(w2860) );
	ym3438_AON222 g_3729 (.A2(w1141), .A1(w2883), .Z(w2860), .B2(w1138), .C1(w1136), .C2(w2817), .B1(w2855) );
	ym3438_FA g_3730 (.CO(w3989), .S(w2883), .CI(w3988), .A(w2881), .B(w2854) );
	ym3438_DLATCH_INV g_3731 (.nQ(w2854), .D(w2853), .nC(w1150), .C(w2545) );
	ym3438_DLATCH_INV g_3732 (.nQ(w2881), .D(w2882), .nC(w1150), .C(w2545) );
	ym3438_AOI22 g_3733 (.A2(w1122), .B1(w1121), .A1(w1135), .Z(w2853), .B2(w2852) );
	ym3438_AOI22 g_3734 (.A1(w1134), .Z(w2882), .B2(w3151), .A2(w1120), .B1(w1121) );
	ym3438_DLATCH_INV g_3735 (.nQ(w3974), .D(w2886), .nC(w1150), .C(w2545) );
	ym3438_FA g_3736 (.CO(w2859), .S(w2886), .CI(w2885), .A(w2862), .B(w3986) );
	ym3438_NOT g_3737 (.A(w3972), .nZ(w2888) );
	ym3438_SR_BIT g_3738 (.Q(w2884), .D(w1128), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3739 (.nQ(w2927), .D(w3987), .C(w2546), .nC(w1149) );
	ym3438_XNOR g_3740 (.Z(w3987), .B(w2710), .A(w2923) );
	ym3438_AON222 g_3741 (.A2(w1141), .A1(w2922), .Z(w2923), .B2(w1138), .C1(w1136), .C2(w2855), .B1(w2883) );
	ym3438_FA g_3742 (.CO(w3988), .S(w2922), .CI(w3966), .A(w2880), .B(w2921) );
	ym3438_DLATCH_INV g_3743 (.nQ(w2921), .D(w2920), .C(w2545), .nC(w1150) );
	ym3438_DLATCH_INV g_3744 (.nQ(w2880), .D(w2879), .C(w2545), .nC(w1150) );
	ym3438_AOI22 g_3745 (.A2(w1123), .B1(w1122), .A1(w1135), .Z(w2920), .B2(w2852) );
	ym3438_AOI22 g_3746 (.A2(w1121), .B1(w1122), .A1(w1134), .Z(w2879), .B2(w3151) );
	ym3438_DLATCH_INV g_3747 (.nQ(w3972), .D(w2887), .C(w2545), .nC(w1150) );
	ym3438_FA g_3748 (.CO(w2885), .S(w2887), .CI(w2928), .A(w2927), .B(w2884) );
	ym3438_NOT g_3749 (.A(w3964), .nZ(w2929) );
	ym3438_DLATCH_INV g_3750 (.nQ(w2926), .D(w2925), .nC(w1149), .C(w2546) );
	ym3438_XNOR g_3751 (.Z(w2925), .B(w2710), .A(w2924) );
	ym3438_AON222 g_3752 (.A2(w1141), .A1(w3965), .Z(w2924), .B2(w1138), .C1(w1136), .C2(w2883), .B1(w2922) );
	ym3438_FA g_3753 (.CO(w3966), .S(w3965), .CI(1'b0), .A(w2946), .B(w2919) );
	ym3438_DLATCH_INV g_3754 (.nQ(w2919), .D(w2918), .nC(w1150), .C(w2545) );
	ym3438_DLATCH_INV g_3755 (.nQ(w2946), .D(w2945), .nC(w1150), .C(w2545) );
	ym3438_AOI22 g_3756 (.A2(w1124), .B1(w1123), .A1(w1135), .Z(w2918), .B2(w2852) );
	ym3438_AOI22 g_3757 (.A2(w1122), .B1(w1123), .A1(w1134), .Z(w2945), .B2(w3151) );
	ym3438_DLATCH_INV g_3758 (.nQ(w3964), .D(w2948), .nC(w1150), .C(w2545) );
	ym3438_FA g_3759 (.CO(w2928), .S(w2948), .CI(w3963), .A(w2926), .B(1'b0) );
	ym3438_SR_BIT g_3760 (.Q(w2711), .D(w1121), .nC1(w1150), .nC2(w1149), .C1(w2545), .C2(w2546) );
	ym3438_DLATCH_INV g_3761 (.nQ(w4002), .D(w2712), .C(w2545), .nC(w1150) );
	ym3438_DLATCH_INV g_3762 (.nQ(w2678), .D(w2715), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3763 (.A(w4002), .nZ(w3970) );
	ym3438_NOT g_3764 (.A(w2710), .nZ(w2715) );
	ym3438_SR_BIT g_3765 (.Q(w2681), .D(w1122), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149) );
	ym3438_DLATCH_INV g_3766 (.nQ(w2722), .D(w2719), .C(w2546), .nC(w1149) );
	ym3438_XNOR g_3767 (.Z(w2719), .B(w2710), .A(w2717) );
	ym3438_AON222 g_3768 (.A2(w1141), .A1(w2716), .Z(w2717), .B2(w1138), .C1(w1136), .C2(1'b0), .B1(1'b0) );
	ym3438_NOT g_3769 (.A(w3971), .nZ(w1149) );
	ym3438_NOT g_3770 (.A(w3973), .nZ(w2546) );
	ym3438_NOT g_3771 (.A(w3976), .nZ(w2545) );
	ym3438_NOT g_3772 (.A(w3978), .nZ(w1150) );
	ym3438_NOT g_3773 (.A(w217), .nZ(w3971) );
	ym3438_NOT g_3774 (.A(w216), .nZ(w3973) );
	ym3438_NOT g_3775 (.A(w213), .nZ(w3976) );
	ym3438_NOT g_3776 (.A(w212), .nZ(w3978) );
	ym3438_SR_BIT g_3777 (.Q(w3087), .D(w847), .nC1(w1150), .nC2(w1149), .C1(w2545), .C2(w2546) );
	ym3438_EDGE_DET g_3778 (.Q(w1140), .D(w3087), .C1(w2545), .nC1(w1150) );
	ym3438_OR g_3779 (.Z(w3955), .B(w1139), .A(w847) );
	ym3438_HA g_3780 (.CO(w3956), .S(w3952), .A(w2981), .B(w3955) );
	ym3438_HA g_3781 (.CO(w3957), .S(w3953), .A(w2982), .B(w3956) );
	ym3438_HA g_3782 (.S(w3940), .A(w2985), .B(w3961) );
	ym3438_HA g_3783 (.CO(w3961), .S(w3943), .A(w2986), .B(w3960) );
	ym3438_HA g_3784 (.CO(w3960), .S(w3945), .A(w2987), .B(w3959) );
	ym3438_HA g_3785 (.CO(w3959), .S(w3947), .A(w2984), .B(w3958) );
	ym3438_HA g_3786 (.CO(w3958), .S(w3954), .A(w2983), .B(w3957) );
	ym3438_XOR g_3787 (.Z(w3939), .A(w2604), .B(w2603) );
	ym3438_SR_BIT g_3788 (.D(w3939), .nC1(w1150), .nC2(w1149), .C1(w2545), .C2(w2546), .Q(w3091) );
	ym3438_DLATCH_INV g_3789 (.nQ(w3962), .D(w2710), .C(w2546), .nC(w1149) );
	ym3438_NOT g_3790 (.A(w3962), .nZ(w3963) );
	ym3438_AON222 g_3791 (.A2(w2888), .A1(w2572), .Z(w2988), .B2(w2741), .C1(1'b0), .C2(w2553), .B1(w2929) );
	ym3438_NOT g_3792 (.A(w3901), .nZ(w3051) );
	ym3438_DLATCH_INV g_3793 (.nQ(w3901), .D(w2996), .C(w2545), .nC(w1150) );
	ym3438_FA g_3794 (.CO(w2994), .S(w2996), .CI(w3136), .A(w3135), .B(w2992) );
	ym3438_DLATCH_INV g_3795 (.nQ(w2992), .D(w2991), .C(w2546), .nC(w1149) );
	ym3438_AOI22 g_3796 (.A2(w2548), .A1(w2989), .Z(w2991), .B2(w2547), .B1(w2890) );
	ym3438_NOT g_3797 (.A(w3906), .nZ(w3052) );
	ym3438_DLATCH_INV g_3798 (.nQ(w3906), .D(w3171), .C(w2545), .nC(w1150) );
	ym3438_FA g_3799 (.CO(w3136), .S(w3171), .CI(w3170), .A(w3134), .B(w3169) );
	ym3438_DLATCH_INV g_3800 (.nQ(w3169), .D(w3165), .C(w2546), .nC(w1149) );
	ym3438_AOI22 g_3801 (.A2(w2548), .A1(w3164), .Z(w3165), .B2(w2547), .B1(w2950) );
	ym3438_NOT g_3802 (.A(w3900), .nZ(w3056) );
	ym3438_DLATCH_INV g_3803 (.nQ(w3900), .D(w3172), .C(w2545), .nC(w1150) );
	ym3438_FA g_3804 (.CO(w3170), .S(w3172), .CI(w2602), .A(w3167), .B(w3168) );
	ym3438_DLATCH_INV g_3805 (.nQ(w3168), .D(w3166), .C(w2546), .nC(w1149) );
	ym3438_SR_BIT g_3806 (.D(w3938), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .Q(w3090) );
	ym3438_SR_BIT g_3807 (.D(w3941), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .Q(w2985) );
	ym3438_XOR g_3808 (.Z(w3938), .A(w2559), .B(w2603) );
	ym3438_AND g_3809 (.Z(w3941), .B(w3088), .A(w3940) );
	ym3438_AND g_3810 (.Z(w3942), .B(w3088), .A(w3943) );
	ym3438_AND g_3811 (.Z(w3944), .B(w3088), .A(w3945) );
	ym3438_AND g_3812 (.Z(w3946), .B(w3088), .A(w3947) );
	ym3438_AND g_3813 (.Z(w3948), .B(w3088), .A(w3954) );
	ym3438_AND g_3814 (.Z(w3949), .B(w3088), .A(w3953) );
	ym3438_AND g_3815 (.Z(w3950), .B(w3088), .A(w3952) );
	ym3438_NOR g_3816 (.Z(w3088), .B(w2980), .A(w3951) );
	ym3438_NOT g_3817 (.A(w214), .nZ(w3951) );
	ym3438_SR_BIT g_3818 (.D(w3949), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .Q(w2982) );
	ym3438_SR_BIT g_3819 (.D(w3950), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .Q(w2981) );
	ym3438_SR_BIT g_3820 (.D(w3948), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .Q(w2983) );
	ym3438_SR_BIT g_3821 (.D(w3946), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .Q(w2984) );
	ym3438_SR_BIT g_3822 (.D(w3942), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .Q(w2986) );
	ym3438_SR_BIT g_3823 (.D(w3944), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .Q(w2987) );
	ym3438_NAND g_3824 (.Z(w3166), .B(w2547), .A(w2949) );
	ym3438_AND g_3825 (.Z(w3164), .B(1'b0), .A(w2572) );
	ym3438_AON22 g_3826 (.A2(w2572), .A1(w2929), .Z(w2989), .B2(w2741), .B1(1'b0) );
	ym3438_XOR g_3827 (.Z(w3937), .B(w2603), .A(w2560) );
	ym3438_AND3 g_3828 (.Z(w3152), .B(w3158), .A(w3126), .C(w3124) );
	ym3438_OR g_3829 (.Z(w3154), .B(w2979), .A(w2978) );
	ym3438_AND3 g_3830 (.Z(w3157), .B(w3125), .A(w3159), .C(w3149) );
	ym3438_AND3 g_3831 (.Z(w3156), .B(w3125), .A(w3159), .C(w3124) );
	ym3438_AND3 g_3832 (.Z(w3155), .B(w3158), .A(w3126), .C(w3149) );
	ym3438_AND3 g_3833 (.Z(w3923), .B(w3158), .A(w3159), .C(w3124) );
	ym3438_AND3 g_3834 (.Z(w3131), .B(w2983), .A(w2981), .C(w3929) );
	ym3438_AND g_3835 (.Z(w3133), .B(w2984), .A(w3930) );
	ym3438_AND4 g_3836 (.Z(w3931), .B(w2986), .A(w2984), .C(w2983), .D(w4149) );
	ym3438_AND6 g_3837 (.Z(w3932), .B(w2983), .A(w2984), .C(w2982), .D(w2987), .E(w2986), .F(w4148) );
	ym3438_AND4 g_3838 (.Z(w4147), .B(w2982), .A(w2985), .C(w2981), .D(w3934) );
	ym3438_AND5 g_3839 (.Z(w3132), .B(w2982), .A(w2981), .C(w2983), .D(w2985), .E(w4146) );
	ym3438_AND5 g_3840 (.Z(w3933), .B(w2983), .A(w2981), .C(w2984), .D(w2985), .E(w3935) );
	ym3438_AND5 g_3841 (.Z(w3130), .B(w2984), .A(w2983), .C(w2986), .D(w2985), .E(w3936) );
	ym3438_SR_BIT g_3842 (.D(w3937), .nC1(w1150), .nC2(w1149), .C1(w2545), .C2(w2546), .Q(w3135) );
	ym3438_SR_BIT g_3843 (.D(w3928), .C1(w2545), .C2(w2546), .nC1(w1150), .nC2(w1149), .Q(w3134) );
	ym3438_SR_BIT g_3844 (.D(w3915), .nC1(w1150), .nC2(w1149), .C1(w2545), .C2(w2546), .Q(w3167) );
	ym3438_DLATCH_INVS g_3845 (.nQ(w1138), .D(w2976), .C(w2545), .nC(w1150) );
	ym3438_DLATCH_INVS g_3846 (.nQ(w1141), .D(w2977), .C(w2545), .nC(w1150) );
	ym3438_DLATCH_INVS g_3847 (.nQ(w1136), .D(w3154), .C(w2545), .nC(w1150) );
	ym3438_AND3 g_3848 (.Z(w2979), .B(w3125), .A(w3126), .C(w3149) );
	ym3438_AND3 g_3849 (.Z(w2978), .B(w3125), .A(w3126), .C(w3124) );
	ym3438_NOT g_3850 (.A(w2979), .nZ(w2976) );
	ym3438_NOT g_3851 (.A(w2978), .nZ(w2977) );
	ym3438_NOT g_3852 (.A(w4364), .nZ(w3151) );
	ym3438_NOT g_3853 (.A(w3922), .nZ(w1134) );
	ym3438_NOT g_3854 (.A(w3927), .nZ(w1135) );
	ym3438_NOT g_3855 (.A(w3925), .nZ(w2852) );
	ym3438_XOR g_3856 (.Z(w3915), .B(w2603), .A(w3150) );
	ym3438_XOR g_3857 (.Z(w3928), .B(w2603), .A(w3123) );
	ym3438_AND3 g_3858 (.Z(w3929), .B(w3129), .A(w3160), .C(w3128) );
	ym3438_AND3 g_3859 (.Z(w3930), .B(w3129), .A(w3160), .C(w3162) );
	ym3438_AND3 g_3860 (.Z(w4149), .B(w3161), .A(w3160), .C(w3128) );
	ym3438_AND3 g_3861 (.Z(w4148), .B(w3161), .A(w3160), .C(w3162) );
	ym3438_OR8 g_3862 (.Z(w2980), .B(w3933), .A(w3130), .C(w3132), .D(w4147), .E(w3932), .F(w3931), .G(w3133), .H(w3131) );
	ym3438_AND3 g_3863 (.Z(w3934), .B(w3129), .A(w3127), .C(w3128) );
	ym3438_AND3 g_3864 (.Z(w4146), .B(w3129), .A(w3127), .C(w3162) );
	ym3438_AND3 g_3865 (.Z(w3935), .B(w3161), .A(w3127), .C(w3128) );
	ym3438_AND3 g_3866 (.Z(w3936), .B(w3161), .A(w3127), .C(w3162) );
	ym3438_COMP_WE g_3867 (.A(w1044), .nZ(w3162), .Z(w3128) );
	ym3438_COMP_WE g_3868 (.A(w1045), .nZ(w3161), .Z(w3129) );
	ym3438_COMP_WE g_3869 (.A(w1137), .nZ(w3127), .Z(w3160) );
	ym3438_OR g_3870 (.Z(w3153), .B(w3152), .A(w3154) );
	ym3438_NAND g_3871 (.Z(w4364), .B(w3153), .A(w3926) );
	ym3438_AOI22 g_3872 (.A2(w3155), .A1(w3926), .Z(w3927), .B2(w3153), .B1(w3067) );
	ym3438_AOI2222 g_3873 (.A2(w3157), .A1(w3068), .Z(w3925), .B2(w3156), .C1(w3155), .C2(w3720), .B1(w3721), .D1(w3719), .D2(w3153) );
	ym3438_AOI222222 g_3874 (.A2(w4143), .B1(w3155), .A1(w3153), .Z(w3922), .B2(w4145), .C1(w3156), .C2(w4144), .D1(w3157), .D2(w4142), .E1(w3923), .E2(w3718), .F1(1'b0), .F2(1'b0) );
	ym3438_HA g_3875 (.S(w3069), .A(w3040), .B(w3921) );
	ym3438_HA g_3876 (.CO(w3921), .S(w3071), .A(w3041), .B(w3920) );
	ym3438_HA g_3877 (.CO(w3920), .S(w3070), .A(w3042), .B(w3919) );
	ym3438_HA g_3878 (.CO(w3916), .S(w3072), .A(w3047), .B(w2980) );
	ym3438_HA g_3879 (.CO(w3917), .S(w3074), .A(w3050), .B(w3916) );
	ym3438_HA g_3880 (.CO(w3918), .S(w3073), .A(w3046), .B(w3917) );
	ym3438_HA g_3881 (.CO(w3919), .S(w3714), .A(w3044), .B(w3918) );
	ym3438_COMP_WE g_3882 (.A(w1148), .nZ(w3149), .Z(w3124) );
	ym3438_COMP_WE g_3883 (.A(w1147), .nZ(w3158), .Z(w3125) );
	ym3438_COMP_WE g_3884 (.A(w1146), .nZ(w3159), .Z(w3126) );
	ym3438_NOT g_3885 (.A(w1112), .nZ(w3288) );
	ym3438_NOT g_3886 (.A(w1115), .nZ(w3290) );
	ym3438_AON22 g_3887 (.A2(w3891), .A1(w2618), .Z(w2559), .B2(w3893), .B1(w3893) );
	ym3438_COMP_WE_STRONG g_7A (.A(w1306), .Z(w1309), .nZ(w1341) );
	ym3438_COMP_WE_STRONG g_7B (.A(w1338), .Z(w1310), .nZ(w830) );
	ym3438_BUF2 g_2 (.A(w1306), .Z(w1307) );
	ym3438_NOT g_2548 (.A(w2442), .nZ(w3270) );
	ym3438_NOT g_2560 (.A(w2440), .nZ(w3278) );
	ym3438_NOR g_2495 (.Z(w3227), .B(w1111), .A(w3226) );
	ym3438_NOR g_2503 (.Z(w3233), .B(w1111), .A(w3232) );
	ym3438_NAND g_1100A (.A(w4426), .Z(w1865), .B(w1863) );
endmodule // ym3438

// ERROR: floating wire w21
// ERROR: conflicting wire w108
// ERROR: conflicting wire w112
// ERROR: conflicting wire w123
// ERROR: conflicting wire w132
// ERROR: floating wire w421
// ERROR: floating wire w525
// ERROR: floating wire w556
// ERROR: floating wire w563
// ERROR: floating wire w620
// ERROR: floating wire w680
// ERROR: floating wire w716
// ERROR: conflicting wire w958
// ERROR: conflicting wire w959
// ERROR: conflicting wire w960
// ERROR: conflicting wire w961
// ERROR: floating wire w968
// ERROR: floating wire w1003
// ERROR: conflicting wire w1078
// ERROR: floating wire w1102
// ERROR: conflicting wire w1155
// ERROR: conflicting wire w1156
// ERROR: floating wire w1336
// ERROR: floating wire w1351
// ERROR: floating wire w1368
// ERROR: floating wire w1386
// ERROR: floating wire w1717
// ERROR: floating wire w1889
// ERROR: floating wire w1953
// ERROR: floating wire w1978
// ERROR: floating wire w2003
// ERROR: floating wire w2017
// ERROR: floating wire w2137
// ERROR: floating wire w2573
// ERROR: floating wire w2578
// ERROR: floating wire w2580
// ERROR: floating wire w2622
// ERROR: floating wire w2635
// ERROR: floating wire w2683
// ERROR: floating wire w2917
// ERROR: floating wire w2947
// ERROR: floating wire w3007
// ERROR: floating wire w3019
// ERROR: floating wire w3054
// ERROR: floating wire w3089
// ERROR: floating wire w3163
// ERROR: floating wire w3173
// ERROR: floating wire w3692
// ERROR: floating wire w3834
// ERROR: floating wire w3835
// ERROR: floating wire w3836
// ERROR: floating wire w3860
// ERROR: floating wire w3861
// ERROR: floating wire w3863
// ERROR: floating wire w3864
// ERROR: floating wire w3866
// ERROR: floating wire w3867
// ERROR: floating wire w3869
// ERROR: floating wire w3870
// ERROR: floating wire w3872
// ERROR: floating wire w3873
// ERROR: floating wire w3875
// ERROR: floating wire w3876
// ERROR: floating wire w3878
// ERROR: floating wire w3879
// ERROR: floating wire w3881
// ERROR: floating wire w3924
// ERROR: floating wire w3968
// ERROR: floating wire w3996
// ERROR: floating wire w4001
// ERROR: floating wire w4005
// ERROR: floating wire w4014
// ERROR: floating wire w4070
// ERROR: floating wire w4325
// ERROR: floating wire w4396
// WARNING: Cell ym3438_AND5:g_45 port Z not connected.
// WARNING: Cell ym3438_AND5:g_46 port Z not connected.
// WARNING: Cell ym3438_AND5:g_91 port Z not connected.
// WARNING: Cell ym3438_AND5:g_92 port Z not connected.
// WARNING: Cell ym3438_AND5:g_93 port Z not connected.
// WARNING: Cell ym3438_AND5:g_94 port Z not connected.
// WARNING: Cell ym3438_AND5:g_95 port Z not connected.
// WARNING: Cell ym3438_AND5:g_96 port Z not connected.
// WARNING: Cell ym3438_COMP_STR:g_124 port nZ not connected.
// WARNING: Cell ym3438_FA:g_315 port CO not connected.
// WARNING: Cell ym3438_CNT_BIT:g_561 port CO not connected.
// WARNING: Cell ym3438_CNT_BIT:g_567 port CO not connected.
// WARNING: Cell ym3438_FA:g_888 port S not connected.
// WARNING: Cell ym3438_HA:g_998 port CO not connected.
// WARNING: Cell ym3438_FA:g_1076 port CO not connected.
// WARNING: Cell ym3438_HA:g_1163 port CO not connected.
// WARNING: Cell ym3438_FA:g_1313 port CO not connected.
// WARNING: Cell ym3438_FA:g_1467 port CO not connected.
// WARNING: Cell ym3438_AND:g_1598 port Z not connected.
// WARNING: Cell ym3438_FA:g_1745 port CO not connected.
// WARNING: Cell ym3438_SYNC_SRFF:g_1972 port nQ not connected.
// WARNING: Cell ym3438_SYNC_SRFF:g_1973 port nQ not connected.
// WARNING: Cell ym3438_FA:g_2316 port CO not connected.
// WARNING: Cell ym3438_FA:g_2368 port CO not connected.
// WARNING: Cell ym3438_AON222222:g_2451 port B2 not connected.
// WARNING: Cell ym3438_SR_BIT:g_2795 port D not connected.
// WARNING: Cell ym3438_FA:g_3454 port CO not connected.
// WARNING: Cell ym3438_FA:g_3457 port CO not connected.
// WARNING: Cell ym3438_FA_SEQ:g_3463 port CO not connected.
// WARNING: Cell ym3438_AND3:g_3485 port Z not connected.
// WARNING: Cell ym3438_AND3:g_3486 port Z not connected.
// WARNING: Cell ym3438_COMP_WE:g_3496 port nZ not connected.
// WARNING: Cell ym3438_AND3:g_3629 port Z not connected.
// WARNING: Cell ym3438_FA:g_3690 port CO not connected.
// WARNING: Cell ym3438_HA:g_3782 port CO not connected.
// WARNING: Cell ym3438_HA:g_3875 port CO not connected.
