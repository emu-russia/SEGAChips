module ym6045c (  VA8_o, VA8_d, VA8_i, VA9_o, VA9_d, VA9_i, VA10_o, VA10_d, VA10_i, VA11_o, VA11_d, VA11_i, VA12_o, VA12_d, VA12_i, VA13_o, VA13_d, VA13_i, VA14_o, VA14_d, VA14_i, VA15_o, VA15_d, VA15_i, VA16_o, VA16_d, VA16_i, VA17_o, VA17_d, VA17_i, VA18_o, VA18_d, VA18_i, VA19_o, VA19_d, VA19_i, VA20_o, VA20_d, VA20_i, VA21_o, VA21_d, VA21_i, VA22_o, VA22_d, VA22_i, VA23_o, VA23_d, VA23_i, FC0, FC1, n_VPA, n_RESET, n_HALT, D8_o, D8_d, D8_i, VCLK, n_TIME, n_CAS0, n_DTACK_o, n_DTACK_d, n_DTACK_i, RW_i, RW_d, RW_o, n_LDS_o, n_LDS_d, n_LDS_i, n_UDS_i, n_UDS_d, n_UDS_o, n_AS_o, n_AS_d, n_AS_i, n_INTAK, n_VDPM, n_BG, n_BGACK_i, n_BGACK_d, n_BGACK_o, n_BR, i_EOE, IA14, n_NOE, EDCK, n_OE0, n_HSYNC, MCLK, TPAL, n_SOUND, ZCLK, n_WRES, n_ZRAM, n_REF, n_M1, n_ZRES, n_ZBR, n_WAIT_o, n_WAIT_d, n_WAIT_i, n_ZBAK, n_ZWR_o, n_ZWR_d, n_ZWR_i, n_ZRD_i, n_ZRD_d, n_ZRD_o, n_IREQ, n_MREQ_i, n_MREQ_d, n_MREQ_o, n_NMI, ZA0_i, ZA0_d, ZA0_o, ZA7, ZA8_i, ZA8_d, ZA8_o, ZA9_o, ZA9_d, ZA9_i, ZA10_i, ZA10_d, ZA10_o, ZA11_o, ZA11_d, ZA11_i, ZA12_o, ZA12_d, ZA12_i, ZA13_i, ZA13_d, ZA13_o, ZA14_o, ZA14_d, ZA14_i, ZA15_i, ZA15_d, ZA15_o, ZD0, n_FDWR, n_FDC, n_ROM, n_ASEL, n_CAS2, n_RAS2, n_CE0, n_VTOZ, n_ZTOV, n_SRES, n_IO, n_M3, n_CART, pin99, pin100);

	output wire VA8_o;
	output wire VA8_d;
	input wire VA8_i;
	output wire VA9_o;
	output wire VA9_d;
	input wire VA9_i;
	output wire VA10_o;
	output wire VA10_d;
	input wire VA10_i;
	output wire VA11_o;
	output wire VA11_d;
	input wire VA11_i;
	output wire VA12_o;
	output wire VA12_d;
	input wire VA12_i;
	output wire VA13_o;
	output wire VA13_d;
	input wire VA13_i;
	output wire VA14_o;
	output wire VA14_d;
	input wire VA14_i;
	output wire VA15_o;
	output wire VA15_d;
	input wire VA15_i;
	output wire VA16_o;
	output wire VA16_d;
	input wire VA16_i;
	output wire VA17_o;
	output wire VA17_d;
	input wire VA17_i;
	output wire VA18_o;
	output wire VA18_d;
	input wire VA18_i;
	output wire VA19_o;
	output wire VA19_d;
	input wire VA19_i;
	output wire VA20_o;
	output wire VA20_d;
	input wire VA20_i;
	output wire VA21_o;
	output wire VA21_d;
	input wire VA21_i;
	output wire VA22_o;
	output wire VA22_d;
	input wire VA22_i;
	output wire VA23_o;
	output wire VA23_d;
	input wire VA23_i;
	input wire FC0;
	input wire FC1;
	output wire n_VPA;
	output wire n_RESET;
	output wire n_HALT;
	output wire D8_o;
	output wire D8_d;
	input wire D8_i;
	input wire VCLK;
	output wire n_TIME;
	input wire n_CAS0;
	output wire n_DTACK_o;
	output wire n_DTACK_d;
	input wire n_DTACK_i;
	input wire RW_i;
	output wire RW_d;
	output wire RW_o;
	output wire n_LDS_o;
	output wire n_LDS_d;
	input wire n_LDS_i;
	input wire n_UDS_i;
	output wire n_UDS_d;
	output wire n_UDS_o;
	output wire n_AS_o;
	output wire n_AS_d;
	input wire n_AS_i;
	output wire n_INTAK;
	output wire n_VDPM;
	input wire n_BG;
	input wire n_BGACK_i;
	output wire n_BGACK_d;
	output wire n_BGACK_o;
	output wire n_BR;
	output wire i_EOE;
	output wire IA14;
	output wire n_NOE;
	output wire EDCK;
	input wire n_OE0;
	input wire n_HSYNC;
	input wire MCLK;
	input wire TPAL;
	output wire n_SOUND;
	input wire ZCLK;
	input wire n_WRES;
	output wire n_ZRAM;
	output wire n_REF;
	input wire n_M1;
	output wire n_ZRES;
	output wire n_ZBR;
	output wire n_WAIT_o;
	output wire n_WAIT_d;
	input wire n_WAIT_i;
	input wire n_ZBAK;
	output wire n_ZWR_o;
	output wire n_ZWR_d;
	input wire n_ZWR_i;
	input wire n_ZRD_i;
	output wire n_ZRD_d;
	output wire n_ZRD_o;
	input wire n_IREQ;
	input wire n_MREQ_i;
	output wire n_MREQ_d;
	output wire n_MREQ_o;
	output wire n_NMI;
	input wire ZA0_i;
	output wire ZA0_d;
	output wire ZA0_o;
	input wire ZA7;
	input wire ZA8_i;
	output wire ZA8_d;
	output wire ZA8_o;
	output wire ZA9_o;
	output wire ZA9_d;
	input wire ZA9_i;
	input wire ZA10_i;
	output wire ZA10_d;
	output wire ZA10_o;
	output wire ZA11_o;
	output wire ZA11_d;
	input wire ZA11_i;
	output wire ZA12_o;
	output wire ZA12_d;
	input wire ZA12_i;
	input wire ZA13_i;
	output wire ZA13_d;
	output wire ZA13_o;
	output wire ZA14_o;
	output wire ZA14_d;
	input wire ZA14_i;
	input wire ZA15_i;
	output wire ZA15_d;
	output wire ZA15_o;
	input wire ZD0;
	output wire n_FDWR;
	output wire n_FDC;
	output wire n_ROM;
	output wire n_ASEL;
	output wire n_CAS2;
	output wire n_RAS2;
	output wire n_CE0;
	output wire n_VTOZ;
	output wire n_ZTOV;
	input wire n_SRES;
	output wire n_IO;
	input wire n_M3;
	input wire n_CART;
	output wire pin99;
	output wire pin100;

	// Wires

	wire w1;
	wire w2;
	wire w3;
	wire w4;
	wire w5;
	wire w6;
	wire w7;
	wire w8;
	wire w9;
	wire w10;
	wire w11;
	wire w12;
	wire w13;
	wire w14;
	wire w15;
	wire w16;
	wire w17;
	wire w18;
	wire w19;
	wire w20;
	wire w21;
	wire w22;
	wire w23;
	wire w24;
	wire w25;
	wire w26;
	wire w27;
	wire w28;
	wire w29;
	wire w30;
	wire w31;
	wire w32;
	wire w33;
	wire w34;
	wire w35;
	wire w36;
	wire w37;
	wire w38;
	wire w39;
	wire w40;
	wire w41;
	wire w42;
	wire w43;
	wire w44;
	wire w45;
	wire w46;
	wire w47;
	wire w48;
	wire w49;
	wire w50;
	wire w51;
	wire w52;
	wire w53;
	wire w54;
	wire w55;
	wire w56;
	wire w57;
	wire w58;
	wire w59;
	wire w60;
	wire w61;
	wire w62;
	wire w63;
	wire w64;
	wire w65;
	wire w66;
	wire w67;
	wire w68;
	wire w69;
	wire w70;
	wire w71;
	wire w72;
	wire w73;
	wire w74;
	wire w75;
	wire w76;
	wire w77;
	wire w78;
	wire w79;
	wire w80;
	wire w81;
	wire w82;
	wire w83;
	wire w84;
	wire w85;
	wire w86;
	wire w87;
	wire w88;
	wire w89;
	wire w90;
	wire w91;
	wire w92;
	wire w93;
	wire w94;
	wire w95;
	wire w96;
	wire w97;
	wire w98;
	wire w99;
	wire w100;
	wire w101;
	wire w102;
	wire w103;
	wire w104;
	wire w105;
	wire w106;
	wire w107;
	wire w108;
	wire w109;
	wire w110;
	wire w111;
	wire w112;
	wire w113;
	wire w114;
	wire w115;
	wire w116;
	wire w117;
	wire w118;
	wire w119;
	wire w120;
	wire w121;
	wire w122;
	wire w123;
	wire w124;
	wire w125;
	wire w126;
	wire w127;
	wire w128;
	wire w129;
	wire w130;
	wire w131;
	wire w132;
	wire w133;
	wire w134;
	wire w135;
	wire w136;
	wire w137;
	wire w138;
	wire w139;
	wire w140;
	wire w141;
	wire w142;
	wire w143;
	wire w144;
	wire w145;
	wire w146;
	wire w147;
	wire w148;
	wire w149;
	wire w150;
	wire w151;
	wire w152;
	wire w153;
	wire w154;
	wire w155;
	wire w156;
	wire w157;
	wire w158;
	wire w159;
	wire w160;
	wire w161;
	wire w162;
	wire w163;
	wire w164;
	wire w165;
	wire w166;
	wire w167;
	wire w168;
	wire w169;
	wire w170;
	wire w171;
	wire w172;
	wire w173;
	wire w174;
	wire w175;
	wire w176;
	wire w177;
	wire w178;
	wire w179;
	wire w180;
	wire w181;
	wire w182;
	wire w183;
	wire w184;
	wire w185;
	wire w186;
	wire w187;
	wire w188;
	wire w189;
	wire w190;
	wire w191;
	wire w192;
	wire w193;
	wire w194;
	wire w195;
	wire w196;
	wire w197;
	wire w198;
	wire w199;
	wire w200;
	wire w201;
	wire w202;
	wire w203;
	wire w204;
	wire w205;
	wire w206;
	wire w207;
	wire w208;
	wire w209;
	wire w210;
	wire w211;
	wire w212;
	wire w213;
	wire w214;
	wire w215;
	wire w216;
	wire w217;
	wire w218;
	wire w219;
	wire w220;
	wire w221;
	wire w222;
	wire w223;
	wire w224;
	wire w225;
	wire w226;
	wire w227;
	wire w228;
	wire w229;
	wire w230;
	wire w231;
	wire w232;
	wire w233;
	wire w234;
	wire w235;
	wire w236;
	wire w237;
	wire w238;
	wire w239;
	wire w240;
	wire w241;
	wire w242;
	wire w243;
	wire w244;
	wire w245;
	wire w246;
	wire w247;
	wire w248;
	wire w249;
	wire w250;
	wire w251;
	wire w252;
	wire w253;
	wire w254;
	wire w255;
	wire w256;
	wire w257;
	wire w258;
	wire w259;
	wire w260;
	wire w261;
	wire w262;
	wire w263;
	wire w264;
	wire w265;
	wire w266;
	wire w267;
	wire w268;
	wire w269;
	wire w270;
	wire w271;
	wire w272;
	wire w273;
	wire w274;
	wire w275;
	wire w276;
	wire w277;
	wire w278;
	wire w279;
	wire w280;
	wire w281;
	wire w282;
	wire w283;
	wire w284;
	wire w285;
	wire w286;
	wire w287;
	wire w288;
	wire w289;
	wire w290;
	wire w291;
	wire w292;
	wire w293;
	wire w294;
	wire w295;
	wire w296;
	wire w297;
	wire w298;
	wire w299;
	wire w300;
	wire w301;
	wire w302;
	wire w303;
	wire w304;
	wire w305;
	wire w306;
	wire w307;
	wire w308;
	wire w309;
	wire w310;
	wire w311;
	wire w312;
	wire w313;
	wire w314;
	wire w315;
	wire w316;
	wire w317;
	wire w318;
	wire w319;
	wire w320;
	wire w321;
	wire w322;
	wire w323;
	wire w324;
	wire w325;
	wire w326;
	wire w327;
	wire w328;
	wire w329;
	wire w330;
	wire w331;
	wire w332;
	wire w333;
	wire w334;
	wire w335;
	wire w336;
	wire w337;
	wire w338;
	wire w339;
	wire w340;
	wire w341;
	wire w342;
	wire w343;
	wire w344;
	wire w345;
	wire w346;
	wire w347;
	wire w348;
	wire w349;
	wire w350;
	wire w351;
	wire w352;
	wire w353;
	wire w354;
	wire w355;
	wire w356;
	wire w357;
	wire w358;
	wire w359;
	wire w360;
	wire w361;
	wire w362;
	wire w363;
	wire w364;
	wire w365;
	wire w366;
	wire w367;
	wire w368;
	wire w369;
	wire w370;
	wire w371;
	wire w372;
	wire w373;
	wire w374;
	wire w375;
	wire w376;
	wire w377;
	wire w378;
	wire w379;
	wire w380;
	wire w381;
	wire w382;
	wire w383;
	wire w384;
	wire w385;
	wire w386;
	wire w387;
	wire w388;
	wire w389;
	wire w390;
	wire w391;
	wire w392;
	wire w393;
	wire w394;
	wire w395;
	wire w396;
	wire w397;
	wire w398;
	wire w399;
	wire w400;
	wire w401;
	wire w402;
	wire w403;
	wire w404;
	wire w405;
	wire w406;
	wire w407;
	wire w408;
	wire w409;
	wire w410;
	wire w411;
	wire w412;
	wire w413;
	wire w414;
	wire w415;
	wire w416;
	wire w417;
	wire w418;
	wire w419;
	wire w420;
	wire w421;
	wire w422;
	wire w423;
	wire w424;
	wire w425;
	wire w426;
	wire w427;
	wire w428;
	wire w429;
	wire w430;
	wire w431;
	wire w432;
	wire w433;
	wire w434;
	wire w435;
	wire w436;
	wire w437;
	wire w438;
	wire w439;
	wire w440;
	wire w441;
	wire w442;
	wire w443;
	wire w444;
	wire w445;
	wire w446;
	wire w447;
	wire w448;
	wire w449;
	wire w450;
	wire w451;
	wire w452;
	wire w453;
	wire w454;
	wire w455;
	wire w456;
	wire w457;
	wire w458;
	wire w459;
	wire w460;
	wire w461;
	wire w462;
	wire w463;
	wire w464;
	wire w465;
	wire w466;

	assign VA8_o = w438;
	assign VA8_d = w455;
	assign w81 = VA8_i;
	assign VA9_o = w439;
	assign VA9_d = w455;
	assign w73 = VA9_i;
	assign VA10_o = w461;
	assign VA10_d = w455;
	assign w142 = VA10_i;
	assign VA11_o = w440;
	assign VA11_d = w455;
	assign w56 = VA11_i;
	assign VA12_o = w441;
	assign VA12_d = w455;
	assign w287 = VA12_i;
	assign VA13_o = w442;
	assign VA13_d = w455;
	assign w304 = VA13_i;
	assign VA14_o = w456;
	assign VA14_d = w455;
	assign w92 = VA14_i;
	assign VA15_o = w443;
	assign VA15_d = w455;
	assign w353 = VA15_i;
	assign VA16_o = w444;
	assign VA16_d = w455;
	assign w265 = VA16_i;
	assign VA17_o = w457;
	assign VA17_d = w455;
	assign w358 = VA17_i;
	assign VA18_o = w445;
	assign VA18_d = w455;
	assign w360 = VA18_i;
	assign VA19_o = w446;
	assign VA19_d = w455;
	assign w359 = VA19_i;
	assign VA20_o = w448;
	assign VA20_d = w455;
	assign w369 = VA20_i;
	assign VA21_o = w451;
	assign VA21_d = w449;
	assign w20 = VA21_i;
	assign VA22_o = w383;
	assign VA22_d = w449;
	assign w281 = VA22_i;
	assign VA23_o = w450;
	assign VA23_d = w449;
	assign w463 = VA23_i;
	assign w385 = FC0;
	assign w384 = FC1;
	assign n_VPA = w386;
	assign n_RESET = w465;
	assign n_HALT = w465;
	assign D8_o = w64;
	assign D8_d = w399;
	assign w173 = D8_i;
	assign w171 = VCLK;
	assign n_TIME = w275;
	assign w278 = n_CAS0;
	assign n_DTACK_o = w147;
	assign n_DTACK_d = w143;
	assign w203 = n_DTACK_i;
	assign w50 = RW_i;
	assign RW_d = w197;
	assign RW_o = w57;
	assign n_LDS_o = w100;
	assign n_LDS_d = w437;
	assign w174 = n_LDS_i;
	assign w175 = n_UDS_i;
	assign n_UDS_d = w437;
	assign n_UDS_o = w96;
	assign n_AS_o = w102;
	assign n_AS_d = w437;
	assign w146 = n_AS_i;
	assign n_INTAK = w268;
	assign n_VDPM = w101;
	assign w105 = n_BG;
	assign w200 = n_BGACK_i;
	assign n_BGACK_d = w99;
	assign n_BGACK_o = w95;
	assign n_BR = w97;
	assign i_EOE = w129;
	assign IA14 = w131;
	assign n_NOE = w139;
	assign EDCK = w133;
	assign w452 = n_OE0;
	assign w436 = n_HSYNC;
	assign w433 = MCLK;
	assign w98 = TPAL;
	assign n_SOUND = w89;
	assign w138 = ZCLK;
	assign w60 = n_WRES;
	assign n_ZRAM = w62;
	assign n_REF = w83;
	assign w87 = n_M1;
	assign n_ZRES = w82;
	assign n_ZBR = w117;
	assign n_WAIT_o = w61;
	assign n_WAIT_d = w116;
	assign w93 = n_WAIT_i;
	assign w64 = n_ZBAK;
	assign n_ZWR_o = w67;
	assign n_ZWR_d = w63;
	assign w57 = n_ZWR_i;
	assign w109 = n_ZRD_i;
	assign n_ZRD_d = w63;
	assign n_ZRD_o = w115;
	assign w91 = n_IREQ;
	assign w182 = n_MREQ_i;
	assign n_MREQ_d = w63;
	assign n_MREQ_o = w90;
	assign n_NMI = w66;
	assign w103 = ZA0_i;
	assign ZA0_d = w63;
	assign ZA0_o = w65;
	assign w25 = ZA7;
	assign w24 = ZA8_i;
	assign ZA8_d = w63;
	assign ZA8_o = w81;
	assign ZA9_o = w73;
	assign ZA9_d = w63;
	assign w18 = ZA9_i;
	assign w17 = ZA10_i;
	assign ZA10_d = w63;
	assign ZA10_o = w142;
	assign ZA11_o = w56;
	assign ZA11_d = w63;
	assign w37 = ZA11_i;
	assign ZA12_o = w287;
	assign ZA12_d = w63;
	assign w38 = ZA12_i;
	assign w236 = ZA13_i;
	assign ZA13_d = w63;
	assign ZA13_o = w304;
	assign ZA14_o = w92;
	assign ZA14_d = w63;
	assign w239 = ZA14_i;
	assign w32 = ZA15_i;
	assign ZA15_d = w63;
	assign ZA15_o = w453;
	assign w230 = ZD0;
	assign n_FDWR = w454;
	assign n_FDC = w155;
	assign n_ROM = w27;
	assign n_ASEL = w1;
	assign n_CAS2 = w46;
	assign n_RAS2 = w58;
	assign n_CE0 = w19;
	assign n_VTOZ = w63;
	assign n_ZTOV = w269;
	assign w88 = n_SRES;
	assign n_IO = w86;
	assign w35 = n_M3;
	assign w288 = n_CART;
	assign pin99 = w76;
	assign pin100 = w315;

	// Instances

	ym6045c_NOT g_1 (.A(w140), .nZ(w139) );
	ym6045c_AND g_2 (.Z(w127), .B(w120), .A(w122) );
	ym6045c_NAND g_3 (.A(w35), .B(w107), .Z(w129) );
	ym6045c_BUF g_4 (.Z(w134), .A(w130) );
	ym6045c_NAND g_5 (.A(w92), .B(w35), .Z(w131) );
	ym6045c_NAND3 g_6 (.A(w121), .B(w128), .C(w124), .Z(w119) );
	ym6045c_BUF g_7 (.Z(w84), .A(w120) );
	ym6045c_CNT_BIT g_8 (.Q(w122), .nQ(w121), .C(w433), .RES(w94), .D(w132), .nLD(w119), .CI(1'b1) );
	ym6045c_CNT_BIT g_9 (.nQ(w128), .C(w433), .RES(w94), .D(1'b1), .nLD(w119), .CI(w127) );
	ym6045c_NOT g_10 (.A(w84), .nZ(w85) );
	ym6045c_NOT g_11 (.A(w436), .nZ(w135) );
	ym6045c_BUF g_12 (.Z(w94), .A(w88) );
	ym6045c_AND6 g_13 (.Z(w59), .F(w75), .E(w20), .D(w265), .C(1'b1), .B(w92), .A(w190) );
	ym6045c_BUF g_14 (.Z(w108), .A(w84) );
	ym6045c_NOR4 g_15 (.Z(w136), .D(w114), .C(w113), .B(w432), .A(w141) );
	ym6045c_CNT_BIT g_16 (.nQ(w114), .C(w108), .RES(w111), .D(1'b0), .nLD(w104), .CI(w112) );
	ym6045c_CNT_BIT g_17 (.nQ(w113), .C(w108), .RES(w111), .D(1'b0), .nLD(w104), .CO(w112), .CI(w123) );
	ym6045c_CNT_BIT g_18 (.nQ(w141), .C(w108), .RES(w111), .D(1'b0), .nLD(w104), .CO(w123), .CI(w110) );
	ym6045c_CNT_BIT g_19 (.Q(w120), .nQ(w124), .C(w433), .RES(w94), .D(1'b0), .nLD(w119), .CI(w122) );
	ym6045c_DFFSPOS g_20 (.C(w84), .D(w136), .nSET(w111), .nQ(w106) );
	ym6045c_JKFF g_21 (.C(w85), .K(w135), .J(1'b0), .nSET(w134), .nQ(w104), .Q(w132) );
	ym6045c_BUF g_22 (.A(w84), .Z(w133) );
	ym6045c_AND g_25 (.Z(w1), .B(w2), .A(w3) );
	ym6045c_DELAY g_26 (.Z(w2), .A(w10) );
	ym6045c_AND4 g_27 (.Z(w19), .D(w4), .C(w13), .B(w6), .A(w77) );
	ym6045c_OR g_28 (.A(w7), .Z(w6), .B(w12) );
	ym6045c_NOR g_29 (.Z(w11), .B(w8), .A(w12) );
	ym6045c_OR3 g_30 (.Z(w4), .C(w11), .B(w14), .A(w16) );
	ym6045c_NOT g_31 (.A(w14), .nZ(w5) );
	ym6045c_NAND4 g_32 (.B(w5), .C(w8), .A(w20), .D(w16), .Z(w15) );
	ym6045c_AND3 g_33 (.Z(w58), .C(w15), .B(w7), .A(w9) );
	ym6045c_DELAY_S g_34 (.Z(w10), .A(w34) );
	ym6045c_OR3 g_35 (.Z(w13), .C(w35), .B(w32), .A(w33) );
	ym6045c_NOT g_36 (.A(w24), .nZ(w28) );
	ym6045c_NOT g_37 (.A(w17), .nZ(w30) );
	ym6045c_NAND6 g_38 (.C(w23), .D(w28), .B(w22), .E(w30), .A(1'b1), .F(w29), .Z(w36) );
	ym6045c_NOT g_39 (.A(w38), .nZ(w22) );
	ym6045c_NOT g_40 (.A(w37), .nZ(w29) );
	ym6045c_NAND6 g_41 (.A(w24), .F(w17), .B(w18), .E(w37), .C(1'b1), .D(w38), .Z(w31) );
	ym6045c_NOT g_42 (.A(w18), .nZ(w23) );
	ym6045c_AND g_43 (.Z(w27), .B(w40), .A(w235) );
	ym6045c_AND3 g_44 (.Z(w46), .C(w49), .B(w267), .A(w462) );
	ym6045c_OR4 g_45 (.Z(w49), .D(w239), .C(w33), .B(w55), .A(w35) );
	ym6045c_DFFPOS g_46 (.nQ(w454), .Q(w48), .D(w47), .C(w171) );
	ym6045c_NOR3 g_47 (.Z(w47), .C(w48), .B(w155), .A(w50) );
	ym6045c_NOT g_48 (.A(w32), .nZ(w55) );
	ym6045c_OR g_49 (.B(w54), .Z(w53), .A(w31) );
	ym6045c_AND g_50 (.Z(w52), .B(w51), .A(w53) );
	ym6045c_NAND4 g_51 (.B(w35), .D(w239), .A(w236), .C(w55), .Z(w54) );
	ym6045c_OR4 g_52 (.Z(w224), .A(w57), .B(w33), .C(w54), .D(w36) );
	ym6045c_DFFRPOS g_53 (.Q(w51), .nRES(w253), .D(w225), .C(w224) );
	ym6045c_DELAY g_54 (.Z(w41), .A(w231) );
	ym6045c_DFFSPOS g_55 (.C(w223), .D(w75), .nSET(w222), .Q(w66) );
	ym6045c_OR g_56 (.B(w50), .Z(w67), .A(w146) );
	ym6045c_AND g_57 (.Z(w65), .B(w175), .A(w221) );
	ym6045c_DFFPOS g_58 (.Q(w221), .D(w175), .C(w176) );
	ym6045c_NOT g_59 (.A(w236), .nZ(w68) );
	ym6045c_NOT g_60 (.A(w33), .nZ(w70) );
	ym6045c_NAND g_61 (.A(w59), .B(w233), .Z(w234) );
	ym6045c_NAND6 g_62 (.C(w68), .D(w55), .B(w70), .E(w239), .A(1'b1), .F(w35), .Z(w89) );
	ym6045c_NAND4 g_63 (.B(w70), .C(w35), .A(w71), .D(w55), .Z(w62) );
	ym6045c_NOT g_64 (.A(w239), .nZ(w71) );
	ym6045c_OR g_65 (.A(w64), .Z(w63), .B(w266) );
	ym6045c_DFFRPOS g_66 (.nQ(w261), .Q(w245), .nRES(w244), .D(w60), .C(w223) );
	ym6045c_DFFRPOS g_67 (.Q(w249), .nRES(w244), .D(w245), .C(w247) );
	ym6045c_NOR g_68 (.Z(w246), .B(w249), .A(w261) );
	ym6045c_AND g_69 (.Z(w86), .B(w157), .A(w264) );
	ym6045c_OR3 g_70 (.Z(w252), .C(w250), .B(w35), .A(w91) );
	ym6045c_AND g_71 (.Z(w264), .B(w252), .A(w251) );
	ym6045c_DFFPOS g_72 (.Q(w251), .D(w252), .C(w138) );
	ym6045c_NOR g_73 (.Z(w256), .B(w175), .A(w50) );
	ym6045c_NOT g_74 (.A(w87), .nZ(w250) );
	ym6045c_DFFPOS g_75 (.nQ(w283), .Q(w253), .D(w88), .C(w171) );
	ym6045c_OR g_76 (.A(w146), .Z(w115), .B(w168) );
	ym6045c_NOR g_77 (.Z(w166), .B(w167), .A(w146) );
	ym6045c_DFFRPOS g_78 (.nQ(w117), .nRES(w253), .D(w173), .C(w169) );
	ym6045c_OR g_79 (.B(w50), .Z(w169), .A(w162) );
	ym6045c_NAND3 g_80 (.A(w170), .B(w151), .C(w172), .Z(w90) );
	ym6045c_DFFPOS g_81 (.Q(w172), .D(w151), .C(w171) );
	ym6045c_OR g_82 (.A(w117), .Z(w153), .B(w64) );
	ym6045c_NAND g_83 (.A(w82), .B(w153), .Z(w150) );
	ym6045c_NOT g_84 (.Z(w176), .A(w171) );
	ym6045c_NOR g_85 (.Z(w83), .B(w204), .A(w206) );
	ym6045c_NOT g_86 (.A(w50), .nZ(w168) );
	ym6045c_NAND g_87 (.A(w174), .B(w175), .Z(w151) );
	ym6045c_AND g_88 (.Z(w177), .B(w154), .A(w452) );
	ym6045c_BUF g_89 (.Z(w208), .A(w94) );
	ym6045c_NOT g_90 (.A(w88), .nZ(w209) );
	ym6045c_OR3 g_91 (.Z(w212), .C(w186), .B(w178), .A(w209) );
	ym6045c_NOT g_92 (.A(w179), .nZ(w178) );
	ym6045c_DFFPOS g_93 (.Q(w189), .D(w179), .C(w171) );
	ym6045c_OR3 g_94 (.Z(w116), .C(w213), .B(w186), .A(w187) );
	ym6045c_OR g_95 (.B(w186), .Z(w180), .A(w189) );
	ym6045c_NOT g_96 (.A(w146), .nZ(w190) );
	ym6045c_BUF g_97 (.Z(w111), .A(w88) );
	ym6045c_CNT_BIT g_98 (.nQ(w432), .C(w108), .RES(w111), .D(1'b1), .nLD(w104), .CO(w110), .CI(w104) );
	ym6045c_NOT g_99 (.A(w146), .nZ(w183) );
	ym6045c_OR4 g_100 (.Z(w184), .D(w183), .C(w186), .B(w181), .A(w105) );
	ym6045c_DFFPOS g_101 (.Q(w194), .D(w180), .C(w171) );
	ym6045c_OR g_102 (.A(w194), .Z(w102), .B(w186) );
	ym6045c_NOT g_103 (.A(w139), .nZ(w107) );
	ym6045c_DFFPOS g_104 (.Q(w466), .D(w102), .C(w171) );
	ym6045c_OR g_105 (.B(w57), .Z(w214), .A(w466) );
	ym6045c_OR g_106 (.A(w102), .B(w109), .Z(w198) );
	ym6045c_AND g_107 (.Z(w191), .B(w214), .A(w198) );
	ym6045c_OR g_108 (.B(w193), .Z(w101), .A(w173) );
	ym6045c_NOT g_109 (.A(w103), .nZ(w192) );
	ym6045c_OR g_110 (.B(w191), .Z(w96), .A(w103) );
	ym6045c_OR g_111 (.B(w191), .Z(w100), .A(w192) );
	ym6045c_BUF g_112 (.Z(w130), .A(w106) );
	ym6045c_DFFPOS g_113 (.Q(w97), .D(w212), .C(w171) );
	ym6045c_NOT g_114 (.A(w98), .nZ(w213) );
	ym6045c_OR g_115 (.B(w197), .Z(w99), .A(w213) );
	ym6045c_MUX4BIT g_118 (.C(w35), .Z0(w241), .B1(w17), .A1(w37), .B2(w18), .A2(w17), .Z1(w243), .Z2(w242), .A3(w18), .B3(w24), .B4(w25), .A4(w24), .Z3(w240) );
	ym6045c_NOT g_119 (.A(w42), .nZ(w16) );
	ym6045c_XNOR g_120 (.A(w288), .B(w281), .Z(w42) );
	ym6045c_NOT g_121 (.A(w20), .nZ(w434) );
	ym6045c_OR3 g_122 (.Z(w39), .C(w34), .B(w42), .A(w434) );
	ym6045c_AND g_123 (.B(w39), .A(w41), .Z(w9) );
	ym6045c_OR3 g_124 (.Z(w40), .C(w42), .B(w14), .A(w20) );
	ym6045c_MUX4BIT g_125 (.C(w35), .Z0(w238), .B1(w239), .A1(w52), .B2(w236), .A2(w239), .Z1(w237), .Z2(w328), .A3(w236), .B3(w38), .B4(w37), .A4(w38), .Z3(w291) );
	ym6045c_NOT g_126 (.nZ(w43), .A(w42) );
	ym6045c_OR3 g_127 (.Z(w235), .C(w74), .B(w20), .A(w42) );
	ym6045c_AND g_128 (.Z(w77), .B(w44), .A(w79) );
	ym6045c_AND g_129 (.Z(w462), .B(w292), .A(w295) );
	ym6045c_OR g_130 (.A(w45), .Z(w44), .B(w43) );
	ym6045c_MUX g_131 (.C(w12), .Z(w45), .A(w34), .B(w74) );
	ym6045c_OR g_132 (.B(w41), .Z(w79), .A(w12) );
	ym6045c_OR g_133 (.A(w289), .Z(w34), .B(w75) );
	ym6045c_OR g_134 (.A(w14), .Z(w158), .B(w290) );
	ym6045c_OR3 g_135 (.Z(w14), .C(w75), .B(w78), .A(w146) );
	ym6045c_NOT g_136 (.A(w35), .nZ(w78) );
	ym6045c_NOR g_137 (.Z(w222), .B(w226), .A(w80) );
	ym6045c_NOR g_138 (.Z(w80), .B(w226), .A(w244) );
	ym6045c_OR8 g_139 (.A(1'b0), .E(w56), .B(w234), .F(w142), .Z(w76), .C(w174), .G(w73), .D(w175), .H(w81) );
	ym6045c_SIPO_8BIT g_140 (.nRES(w253), .Q0(w225), .Q1(w303), .Q2(w227), .Q3(w300), .Q4(w228), .Q5(w229), .Q6(w286), .Q7(w285), .D(w230), .C(w224) );
	ym6045c_OR g_141 (.A(w284), .Z(w231), .B(w232) );
	ym6045c_DELAY g_142 (.Z(w232), .A(w267) );
	ym6045c_NOR g_143 (.Z(w302), .B(w246), .A(w301) );
	ym6045c_DEC_2TO4 g_144 (.A1(w304), .Z3(w248), .Z2(w259), .A0(w287), .Z0(w263), .Z1(w262) );
	ym6045c_NAND3 g_145 (.A(w262), .B(w305), .C(w265), .Z(w156) );
	ym6045c_NAND4 g_146 (.B(w259), .C(w305), .A(w255), .D(w265), .Z(w260) );
	ym6045c_NAND4 g_147 (.B(w248), .C(w305), .A(w255), .D(w265), .Z(w163) );
	ym6045c_NAND4 g_148 (.B(w263), .C(w305), .A(w255), .D(w265), .Z(w157) );
	ym6045c_OR g_149 (.B(w146), .Z(w155), .A(w260) );
	ym6045c_NOT g_150 (.A(w35), .nZ(w258) );
	ym6045c_OR3 g_151 (.Z(w218), .C(w33), .B(w258), .A(w55) );
	ym6045c_NAND3 g_153 (.A(w220), .B(w256), .C(w257), .Z(w282) );
	ym6045c_NAND3 g_154 (.A(w255), .B(w220), .C(w256), .Z(w254) );
	ym6045c_DFFRPOS g_155 (.nQ(w12), .nRES(w253), .D(w173), .C(w254) );
	ym6045c_OR g_156 (.A(w33), .Z(w219), .i4(w53) );
	ym6045c_AND g_157 (.Z(w199), .B(w219), .A(w218) );
	ym6045c_NOR g_158 (.Z(w160), .B(w165), .A(w166) );
	ym6045c_NOT g_159 (.A(w156), .nZ(w220) );
	ym6045c_NAND3 g_160 (.A(w220), .B(w164), .C(w161), .Z(w162) );
	ym6045c_NOT g_161 (.A(w175), .nZ(w161) );
	ym6045c_DFFSPOS g_162 (.C(w176), .D(w160), .nSET(w150), .nQ(w159), .Q(w167) );
	ym6045c_OR g_163 (.B(w146), .Z(w152), .A(w266) );
	ym6045c_OR g_164 (.B(w146), .Z(w277), .A(w156) );
	ym6045c_NAND6 g_165 (.C(w157), .D(w276), .B(w155), .E(w275), .A(w158), .F(w277), .Z(w148) );
	ym6045c_OR g_166 (.A(w163), .Z(w275), .B(w146) );
	ym6045c_OR g_167 (.B(w205), .Z(w276), .A(w152) );
	ym6045c_NAND g_168 (.A(w201), .B(w93), .Z(w205) );
	ym6045c_OR g_169 (.B(w177), .Z(w211), .A(w274) );
	ym6045c_OAI21 g_170 (.Z(w140), .A2(w280), .B(w211), .A1(w279) );
	ym6045c_OR4 g_171 (.Z(w193), .D(w35), .C(w182), .B(w173), .A(w281) );
	ym6045c_NOR3 g_172 (.Z(w204), .C(w272), .B(w207), .A(w182) );
	ym6045c_NOR g_173 (.Z(w206), .B(w207), .A(w273) );
	ym6045c_NOT g_174 (.A(w35), .nZ(w207) );
	ym6045c_AND g_175 (.Z(w269), .B(w35), .A(w210) );
	ym6045c_OR g_176 (.A(w209), .Z(w210), .B(w188) );
	ym6045c_OR3 g_177 (.Z(w179), .C(w186), .B(w188), .A(w209) );
	ym6045c_NAND g_178 (.A(w159), .B(w146), .Z(w217) );
	ym6045c_NOR g_179 (.Z(w187), .B(w179), .A(w203) );
	ym6045c_DFFPOS g_180 (.Q(w202), .D(w87), .C(w138) );
	ym6045c_DFFPOS g_181 (.Q(w216), .D(w202), .C(w138) );
	ym6045c_AND g_182 (.Z(w196), .B(w179), .A(w184) );
	ym6045c_DFFPOS g_183 (.D(w196), .C(w176), .Q(w188) );
	ym6045c_DFFPOS g_184 (.nQ(w170), .Q(w149), .D(w271), .C(w176) );
	ym6045c_NOT g_185 (.A(w200), .nZ(w181) );
	ym6045c_DFFPOS g_186 (.Q(w195), .D(w199), .C(w138) );
	ym6045c_AND g_187 (.Z(w186), .B(w195), .A(w199) );
	ym6045c_BUF g_188 (.Z(w197), .A(w210) );
	ym6045c_AND g_189 (.Z(w270), .B(w269), .A(w215) );
	ym6045c_OR g_190 (.B(w200), .Z(w215), .A(w270) );
	ym6045c_DFFPOS g_191 (.nQ(w201), .D(w145), .C(w171) );
	ym6045c_OR3 g_192 (.Z(w145), .C(w144), .B(w146), .A(w149) );
	ym6045c_DFFPOS g_193 (.Q(w144), .D(w146), .C(w171) );
	ym6045c_NAND g_194 (.A(w148), .B(w268), .Z(w143) );
	ym6045c_NOR4 g_195 (.Z(w330), .D(w307), .C(w316), .B(w314), .A(w319) );
	ym6045c_NAND g_196 (.A(w320), .B(w321), .Z(w308) );
	ym6045c_AND g_197 (.Z(w309), .B(w308), .A(w327) );
	ym6045c_DFFSPOS g_198 (.C(w171), .D(w309), .nSET(w298), .nQ(w320), .Q(w322) );
	ym6045c_DFFPOS g_199 (.Q(w324), .D(w3), .C(w176) );
	ym6045c_DFFPOS g_200 (.nQ(w299), .Q(w321), .D(w323), .C(w176) );
	ym6045c_OR g_201 (.B(w292), .Z(w323), .A(w322) );
	ym6045c_NOR g_202 (.Z(w8), .A(w325), .B(w299) );
	ym6045c_OR g_203 (.A(w324), .Z(w292), .B(w325) );
	ym6045c_DFFPOS g_204 (.Q(w326), .D(w325), .C(w171) );
	ym6045c_OR g_205 (.B(w325), .Z(w3), .A(w326) );
	ym6045c_OR g_206 (.B(w320), .Z(w290), .A(w3) );
	ym6045c_OR g_207 (.B(w335), .Z(w327), .A(w75) );
	ym6045c_NOT g_208 (.A(w20), .nZ(w293) );
	ym6045c_NAND4 g_209 (.B(w190), .C(w75), .A(w281), .D(w293), .Z(w315) );
	ym6045c_DFFRPOS g_210 (.nQ(w294), .nRES(w298), .D(w299), .C(w176) );
	ym6045c_NOR g_211 (.Z(w7), .B(w294), .A(w350) );
	ym6045c_OR g_212 (.A(w349), .Z(w74), .B(w289) );
	ym6045c_OR3 g_213 (.Z(w325), .C(w296), .B(w75), .A(w351) );
	ym6045c_NAND g_214 (.A(w297), .B(w295), .Z(w296) );
	ym6045c_DFFSPOS g_215 (.C(w176), .D(w295), .nSET(w298), .Q(w297) );
	ym6045c_OR4 g_216 (.Z(w354), .D(w353), .C(w92), .B(w142), .A(w56) );
	ym6045c_DFFSPOS g_217 (.C(w176), .D(w348), .nSET(w298), .nQ(w350), .Q(w352) );
	ym6045c_AND g_218 (.Z(w295), .A(w348), .B(w352) );
	ym6045c_AND g_219 (.Z(w298), .A(w35), .B(w253) );
	ym6045c_AND g_220 (.Z(w342), .A(w225), .B(w53) );
	ym6045c_AND g_221 (.Z(w356), .A(w53), .B(w300) );
	ym6045c_AND g_222 (.Z(w343), .A(w227), .B(w53) );
	ym6045c_AND g_223 (.Z(w357), .A(w303), .B(w53) );
	ym6045c_NOR8 g_224 (.A(w353), .B(w287), .C(w304), .D(w358), .Z(w233), .E(w360), .F(w359), .G(w369), .H(w281) );
	ym6045c_OR4 g_225 (.Z(w370), .D(w359), .C(w369), .B(w358), .A(w360) );
	ym6045c_NOT g_226 (.A(w53), .nZ(w347) );
	ym6045c_DFFRPOS g_227 (.nQ(w301), .nRES(w244), .D(w368), .C(w223) );
	ym6045c_DFFRPOS g_228 (.Q(w368), .nRES(w244), .D(w244), .C(w223) );
	ym6045c_NOR3 g_229 (.Z(w305), .C(w354), .B(w370), .A(w361) );
	ym6045c_OR3 g_230 (.Z(w266), .C(w265), .B(w361), .A(w370) );
	ym6045c_TFF g_231 (.nQ(w223), .C(w371), .T(w244) );
	ym6045c_BUF g_232 (.Z(w244), .A(w253) );
	ym6045c_NOT g_233 (.A(w332), .nZ(w247) );
	ym6045c_AND g_234 (.Z(w373), .A(w53), .B(w285) );
	ym6045c_AND g_235 (.Z(w372), .A(w53), .B(w286) );
	ym6045c_AND g_236 (.Z(w374), .A(w53), .B(w229) );
	ym6045c_AND g_237 (.Z(w376), .A(w53), .B(w228) );
	ym6045c_BUF g_238 (.Z(w317), .A(w458) );
	ym6045c_NOR g_239 (.Z(w458), .B(w355), .A(w283) );
	ym6045c_NOR g_240 (.Z(w459), .B(w365), .A(w355) );
	ym6045c_NOR g_241 (.Z(w165), .B(w283), .A(w459) );
	ym6045c_DFFSPOS g_242 (.C(w338), .D(w378), .nSET(w375), .nQ(w378), .Q(w284) );
	ym6045c_NOT g_243 (.A(w278), .nZ(w338) );
	ym6045c_OR g_244 (.B(w289), .Z(w267), .A(w278) );
	ym6045c_BUF g_245 (.Z(w460), .A(w210) );
	ym6045c_NOT g_246 (.A(w427), .nZ(w379) );
	ym6045c_DFFRPOS g_247 (.Q(w380), .nRES(w379), .D(w93), .C(w381) );
	ym6045c_AND g_248 (.Z(w274), .B(w278), .A(w382) );
	ym6045c_DFFRPOS g_249 (.nQ(w154), .Q(w426), .nRES(w380), .D(w419), .C(w400) );
	ym6045c_DFFRPOS g_250 (.nQ(w424), .Q(w280), .nRES(w208), .D(w382), .C(w400) );
	ym6045c_OAI21 g_251 (.Z(w427), .A1(w424), .B(w208), .A2(w382) );
	ym6045c_DFFRPOS g_252 (.nQ(w279), .Q(w419), .nRES(w380), .D(w381), .C(w171) );
	ym6045c_OR g_253 (.B(w162), .Z(w399), .A(w168) );
	ym6045c_NOT g_254 (.A(w171), .nZ(w400) );
	ym6045c_NOT g_255 (.A(w200), .nZ(w381) );
	ym6045c_NOT g_256 (.A(w35), .nZ(w393) );
	ym6045c_OR3 g_257 (.Z(w289), .C(w395), .B(w200), .A(w393) );
	ym6045c_NOT g_258 (.A(w270), .nZ(w395) );
	ym6045c_NOT g_259 (.A(w138), .nZ(w398) );
	ym6045c_DFFPOS g_260 (.nQ(w401), .Q(w272), .D(w216), .C(w398) );
	ym6045c_DFFPOS g_261 (.nQ(w397), .D(w396), .C(w176) );
	ym6045c_NAND g_262 (.A(w217), .B(w273), .Z(w396) );
	ym6045c_NAND3 g_263 (.A(w397), .B(w273), .C(w217), .Z(w271) );
	ym6045c_DFFPOS g_264 (.Q(w273), .D(w217), .C(w176) );
	ym6045c_MUX g_265 (.C(w35), .Z(w82), .A(w302), .B(w407) );
	ym6045c_DFFRPOS g_266 (.Q(w407), .nRES(w302), .D(w173), .C(w282) );
	ym6045c_TFF g_267 (.Q(w405), .C(w394), .T(w402) );
	ym6045c_TFF g_268 (.Q(w417), .C(w405), .T(w402) );
	ym6045c_DELAY g_269 (.Z(w403), .A(w289) );
	ym6045c_NAND g_270 (.A(w289), .B(w403), .Z(w404) );
	ym6045c_AND g_273 (.Z(w440), .B(w306), .A(w241) );
	ym6045c_AND g_274 (.Z(w438), .B(w306), .A(w240) );
	ym6045c_AND g_275 (.Z(w439), .B(w306), .A(w242) );
	ym6045c_AND g_276 (.Z(w461), .B(w306), .A(w243) );
	ym6045c_CNT_BIT g_277 (.nQ(w307), .C(w171), .RES(1'b1), .D(1'b0), .nLD(w317), .CO(w311), .CI(w312) );
	ym6045c_CNT_BIT g_278 (.nQ(w319), .C(w171), .RES(1'b1), .D(1'b0), .nLD(w317), .CO(w329), .CI(w311) );
	ym6045c_CNT_BIT g_279 (.nQ(w314), .C(w171), .RES(1'b1), .D(1'b0), .nLD(w317), .CO(w318), .CI(w329) );
	ym6045c_CNT_BIT g_280 (.nQ(w316), .C(w171), .RES(1'b1), .D(w35), .nLD(w317), .CI(w318) );
	ym6045c_AND g_281 (.Z(w441), .B(w306), .A(w291) );
	ym6045c_AND g_282 (.Z(w442), .B(w306), .A(w328) );
	ym6045c_AND g_283 (.Z(w456), .B(w237), .A(w306) );
	ym6045c_AND g_284 (.Z(w443), .B(w238), .A(w306) );
	ym6045c_AND3 g_285 (.Z(w312), .A(w317), .B(w334), .C(w334) );
	ym6045c_NAND g_286 (.A(w333), .B(w75), .Z(w336) );
	ym6045c_AND g_287 (.Z(w337), .B(w336), .A(w435) );
	ym6045c_NAND3 g_288 (.A(w332), .B(w335), .C(w334), .Z(w435) );
	ym6045c_DFFRPOS g_289 (.nQ(w335), .Q(w333), .nRES(w332), .D(w332), .C(w331) );
	ym6045c_NOT g_290 (.A(w351), .nZ(w331) );
	ym6045c_NOT g_291 (.A(w35), .nZ(w464) );
	ym6045c_OR g_292 (.B(w146), .Z(w351), .A(w464) );
	ym6045c_NOT g_293 (.A(w347), .nZ(w306) );
	ym6045c_DFFSPOS g_294 (.C(w171), .D(w337), .nSET(w298), .Q(w348) );
	ym6045c_AND g_295 (.Z(w355), .B(w334), .A(w330) );
	ym6045c_AND3 g_296 (.Z(w349), .C(w75), .B(w341), .A(w338) );
	ym6045c_DFFSPOS g_297 (.C(w338), .D(w75), .nSET(w340), .Q(w341) );
	ym6045c_NOT g_298 (.A(w289), .nZ(w340) );
	ym6045c_OR g_299 (.B(w20), .Z(w339), .A(w182) );
	ym6045c_MUX4BIT g_300 (.C(w35), .Z0(w446), .B1(w91), .A1(w356), .B2(w182), .A2(w343), .Z1(w445), .Z2(w457), .A3(w357), .B3(w339), .B4(w32), .A4(w342), .Z3(w444) );
	ym6045c_NOT g_301 (.A(w289), .nZ(w344) );
	ym6045c_NOR4 g_302 (.Z(w345), .D(w333), .C(w344), .B(w334), .A(w346) );
	ym6045c_DFFSPOS g_303 (.C(w171), .D(w367), .nSET(w253), .nQ(w332), .Q(w346) );
	ym6045c_NOR3 g_304 (.Z(w367), .C(w345), .B(w355), .A(w365) );
	ym6045c_NOT g_305 (.A(w281), .nZ(w447) );
	ym6045c_NAND4 g_306 (.B(w35), .C(w447), .A(w75), .D(w20), .Z(w361) );
	ym6045c_TFF g_307 (.Q(w366), .C(w363), .T(w362) );
	ym6045c_TFF g_308 (.Q(w363), .C(w364), .T(w362) );
	ym6045c_TFF g_309 (.Q(w364), .C(w430), .T(w362) );
	ym6045c_NOR g_310 (.Z(w430), .B(w332), .A(w425) );
	ym6045c_TFF g_311 (.Q(w422), .C(w366), .T(w362) );
	ym6045c_OR g_312 (.B(w347), .Z(w377), .A(w373) );
	ym6045c_OR g_313 (.A(w372), .o3(w429), .B(w347) );
	ym6045c_MUX4BIT g_314 (.C(w35), .Z0(w450), .B1(1'b0), .A1(w377), .B2(1'b0), .A2(w429), .Z1(w383), .Z2(w451), .A3(w374), .B3(1'b0), .B4(w82), .A4(w376), .Z3(w448) );
	ym6045c_NOT g_315 (.A(w283), .nZ(w362) );
	ym6045c_OR g_316 (.A(w213), .Z(w455), .B(w269) );
	ym6045c_OR g_317 (.A(w460), .Z(w449), .B(w213) );
	ym6045c_OR g_318 (.A(w401), .Z(w33), .B(w182) );
	ym6045c_NOR g_319 (.Z(w365), .B(w226), .A(w392) );
	ym6045c_NOT g_320 (.A(w283), .nZ(w402) );
	ym6045c_DFFRPOS g_321 (.Q(w382), .nRES(w380), .D(w426), .C(w171) );
	ym6045c_TFF g_322 (.Q(w371), .C(w417), .T(w402) );
	ym6045c_AND g_323 (.Z(w375), .B(w463), .A(w404) );
	ym6045c_BUF g_324 (.Z(w226), .A(w35) );
	ym6045c_NOR g_325 (.Z(w425), .B(w226), .A(w421) );
	ym6045c_OR g_326 (.A(w423), .Z(w387), .B(w422) );
	ym6045c_NOR g_327 (.Z(w423), .B(w226), .A(w420) );
	ym6045c_NOT g_328 (.A(w391), .nZ(w392) );
	ym6045c_NOT g_329 (.A(w389), .nZ(w420) );
	ym6045c_NOT g_330 (.A(w390), .nZ(w421) );
	ym6045c_DEC_2TO4 g_331 (.A1(w384), .Z3(w388), .Z1(w389), .A0(w385), .Z2(w390), .Z0(w391) );
	ym6045c_NAND g_332 (.A(w388), .B(w269), .Z(w268) );
	ym6045c_OR g_333 (.B(w268), .Z(w386), .A(w146) );
	ym6045c_TFF g_334 (.Q(w394), .C(w387), .T(w402) );
	ym6045c_AND g_335 (.Z(w465), .B(w302), .A(w35) );
	ym6045c_AND g_336 (.Z(w334), .B(1'b1), .A(w418) );
	ym6045c_CNT_BIT g_337 (.nQ(w410), .C(w171), .RES(1'b1), .D(1'b0), .nLD(w317), .CI(w408) );
	ym6045c_CNT_BIT g_338 (.nQ(w413), .C(w171), .RES(1'b1), .D(1'b0), .nLD(w317), .CO(w408), .CI(w409) );
	ym6045c_NOR4 g_339 (.Z(w418), .D(w410), .C(w413), .B(w416), .A(w406) );
	ym6045c_CNT_BIT g_340 (.nQ(w416), .C(w171), .RES(1'b1), .D(1'b0), .nLD(w317), .CO(w409), .CI(w412) );
	ym6045c_CNT_BIT g_341 (.nQ(w406), .C(w171), .RES(1'b1), .D(1'b0), .nLD(w317), .CO(w412), .CI(w415) );
	ym6045c_AND3 g_342 (.Z(w415), .C(w317), .B(1'b1), .A(1'b1) );
	ym6045c_OR g_343 (.A(w213), .Z(w437), .B(w197) );
	ym6045c_DEC_2TO4 g_152 (.A0(w81), .A1(w73), .Z2(w257), .Z0(w255), .Z1(w164) );
endmodule // ym6045c

// Module Definitions [It is possible to wrap here on your primitives]

module ym6045c_NOT (  A, nZ);

	input wire A;
	output wire nZ;

endmodule // ym6045c_NOT

module ym6045c_AND (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // ym6045c_AND

module ym6045c_NAND (  A, B, Z);

	input wire A;
	input wire B;
	output wire Z;

endmodule // ym6045c_NAND

module ym6045c_BUF (  Z, A);

	output wire Z;
	input wire A;

endmodule // ym6045c_BUF

module ym6045c_NAND3 (  A, B, C, Z);

	input wire A;
	input wire B;
	input wire C;
	output wire Z;

endmodule // ym6045c_NAND3

module ym6045c_CNT_BIT (  Q, nQ, C, RES, D, nLD, CO, CI);

	output wire Q;
	output wire nQ;
	input wire C;
	input wire RES;
	input wire D;
	input wire nLD;
	output wire CO;
	input wire CI;

endmodule // ym6045c_CNT_BIT

module ym6045c_AND6 (  Z, F, E, D, C, B, A);

	output wire Z;
	input wire F;
	input wire E;
	input wire D;
	input wire C;
	input wire B;
	input wire A;

endmodule // ym6045c_AND6

module ym6045c_NOR4 (  Z, D, C, B, A);

	output wire Z;
	input wire D;
	input wire C;
	input wire B;
	input wire A;

endmodule // ym6045c_NOR4

module ym6045c_DFFSPOS (  C, D, nSET, nQ, Q);

	input wire C;
	input wire D;
	input wire nSET;
	output wire nQ;
	output wire Q;

endmodule // ym6045c_DFFSPOS

module ym6045c_JKFF (  C, K, J, nSET, nQ, Q);

	input wire C;
	input wire K;
	input wire J;
	input wire nSET;
	output wire nQ;
	output wire Q;

endmodule // ym6045c_JKFF

module ym6045c_DELAY (  Z, A);

	output wire Z;
	input wire A;

endmodule // ym6045c_DELAY

module ym6045c_AND4 (  Z, D, C, B, A);

	output wire Z;
	input wire D;
	input wire C;
	input wire B;
	input wire A;

endmodule // ym6045c_AND4

module ym6045c_OR (  A, Z, B);

	input wire A;
	output wire Z;
	input wire B;

endmodule // ym6045c_OR

module ym6045c_NOR (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // ym6045c_NOR

module ym6045c_OR3 (  Z, C, B, A);

	output wire Z;
	input wire C;
	input wire B;
	input wire A;

endmodule // ym6045c_OR3

module ym6045c_NAND4 (  B, C, A, D, Z);

	input wire B;
	input wire C;
	input wire A;
	input wire D;
	output wire Z;

endmodule // ym6045c_NAND4

module ym6045c_AND3 (  Z, C, B, A);

	output wire Z;
	input wire C;
	input wire B;
	input wire A;

endmodule // ym6045c_AND3

module ym6045c_DELAY_S (  Z, A);

	output wire Z;
	input wire A;

endmodule // ym6045c_DELAY_S

module ym6045c_NAND6 (  C, D, B, E, A, F, Z);

	input wire C;
	input wire D;
	input wire B;
	input wire E;
	input wire A;
	input wire F;
	output wire Z;

endmodule // ym6045c_NAND6

module ym6045c_OR4 (  Z, D, C, B, A);

	output wire Z;
	input wire D;
	input wire C;
	input wire B;
	input wire A;

endmodule // ym6045c_OR4

module ym6045c_DFFPOS (  nQ, Q, D, C);

	output wire nQ;
	output wire Q;
	input wire D;
	input wire C;

endmodule // ym6045c_DFFPOS

module ym6045c_NOR3 (  Z, C, B, A);

	output wire Z;
	input wire C;
	input wire B;
	input wire A;

endmodule // ym6045c_NOR3

module ym6045c_DFFRPOS (  nQ, Q, nRES, D, C);

	output wire nQ;
	output wire Q;
	input wire nRES;
	input wire D;
	input wire C;

endmodule // ym6045c_DFFRPOS

module ym6045c_MUX4BIT (  C, Z0, B1, A1, B2, A2, Z1, Z2, A3, B3, B4, A4, Z3);

	input wire C;
	output wire Z0;
	input wire B1;
	input wire A1;
	input wire B2;
	input wire A2;
	output wire Z1;
	output wire Z2;
	input wire A3;
	input wire B3;
	input wire B4;
	input wire A4;
	output wire Z3;

endmodule // ym6045c_MUX4BIT

module ym6045c_XNOR (  A, B, Z);

	input wire A;
	input wire B;
	output wire Z;

endmodule // ym6045c_XNOR

module ym6045c_MUX (  C, Z, A, B);

	input wire C;
	output wire Z;
	input wire A;
	input wire B;

endmodule // ym6045c_MUX

module ym6045c_OR8 (  A, E, B, F, Z, C, G, D, H);

	input wire A;
	input wire E;
	input wire B;
	input wire F;
	output wire Z;
	input wire C;
	input wire G;
	input wire D;
	input wire H;

endmodule // ym6045c_OR8

module ym6045c_SIPO_8BIT (  nRES, Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7, D, C);

	input wire nRES;
	output wire Q0;
	output wire Q1;
	output wire Q2;
	output wire Q3;
	output wire Q4;
	output wire Q5;
	output wire Q6;
	output wire Q7;
	input wire D;
	input wire C;

endmodule // ym6045c_SIPO_8BIT

module ym6045c_DEC_2TO4 (  A1, Z3, Z2, A0, Z0, Z1);

	input wire A1;
	output wire Z3;
	output wire Z2;
	input wire A0;
	output wire Z0;
	output wire Z1;

endmodule // ym6045c_DEC_2TO4

module ym6045c_OAI21 (  Z, A2, B, A1);

	output wire Z;
	input wire A2;
	input wire B;
	input wire A1;

endmodule // ym6045c_OAI21

module ym6045c_NOR8 (  A, B, C, D, Z, E, F, G, H);

	input wire A;
	input wire B;
	input wire C;
	input wire D;
	output wire Z;
	input wire E;
	input wire F;
	input wire G;
	input wire H;

endmodule // ym6045c_NOR8

module ym6045c_TFF (  Q, nQ, C, T);

	output wire Q;
	output wire nQ;
	input wire C;
	input wire T;

endmodule // ym6045c_TFF




