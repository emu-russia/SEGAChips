module VDP (  CH0_EN, CH0VOL[0], CH0VOL[1], CH1_EN, CH1VOL[0], CH1VOL[1], CH2_EN, CH2VOL[0], CH2VOL[1], CH3_EN, CH3VOL[0], CH3VOL[1], PSGDAC0[0], PSGDAC0[1], PSGDAC0[2], PSGDAC0[3], PSGDAC0[4], PSGDAC0[5], PSGDAC0[6], PSGDAC0[7], PSGDAC1[0], PSGDAC1[1], PSGDAC1[2], PSGDAC1[3], PSGDAC1[4], PSGDAC1[5], PSGDAC1[6], PSGDAC1[7], PSGDAC2[0], PSGDAC2[1], PSGDAC2[2], PSGDAC2[3], PSGDAC2[4], PSGDAC2[5], PSGDAC2[6], PSGDAC2[7], PSGDAC3[0], PSGDAC3[1], PSGDAC3[2], PSGDAC3[3], PSGDAC3[4], PSGDAC3[5], PSGDAC3[6], PSGDAC3[7], CAi[22], CAo[22], CA[19], DTACK_OUT, Z80_INT, RA[7], RA[6], RA[5], RA[4], RA[2], RA[1], RA[0], nRAS0, RA[3], nCAS0, nOE0, nLWR, nUWR, DTACK_IN, RnW, nLDS, nUDS, nAS, nM1, nWR, nRD, nIORQ, nILP2, nILP1, nINTAK, nMREQ, nBG, BGACK_OUT, BGACK_IN, nBR, VSYNC, nCSYNC, nCSYNC_IN, nHSYNC, nHSYNC_IN, DB[15], DB[14], DB[13], DB[12], DB[11], DB[10], DB[9], DB[8], DB[7], DB[6], DB[5], DB[4], DB[3], DB[2], DB[1], DB[0], CA[0], CA[1], CA[2], CA[3], CA[4], CA[5], CA[6], CA[7], CA[8], CA[9], CA[10], CA[11], CA[12], CA[13], CA[14], CA[15], CA[16], CA[17], CA[18], CA[20], CA[21], R_DAC[0], R_DAC[1], R_DAC[2], R_DAC[3], R_DAC[4], R_DAC[5], R_DAC[6], R_DAC[7], R_DAC[8], G_DAC[0], G_DAC[1], G_DAC[2], G_DAC[3], G_DAC[4], G_DAC[5], G_DAC[6], G_DAC[7], G_DAC[8], R_DAC[9], R_DAC[10], R_DAC[11], R_DAC[12], R_DAC[13], R_DAC[14], R_DAC[15], R_DAC[16], B_DAC[0], B_DAC[1], B_DAC[2], B_DAC[3], B_DAC[4], B_DAC[5], B_DAC[6], B_DAC[7], B_DAC[8], G_DAC[9], G_DAC[10], G_DAC[11], G_DAC[12], G_DAC[13], G_DAC[14], G_DAC[15], G_DAC[16], B_DAC[9], B_DAC[10], B_DAC[11], B_DAC[12], B_DAC[13], B_DAC[14], B_DAC[15], B_DAC[16], nOE1, nWE0, nWE1, nCAS1, nRAS1, AD_RD_DIR, nYS, nSC, nSE0_1, ADo[7], ADo[6], ADo[5], ADo[4], ADo[3], ADo[2], ADo[1], ADo[0], RDo[6], RDo[5], RDo[4], RDo[3], RDo[2], RDo[1], RDo[0], RDi[6], RDi[7], RDi[4], RDi[5], RDi[2], RDi[3], RDi[0], RDi[1], ADi[6], ADi[7], ADi[4], ADi[5], ADi[2], ADi[3], ADi[0], ADi[1], RDo[7], SD[7], SD[6], SD[5], SD[4], SD[3], SD[2], SD[1], SD[0], CLK1, CLK0, EDCLKi, EDCLKo, MCLK, SUB_CLK, nRES_PAD, 68kCLKi, EDCLKd, CA_PAD_DIR, DB_PAD_DIR, SEL0_M3, nPAL, nHL, SPA/Bo, SPA/Bi);

	output wire CH0_EN;
	output wire CH0VOL[0];
	output wire CH0VOL[1];
	output wire CH1_EN;
	output wire CH1VOL[0];
	output wire CH1VOL[1];
	output wire CH2_EN;
	output wire CH2VOL[0];
	output wire CH2VOL[1];
	output wire CH3_EN;
	output wire CH3VOL[0];
	output wire CH3VOL[1];
	output wire PSGDAC0[0];
	output wire PSGDAC0[1];
	output wire PSGDAC0[2];
	output wire PSGDAC0[3];
	output wire PSGDAC0[4];
	output wire PSGDAC0[5];
	output wire PSGDAC0[6];
	output wire PSGDAC0[7];
	output wire PSGDAC1[0];
	output wire PSGDAC1[1];
	output wire PSGDAC1[2];
	output wire PSGDAC1[3];
	output wire PSGDAC1[4];
	output wire PSGDAC1[5];
	output wire PSGDAC1[6];
	output wire PSGDAC1[7];
	output wire PSGDAC2[0];
	output wire PSGDAC2[1];
	output wire PSGDAC2[2];
	output wire PSGDAC2[3];
	output wire PSGDAC2[4];
	output wire PSGDAC2[5];
	output wire PSGDAC2[6];
	output wire PSGDAC2[7];
	output wire PSGDAC3[0];
	output wire PSGDAC3[1];
	output wire PSGDAC3[2];
	output wire PSGDAC3[3];
	output wire PSGDAC3[4];
	output wire PSGDAC3[5];
	output wire PSGDAC3[6];
	output wire PSGDAC3[7];
	input wire CAi[22];
	output wire CAo[22];
	output wire CA[19];
	output wire DTACK_OUT;
	output wire Z80_INT;
	output wire RA[7];
	output wire RA[6];
	output wire RA[5];
	output wire RA[4];
	output wire RA[2];
	output wire RA[1];
	output wire RA[0];
	output wire nRAS0;
	output wire RA[3];
	output wire nCAS0;
	output wire nOE0;
	output wire nLWR;
	output wire nUWR;
	input wire DTACK_IN;
	input wire RnW;
	input wire nLDS;
	input wire nUDS;
	input wire nAS;
	input wire nM1;
	input wire nWR;
	input wire nRD;
	input wire nIORQ;
	output wire nILP2;
	output wire nILP1;
	input wire nINTAK;
	input wire nMREQ;
	input wire nBG;
	output wire BGACK_OUT;
	input wire BGACK_IN;
	output wire nBR;
	output wire VSYNC;
	output wire nCSYNC;
	input wire nCSYNC_IN;
	output wire nHSYNC;
	input wire nHSYNC_IN;
	inout wire DB[15];
	inout wire DB[14];
	inout wire DB[13];
	inout wire DB[12];
	inout wire DB[11];
	inout wire DB[10];
	inout wire DB[9];
	inout wire DB[8];
	inout wire DB[7];
	inout wire DB[6];
	inout wire DB[5];
	inout wire DB[4];
	inout wire DB[3];
	inout wire DB[2];
	inout wire DB[1];
	inout wire DB[0];
	inout wire CA[0];
	inout wire CA[1];
	inout wire CA[2];
	inout wire CA[3];
	inout wire CA[4];
	inout wire CA[5];
	inout wire CA[6];
	inout wire CA[7];
	inout wire CA[8];
	inout wire CA[9];
	inout wire CA[10];
	inout wire CA[11];
	inout wire CA[12];
	inout wire CA[13];
	inout wire CA[14];
	inout wire CA[15];
	inout wire CA[16];
	inout wire CA[17];
	output wire CA[18];
	inout wire CA[20];
	inout wire CA[21];
	output wire R_DAC[0];
	output wire R_DAC[1];
	output wire R_DAC[2];
	output wire R_DAC[3];
	output wire R_DAC[4];
	output wire R_DAC[5];
	output wire R_DAC[6];
	output wire R_DAC[7];
	output wire R_DAC[8];
	output wire G_DAC[0];
	output wire G_DAC[1];
	output wire G_DAC[2];
	output wire G_DAC[3];
	output wire G_DAC[4];
	output wire G_DAC[5];
	output wire G_DAC[6];
	output wire G_DAC[7];
	output wire G_DAC[8];
	output wire R_DAC[9];
	output wire R_DAC[10];
	output wire R_DAC[11];
	output wire R_DAC[12];
	output wire R_DAC[13];
	output wire R_DAC[14];
	output wire R_DAC[15];
	output wire R_DAC[16];
	output wire B_DAC[0];
	output wire B_DAC[1];
	output wire B_DAC[2];
	output wire B_DAC[3];
	output wire B_DAC[4];
	output wire B_DAC[5];
	output wire B_DAC[6];
	output wire B_DAC[7];
	output wire B_DAC[8];
	output wire G_DAC[9];
	output wire G_DAC[10];
	output wire G_DAC[11];
	output wire G_DAC[12];
	output wire G_DAC[13];
	output wire G_DAC[14];
	output wire G_DAC[15];
	output wire G_DAC[16];
	output wire B_DAC[9];
	output wire B_DAC[10];
	output wire B_DAC[11];
	output wire B_DAC[12];
	output wire B_DAC[13];
	output wire B_DAC[14];
	output wire B_DAC[15];
	output wire B_DAC[16];
	output wire nOE1;
	output wire nWE0;
	output wire nWE1;
	output wire nCAS1;
	output wire nRAS1;
	output wire AD_RD_DIR;
	output wire nYS;
	output wire nSC;
	output wire nSE0_1;
	output wire ADo[7];
	output wire ADo[6];
	output wire ADo[5];
	output wire ADo[4];
	output wire ADo[3];
	output wire ADo[2];
	output wire ADo[1];
	output wire ADo[0];
	output wire RDo[6];
	output wire RDo[5];
	output wire RDo[4];
	output wire RDo[3];
	output wire RDo[2];
	output wire RDo[1];
	output wire RDo[0];
	input wire RDi[6];
	input wire RDi[7];
	input wire RDi[4];
	input wire RDi[5];
	input wire RDi[2];
	input wire RDi[3];
	input wire RDi[0];
	input wire RDi[1];
	input wire ADi[6];
	input wire ADi[7];
	input wire ADi[4];
	input wire ADi[5];
	input wire ADi[2];
	input wire ADi[3];
	input wire ADi[0];
	input wire ADi[1];
	output wire RDo[7];
	input wire SD[7];
	input wire SD[6];
	input wire SD[5];
	input wire SD[4];
	input wire SD[3];
	input wire SD[2];
	input wire SD[1];
	input wire SD[0];
	output wire CLK1;
	output wire CLK0;
	input wire EDCLKi;
	output wire EDCLKo;
	input wire MCLK;
	output wire SUB_CLK;
	input wire nRES_PAD;
	input wire 68kCLKi;
	output wire EDCLKd;
	output wire CA_PAD_DIR;
	output wire DB_PAD_DIR;
	input wire SEL0_M3;
	input wire nPAL;
	input wire nHL;
	output wire SPA/Bo;
	input wire SPA/Bi;

	// Wires

	wire w1;
	wire H40;
	wire w3;
	wire w4;
	wire w5;
	wire w6;
	wire w7;
	wire w8;
	wire w9;
	wire w10;
	wire w11;
	wire w12;
	wire w13;
	wire w14;
	wire w15;
	wire w16;
	wire w17;
	wire w18;
	wire w19;
	wire w20;
	wire w21;
	wire w22;
	wire w23;
	wire w24;
	wire w25;
	wire w26;
	wire w27;
	wire w28;
	wire w29;
	wire w30;
	wire w31;
	wire w32;
	wire w33;
	wire w34;
	wire w35;
	wire w36;
	wire w37;
	wire w38;
	wire w39;
	wire w40;
	wire w41;
	wire w42;
	wire w43;
	wire w44;
	wire w45;
	wire w46;
	wire w47;
	wire w48;
	wire ODD_EVEN;
	wire w50;
	wire w51;
	wire w52;
	wire w53;
	wire w54;
	wire w55;
	wire w56;
	wire w57;
	wire w58;
	wire w59;
	wire FIFOo[7];
	wire FIFOo[6];
	wire FIFOo[5];
	wire FIFOo[4];
	wire FIFOo[3];
	wire FIFOo[2];
	wire FIFOo[1];
	wire FIFOo[0];
	wire w68;
	wire w69;
	wire w70;
	wire w71;
	wire w72;
	wire w73;
	wire w74;
	wire w75;
	wire w76;
	wire w77;
	wire w78;
	wire w79;
	wire w80;
	wire w81;
	wire w82;
	wire w83;
	wire w84;
	wire w85;
	wire w86;
	wire w87;
	wire w88;
	wire w89;
	wire w90;
	wire w91;
	wire w92;
	wire w93;
	wire w94;
	wire w95;
	wire w96;
	wire VPOS[9];
	wire w98;
	wire w99;
	wire w100;
	wire w101;
	wire HPOS[0];
	wire w103;
	wire w104;
	wire w105;
	wire w106;
	wire w107;
	wire w108;
	wire w109;
	wire w110;
	wire w111;
	wire VPOS[8];
	wire w113;
	wire w114;
	wire w115;
	wire w116;
	wire w117;
	wire w118;
	wire w119;
	wire w120;
	wire w121;
	wire w122;
	wire w123;
	wire w124;
	wire w125;
	wire w126;
	wire w127;
	wire w128;
	wire w129;
	wire AD_DATA[7];
	wire AD_DATA[6];
	wire AD_DATA[4];
	wire RD_DATA[2];
	wire RD_DATA[1];
	wire RD_DATA[0];
	wire AD_DATA[5];
	wire w137;
	wire w138;
	wire DCLK1;
	wire DCLK2;
	wire nDCLK1;
	wire nDCLK2;
	wire HCLK1;
	wire HCLK2;
	wire nHCLK1;
	wire nHCLK2;
	wire SYSRES;
	wire DB[0];
	wire DB[1];
	wire DB[2];
	wire DB[3];
	wire DB[4];
	wire DB[5];
	wire DB[6];
	wire DB[7];
	wire DB[8];
	wire DB[9];
	wire AD_DATA[3];
	wire AD_DATA[2];
	wire AD_DATA[1];
	wire AD_DATA[0];
	wire DB[14];
	wire DB[13];
	wire DB[12];
	wire DB[11];
	wire DB[10];
	wire M5;
	wire w168;
	wire w169;
	wire w170;
	wire w171;
	wire w172;
	wire w173;
	wire w174;
	wire HPOS[1];
	wire w176;
	wire w177;
	wire w178;
	wire w179;
	wire w180;
	wire w181;
	wire w182;
	wire w183;
	wire w184;
	wire w185;
	wire w186;
	wire w187;
	wire w188;
	wire VPOS[2];
	wire HPOS[3];
	wire w191;
	wire w192;
	wire w193;
	wire w194;
	wire w195;
	wire w196;
	wire w197;
	wire w198;
	wire w199;
	wire w200;
	wire w201;
	wire w202;
	wire w203;
	wire VPOS[4];
	wire w205;
	wire RD_DATA[4];
	wire HPOS[5];
	wire w208;
	wire w209;
	wire w210;
	wire w211;
	wire w212;
	wire w213;
	wire w214;
	wire w215;
	wire w216;
	wire w217;
	wire w218;
	wire w219;
	wire w220;
	wire RD_DATA[6];
	wire HPOS[7];
	wire w223;
	wire w224;
	wire w225;
	wire w226;
	wire w227;
	wire w228;
	wire w229;
	wire w230;
	wire w231;
	wire w232;
	wire w233;
	wire w234;
	wire w235;
	wire w236;
	wire w237;
	wire w238;
	wire w239;
	wire w240;
	wire w241;
	wire w242;
	wire w243;
	wire w244;
	wire w245;
	wire w246;
	wire w247;
	wire w248;
	wire w249;
	wire w250;
	wire w251;
	wire w252;
	wire w253;
	wire w254;
	wire w255;
	wire w256;
	wire w257;
	wire w258;
	wire w259;
	wire w260;
	wire w261;
	wire w262;
	wire w263;
	wire w264;
	wire w265;
	wire w266;
	wire w267;
	wire w268;
	wire w269;
	wire w270;
	wire w271;
	wire w272;
	wire w273;
	wire w274;
	wire w275;
	wire w276;
	wire w277;
	wire w278;
	wire w279;
	wire w280;
	wire w281;
	wire w282;
	wire w283;
	wire w284;
	wire w285;
	wire w286;
	wire w287;
	wire w288;
	wire w289;
	wire w290;
	wire w291;
	wire w292;
	wire w293;
	wire w294;
	wire w295;
	wire w296;
	wire w297;
	wire w298;
	wire w299;
	wire w300;
	wire w301;
	wire w302;
	wire w303;
	wire w304;
	wire w305;
	wire w306;
	wire HPOS[2];
	wire VPOS[1];
	wire w309;
	wire w310;
	wire w311;
	wire w312;
	wire w313;
	wire w314;
	wire w315;
	wire w316;
	wire w317;
	wire w318;
	wire w319;
	wire VPOS[3];
	wire w321;
	wire HPOS[4];
	wire w323;
	wire w324;
	wire w325;
	wire w326;
	wire w327;
	wire w328;
	wire w329;
	wire w330;
	wire w331;
	wire w332;
	wire w333;
	wire w334;
	wire w335;
	wire VPOS[5];
	wire RD_DATA[5];
	wire HPOS[6];
	wire w339;
	wire w340;
	wire w341;
	wire w342;
	wire w343;
	wire w344;
	wire w345;
	wire w346;
	wire w347;
	wire w348;
	wire w349;
	wire w350;
	wire w351;
	wire HPOS[8];
	wire VPOS[7];
	wire DB[15];
	wire w355;
	wire w356;
	wire w357;
	wire w358;
	wire w359;
	wire w360;
	wire w361;
	wire w362;
	wire w363;
	wire w364;
	wire w365;
	wire w366;
	wire w367;
	wire w368;
	wire w369;
	wire w370;
	wire w371;
	wire w372;
	wire w373;
	wire w374;
	wire w375;
	wire w376;
	wire w377;
	wire w378;
	wire w379;
	wire w380;
	wire w381;
	wire w382;
	wire w383;
	wire w384;
	wire w385;
	wire w386;
	wire w387;
	wire w388;
	wire w389;
	wire w390;
	wire w391;
	wire w392;
	wire w393;
	wire w394;
	wire w395;
	wire w396;
	wire w397;
	wire w398;
	wire w399;
	wire w400;
	wire w401;
	wire w402;
	wire w403;
	wire w404;
	wire w405;
	wire w406;
	wire w407;
	wire w408;
	wire w409;
	wire w410;
	wire w411;
	wire w412;
	wire w413;
	wire w414;
	wire w415;
	wire w416;
	wire w417;
	wire w418;
	wire w419;
	wire w420;
	wire w421;
	wire w422;
	wire w423;
	wire w424;
	wire w425;
	wire w426;
	wire w427;
	wire w428;
	wire w429;
	wire w430;
	wire w431;
	wire w432;
	wire 128k;
	wire w434;
	wire w435;
	wire w436;
	wire w437;
	wire w438;
	wire w439;
	wire w440;
	wire w441;
	wire w442;
	wire w443;
	wire w444;
	wire w445;
	wire w446;
	wire w447;
	wire w448;
	wire w449;
	wire w450;
	wire w451;
	wire w452;
	wire w453;
	wire w454;
	wire w455;
	wire w456;
	wire w457;
	wire w458;
	wire w459;
	wire w460;
	wire w461;
	wire w462;
	wire w463;
	wire w464;
	wire w465;
	wire w466;
	wire w467;
	wire w468;
	wire w469;
	wire CA[0];
	wire w471;
	wire w472;
	wire w473;
	wire w474;
	wire w475;
	wire w476;
	wire w477;
	wire w478;
	wire w479;
	wire w480;
	wire w481;
	wire w482;
	wire w483;
	wire w484;
	wire w485;
	wire w486;
	wire w487;
	wire w488;
	wire w489;
	wire w490;
	wire w491;
	wire w492;
	wire w493;
	wire w494;
	wire w495;
	wire w496;
	wire w497;
	wire w498;
	wire w499;
	wire w500;
	wire w501;
	wire w502;
	wire w503;
	wire w504;
	wire w505;
	wire w506;
	wire w507;
	wire w508;
	wire w509;
	wire w510;
	wire w511;
	wire w512;
	wire w513;
	wire w514;
	wire w515;
	wire w516;
	wire w517;
	wire w518;
	wire w519;
	wire w520;
	wire w521;
	wire w522;
	wire w523;
	wire w524;
	wire w525;
	wire w526;
	wire w527;
	wire w528;
	wire w529;
	wire w530;
	wire w531;
	wire w532;
	wire w533;
	wire w534;
	wire w535;
	wire w536;
	wire w537;
	wire w538;
	wire w539;
	wire w540;
	wire w541;
	wire w542;
	wire w543;
	wire w544;
	wire w545;
	wire w546;
	wire w547;
	wire w548;
	wire w549;
	wire w550;
	wire w551;
	wire w552;
	wire w553;
	wire w554;
	wire w555;
	wire w556;
	wire w557;
	wire w558;
	wire w559;
	wire w560;
	wire VRAMA[0];
	wire w562;
	wire w563;
	wire w564;
	wire w565;
	wire w566;
	wire w567;
	wire w568;
	wire w569;
	wire w570;
	wire w571;
	wire w572;
	wire w573;
	wire w574;
	wire w575;
	wire w576;
	wire w577;
	wire w578;
	wire w579;
	wire w580;
	wire w581;
	wire w582;
	wire w583;
	wire w584;
	wire w585;
	wire w586;
	wire w587;
	wire w588;
	wire w589;
	wire w590;
	wire w591;
	wire w592;
	wire w593;
	wire w594;
	wire w595;
	wire w596;
	wire w597;
	wire DMA_BUSY;
	wire w599;
	wire w600;
	wire w601;
	wire w602;
	wire w603;
	wire w604;
	wire w605;
	wire REG_BUS[0];
	wire w607;
	wire w608;
	wire w609;
	wire w610;
	wire REG_BUS[7];
	wire VRAMA[8];
	wire w613;
	wire w614;
	wire w615;
	wire w616;
	wire w617;
	wire w618;
	wire w619;
	wire w620;
	wire w621;
	wire w622;
	wire w623;
	wire w624;
	wire w625;
	wire w626;
	wire w627;
	wire w628;
	wire w629;
	wire w630;
	wire w631;
	wire w632;
	wire w633;
	wire w634;
	wire w635;
	wire w636;
	wire CA[8];
	wire CA[7];
	wire w639;
	wire w640;
	wire w641;
	wire w642;
	wire w643;
	wire w644;
	wire w645;
	wire w646;
	wire w647;
	wire w648;
	wire w649;
	wire w650;
	wire w651;
	wire CA[9];
	wire w653;
	wire VRAMA[7];
	wire w655;
	wire REG_BUS[6];
	wire VRAMA[9];
	wire w658;
	wire CA[6];
	wire w660;
	wire w661;
	wire w662;
	wire w663;
	wire w664;
	wire w665;
	wire w666;
	wire w667;
	wire w668;
	wire w669;
	wire w670;
	wire w671;
	wire w672;
	wire w673;
	wire w674;
	wire REG_BUS[5];
	wire VRAMA[10];
	wire VRAMA[6];
	wire w678;
	wire REG_BUS[1];
	wire w680;
	wire w681;
	wire w682;
	wire w683;
	wire CA[10];
	wire w685;
	wire w686;
	wire w687;
	wire w688;
	wire w689;
	wire w690;
	wire w691;
	wire REG_BUS[2];
	wire w693;
	wire CA[11];
	wire w695;
	wire w696;
	wire w697;
	wire w698;
	wire w699;
	wire w700;
	wire w701;
	wire w702;
	wire w703;
	wire w704;
	wire VRAMA[5];
	wire w706;
	wire w707;
	wire VRAMA[11];
	wire CA[5];
	wire w710;
	wire w711;
	wire w712;
	wire REG_BUS[3];
	wire VRAMA[12];
	wire VRAMA[4];
	wire w716;
	wire w717;
	wire w718;
	wire REG_BUS[4];
	wire w720;
	wire CA[12];
	wire w722;
	wire w723;
	wire CA[4];
	wire w725;
	wire w726;
	wire w727;
	wire w728;
	wire CA[19];
	wire w730;
	wire w731;
	wire w732;
	wire w733;
	wire w734;
	wire VRAMA[13];
	wire w736;
	wire w737;
	wire w738;
	wire VRAMA[3];
	wire CA[3];
	wire w741;
	wire w742;
	wire CA[13];
	wire CA[20];
	wire w745;
	wire w746;
	wire w747;
	wire w748;
	wire w749;
	wire w750;
	wire VRAMA[14];
	wire VRAMA[2];
	wire w753;
	wire w754;
	wire w755;
	wire w756;
	wire w757;
	wire CA[2];
	wire w759;
	wire w760;
	wire w761;
	wire CA[21];
	wire w763;
	wire w764;
	wire w765;
	wire w766;
	wire w767;
	wire CA[14];
	wire w769;
	wire w770;
	wire VRAMA[15];
	wire CA[15];
	wire VRAMA[1];
	wire w774;
	wire w775;
	wire w776;
	wire w777;
	wire w778;
	wire w779;
	wire w780;
	wire w781;
	wire w782;
	wire w783;
	wire w784;
	wire CA[17];
	wire CA[1];
	wire VRAMA[16];
	wire w788;
	wire w789;
	wire CA[16];
	wire w791;
	wire w792;
	wire w793;
	wire w794;
	wire w795;
	wire w796;
	wire w797;
	wire w798;
	wire w799;
	wire w800;
	wire w801;
	wire w802;
	wire w803;
	wire w804;
	wire w805;
	wire w806;
	wire w807;
	wire w808;
	wire w809;
	wire w810;
	wire w811;
	wire w812;
	wire w813;
	wire w814;
	wire w815;
	wire w816;
	wire w817;
	wire w818;
	wire w819;
	wire w820;
	wire w821;
	wire w822;
	wire w823;
	wire w824;
	wire w825;
	wire w826;
	wire w827;
	wire w828;
	wire w829;
	wire w830;
	wire w831;
	wire w832;
	wire w833;
	wire w834;
	wire w835;
	wire w836;
	wire w837;
	wire w838;
	wire w839;
	wire w840;
	wire w841;
	wire w842;
	wire w843;
	wire w844;
	wire w845;
	wire w846;
	wire w847;
	wire w848;
	wire w849;
	wire w850;
	wire w851;
	wire w852;
	wire w853;
	wire w854;
	wire w855;
	wire w856;
	wire w857;
	wire w858;
	wire w859;
	wire w860;
	wire w861;
	wire w862;
	wire w863;
	wire w864;
	wire w865;
	wire w866;
	wire w867;
	wire w868;
	wire w869;
	wire w870;
	wire w871;
	wire w872;
	wire w873;
	wire w874;
	wire w875;
	wire w876;
	wire w877;
	wire w878;
	wire w879;
	wire w880;
	wire w881;
	wire w882;
	wire w883;
	wire w884;
	wire w885;
	wire w886;
	wire w887;
	wire w888;
	wire w889;
	wire w890;
	wire w891;
	wire w892;
	wire w893;
	wire w894;
	wire w895;
	wire w896;
	wire w897;
	wire w898;
	wire w899;
	wire w900;
	wire w901;
	wire w902;
	wire w903;
	wire w904;
	wire w905;
	wire w906;
	wire w907;
	wire w908;
	wire w909;
	wire w910;
	wire w911;
	wire w912;
	wire w913;
	wire w914;
	wire w915;
	wire w916;
	wire w917;
	wire w918;
	wire w919;
	wire w920;
	wire w921;
	wire w922;
	wire w923;
	wire w924;
	wire w925;
	wire w926;
	wire w927;
	wire w928;
	wire w929;
	wire w930;
	wire w931;
	wire w932;
	wire w933;
	wire w934;
	wire w935;
	wire w936;
	wire w937;
	wire w938;
	wire w939;
	wire w940;
	wire w941;
	wire w942;
	wire w943;
	wire w944;
	wire w945;
	wire w946;
	wire w947;
	wire w948;
	wire w949;
	wire w950;
	wire w951;
	wire w952;
	wire w953;
	wire w954;
	wire w955;
	wire w956;
	wire w957;
	wire w958;
	wire w959;
	wire w960;
	wire w961;
	wire w962;
	wire w963;
	wire w964;
	wire w965;
	wire w966;
	wire w967;
	wire w968;
	wire w969;
	wire w970;
	wire w971;
	wire w972;
	wire w973;
	wire w974;
	wire w975;
	wire w976;
	wire w977;
	wire w978;
	wire w979;
	wire w980;
	wire w981;
	wire w982;
	wire w983;
	wire w984;
	wire w985;
	wire w986;
	wire w987;
	wire w988;
	wire w989;
	wire w990;
	wire w991;
	wire w992;
	wire w993;
	wire w994;
	wire w995;
	wire w996;
	wire w997;
	wire w998;
	wire w999;
	wire w1000;
	wire w1001;
	wire w1002;
	wire w1003;
	wire w1004;
	wire w1005;
	wire w1006;
	wire w1007;
	wire w1008;
	wire w1009;
	wire w1010;
	wire w1011;
	wire w1012;
	wire w1013;
	wire w1014;
	wire w1015;
	wire w1016;
	wire w1017;
	wire w1018;
	wire w1019;
	wire w1020;
	wire w1021;
	wire w1022;
	wire w1023;
	wire w1024;
	wire w1025;
	wire w1026;
	wire w1027;
	wire w1028;
	wire w1029;
	wire w1030;
	wire w1031;
	wire w1032;
	wire w1033;
	wire w1034;
	wire w1035;
	wire w1036;
	wire w1037;
	wire w1038;
	wire w1039;
	wire w1040;
	wire w1041;
	wire w1042;
	wire w1043;
	wire w1044;
	wire w1045;
	wire w1046;
	wire w1047;
	wire w1048;
	wire w1049;
	wire w1050;
	wire w1051;
	wire w1052;
	wire PSG_Z80_CLK;
	wire LS0;
	wire w1055;
	wire VPOS[0];
	wire w1057;
	wire w1058;
	wire w1059;
	wire w1060;
	wire w1061;
	wire w1062;
	wire w1063;
	wire w1064;
	wire w1065;
	wire w1066;
	wire w1067;
	wire w1068;
	wire w1069;
	wire w1070;
	wire w1071;
	wire w1072;
	wire w1073;
	wire w1074;
	wire w1075;
	wire w1076;
	wire w1077;
	wire COL[0];
	wire COL[1];
	wire COL[2];
	wire COL[3];
	wire COL[4];
	wire COL[5];
	wire COL[6];
	wire w1085;
	wire w1086;
	wire w1087;
	wire w1088;
	wire w1089;
	wire w1090;
	wire w1091;
	wire w1092;
	wire w1093;
	wire w1094;
	wire w1095;
	wire w1096;
	wire w1097;
	wire w1098;
	wire w1099;
	wire w1100;
	wire w1101;
	wire w1102;
	wire w1103;
	wire w1104;
	wire w1105;
	wire w1106;
	wire w1107;
	wire w1108;
	wire w1109;
	wire w1110;
	wire w1111;
	wire w1112;
	wire w1113;
	wire w1114;
	wire w1115;
	wire w1116;
	wire w1117;
	wire w1118;
	wire w1119;
	wire w1120;
	wire w1121;
	wire w1122;
	wire w1123;
	wire w1124;
	wire w1125;
	wire w1126;
	wire w1127;
	wire w1128;
	wire w1129;
	wire w1130;
	wire w1131;
	wire w1132;
	wire w1133;
	wire w1134;
	wire w1135;
	wire w1136;
	wire w1137;
	wire w1138;
	wire w1139;
	wire w1140;
	wire w1141;
	wire w1142;
	wire PSG_TEST_OE;
	wire w1144;
	wire w1145;
	wire w1146;
	wire w1147;
	wire w1148;
	wire w1149;
	wire w1150;
	wire w1151;
	wire w1152;
	wire w1153;
	wire w1154;
	wire w1155;
	wire w1156;
	wire w1157;
	wire w1158;
	wire w1159;
	wire w1160;
	wire w1161;
	wire w1162;
	wire w1163;
	wire w1164;
	wire w1165;
	wire w1166;
	wire w1167;
	wire w1168;
	wire w1169;
	wire w1170;
	wire w1171;
	wire w1172;
	wire w1173;
	wire w1174;
	wire w1175;
	wire w1176;
	wire w1177;
	wire w1178;
	wire w1179;
	wire w1180;
	wire w1181;
	wire w1182;
	wire w1183;
	wire w1184;
	wire w1185;
	wire w1186;
	wire w1187;
	wire w1188;
	wire w1189;
	wire w1190;
	wire w1191;
	wire w1192;
	wire w1193;
	wire w1194;
	wire w1195;
	wire PAL;
	wire w1197;
	wire w1198;
	wire w1199;
	wire w1200;
	wire w1201;
	wire w1202;
	wire w1203;
	wire w1204;
	wire w1205;
	wire w1206;
	wire w1207;
	wire w1208;
	wire w1209;
	wire w1210;
	wire w1211;
	wire w1212;
	wire w1213;
	wire w1214;
	wire w1215;
	wire w1216;
	wire w1217;
	wire w1218;
	wire w1219;
	wire w1220;
	wire w1221;
	wire w1222;
	wire w1223;
	wire w1224;
	wire w1225;
	wire w1226;
	wire w1227;
	wire w1228;
	wire w1229;
	wire w1230;
	wire w1231;
	wire w1232;
	wire w1233;
	wire w1234;
	wire w1235;
	wire w1236;
	wire w1237;
	wire w1238;
	wire w1239;
	wire w1240;
	wire w1241;
	wire w1242;
	wire w1243;
	wire w1244;
	wire w1245;
	wire w1246;
	wire w1247;
	wire w1248;
	wire w1249;
	wire w1250;
	wire w1251;
	wire w1252;
	wire w1253;
	wire w1254;
	wire w1255;
	wire w1256;
	wire w1257;
	wire w1258;
	wire w1259;
	wire w1260;
	wire w1261;
	wire w1262;
	wire w1263;
	wire w1264;
	wire w1265;
	wire w1266;
	wire w1267;
	wire w1268;
	wire w1269;
	wire w1270;
	wire w1271;
	wire w1272;
	wire w1273;
	wire w1274;
	wire w1275;
	wire w1276;
	wire w1277;
	wire w1278;
	wire w1279;
	wire w1280;
	wire w1281;
	wire w1282;
	wire w1283;
	wire w1284;
	wire w1285;
	wire w1286;
	wire w1287;
	wire w1288;
	wire w1289;
	wire w1290;
	wire w1291;
	wire w1292;
	wire w1293;
	wire w1294;
	wire w1295;
	wire w1296;
	wire w1297;
	wire w1298;
	wire w1299;
	wire w1300;
	wire w1301;
	wire w1302;
	wire w1303;
	wire w1304;
	wire w1305;
	wire w1306;
	wire w1307;
	wire w1308;
	wire w1309;
	wire w1310;
	wire w1311;
	wire w1312;
	wire w1313;
	wire w1314;
	wire w1315;
	wire w1316;
	wire w1317;
	wire w1318;
	wire w1319;
	wire w1320;
	wire w1321;
	wire w1322;
	wire w1323;
	wire w1324;
	wire w1325;
	wire w1326;
	wire w1327;
	wire w1328;
	wire w1329;
	wire w1330;
	wire w1331;
	wire w1332;
	wire w1333;
	wire w1334;
	wire w1335;
	wire w1336;
	wire w1337;
	wire w1338;
	wire w1339;
	wire w1340;
	wire w1341;
	wire w1342;
	wire w1343;
	wire w1344;
	wire w1345;
	wire w1346;
	wire w1347;
	wire w1348;
	wire w1349;
	wire w1350;
	wire w1351;
	wire w1352;
	wire w1353;
	wire w1354;
	wire w1355;
	wire w1356;
	wire w1357;
	wire w1358;
	wire w1359;
	wire w1360;
	wire w1361;
	wire w1362;
	wire w1363;
	wire w1364;
	wire w1365;
	wire w1366;
	wire w1367;
	wire w1368;
	wire w1369;
	wire w1370;
	wire w1371;
	wire w1372;
	wire w1373;
	wire w1374;
	wire w1375;
	wire w1376;
	wire w1377;
	wire w1378;
	wire w1379;
	wire w1380;
	wire w1381;
	wire w1382;
	wire w1383;
	wire w1384;
	wire w1385;
	wire w1386;
	wire VRAM_REFRESH;
	wire w1388;
	wire w1389;
	wire w1390;
	wire w1391;
	wire w1392;
	wire w1393;
	wire w1394;
	wire w1395;
	wire w1396;
	wire w1397;
	wire w1398;
	wire w1399;
	wire w1400;
	wire w1401;
	wire w1402;
	wire w1403;
	wire w1404;
	wire w1405;
	wire w1406;
	wire w1407;
	wire w1408;
	wire w1409;
	wire w1410;
	wire w1411;
	wire w1412;
	wire w1413;
	wire w1414;
	wire w1415;
	wire w1416;
	wire w1417;
	wire w1418;
	wire w1419;
	wire w1420;
	wire w1421;
	wire w1422;
	wire w1423;
	wire w1424;
	wire w1425;
	wire w1426;
	wire w1427;
	wire w1428;
	wire w1429;
	wire w1430;
	wire w1431;
	wire w1432;
	wire w1433;
	wire w1434;
	wire w1435;
	wire w1436;
	wire w1437;
	wire w1438;
	wire w1439;
	wire w1440;
	wire w1441;
	wire w1442;
	wire w1443;
	wire w1444;
	wire w1445;
	wire w1446;
	wire w1447;
	wire w1448;
	wire w1449;
	wire w1450;
	wire w1451;
	wire w1452;
	wire w1453;
	wire w1454;
	wire w1455;
	wire w1456;
	wire w1457;
	wire w1458;
	wire w1459;
	wire w1460;
	wire w1461;
	wire w1462;
	wire w1463;
	wire w1464;
	wire w1465;
	wire w1466;
	wire w1467;
	wire w1468;
	wire w1469;
	wire w1470;
	wire w1471;
	wire w1472;
	wire w1473;
	wire w1474;
	wire w1475;
	wire w1476;
	wire w1477;
	wire w1478;
	wire w1479;
	wire w1480;
	wire w1481;
	wire w1482;
	wire w1483;
	wire w1484;
	wire w1485;
	wire w1486;
	wire w1487;
	wire w1488;
	wire w1489;
	wire w1490;
	wire w1491;
	wire w1492;
	wire w1493;
	wire w1494;
	wire w1495;
	wire w1496;
	wire w1497;
	wire w1498;
	wire w1499;
	wire CA[18];
	wire w1501;
	wire w1502;
	wire w1503;
	wire w1504;
	wire w1505;
	wire w1506;
	wire w1507;
	wire w1508;
	wire w1509;
	wire w1510;
	wire w1511;
	wire w1512;
	wire w1513;
	wire w1514;
	wire w1515;
	wire w1516;
	wire w1517;
	wire w1518;
	wire w1519;
	wire w1520;
	wire w1521;
	wire w1522;
	wire w1523;
	wire w1524;
	wire w1525;
	wire w1526;
	wire w1527;
	wire w1528;
	wire w1529;
	wire w1530;
	wire w1531;
	wire w1532;
	wire w1533;
	wire w1534;
	wire w1535;
	wire w1536;
	wire w1537;
	wire w1538;
	wire w1539;
	wire w1540;
	wire w1541;
	wire w1542;
	wire w1543;
	wire w1544;
	wire w1545;
	wire w1546;
	wire w1547;
	wire w1548;
	wire w1549;
	wire w1550;
	wire w1551;
	wire w1552;
	wire w1553;
	wire w1554;
	wire w1555;
	wire w1556;
	wire w1557;
	wire w1558;
	wire w1559;
	wire w1560;
	wire w1561;
	wire VPOS[6];
	wire w1563;
	wire w1564;
	wire w1565;
	wire w1566;
	wire w1567;
	wire w1568;
	wire w1569;
	wire w1570;
	wire w1571;
	wire w1572;
	wire w1573;
	wire w1574;
	wire w1575;
	wire w1576;
	wire w1577;
	wire w1578;
	wire w1579;
	wire w1580;
	wire w1581;
	wire w1582;
	wire w1583;
	wire w1584;
	wire w1585;
	wire w1586;
	wire w1587;
	wire w1588;
	wire w1589;
	wire w1590;
	wire w1591;
	wire w1592;
	wire w1593;
	wire w1594;
	wire w1595;
	wire w1596;
	wire w1597;
	wire w1598;
	wire w1599;
	wire w1600;
	wire w1601;
	wire w1602;
	wire w1603;
	wire w1604;
	wire w1605;
	wire w1606;
	wire w1607;
	wire w1608;
	wire w1609;
	wire w1610;
	wire w1611;
	wire w1612;
	wire w1613;
	wire w1614;
	wire w1615;
	wire w1616;
	wire w1617;
	wire w1618;
	wire w1619;
	wire w1620;
	wire w1621;
	wire w1622;
	wire w1623;
	wire w1624;
	wire w1625;
	wire w1626;
	wire w1627;
	wire w1628;
	wire w1629;
	wire w1630;
	wire w1631;
	wire w1632;
	wire w1633;
	wire w1634;
	wire w1635;
	wire w1636;
	wire w1637;
	wire w1638;
	wire w1639;
	wire w1640;
	wire w1641;
	wire w1642;
	wire w1643;
	wire w1644;
	wire w1645;
	wire w1646;
	wire w1647;
	wire w1648;
	wire w1649;
	wire w1650;
	wire w1651;
	wire w1652;
	wire w1653;
	wire w1654;
	wire w1655;
	wire w1656;
	wire w1657;
	wire w1658;
	wire w1659;
	wire w1660;
	wire w1661;
	wire w1662;
	wire w1663;
	wire w1664;
	wire w1665;
	wire w1666;
	wire w1667;
	wire w1668;
	wire w1669;
	wire w1670;
	wire w1671;
	wire w1672;
	wire w1673;
	wire w1674;
	wire w1675;
	wire w1676;
	wire w1677;
	wire w1678;
	wire w1679;
	wire w1680;
	wire w1681;
	wire w1682;
	wire w1683;
	wire w1684;
	wire w1685;
	wire w1686;
	wire w1687;
	wire w1688;
	wire w1689;
	wire w1690;
	wire w1691;
	wire w1692;
	wire w1693;
	wire w1694;
	wire w1695;
	wire w1696;
	wire w1697;
	wire w1698;
	wire w1699;
	wire w1700;
	wire w1701;
	wire w1702;
	wire w1703;
	wire w1704;
	wire w1705;
	wire w1706;
	wire w1707;
	wire w1708;
	wire w1709;
	wire w1710;
	wire w1711;
	wire w1712;
	wire w1713;
	wire w1714;
	wire w1715;
	wire w1716;
	wire w1717;
	wire w1718;
	wire w1719;
	wire w1720;
	wire w1721;
	wire w1722;
	wire w1723;
	wire w1724;
	wire w1725;
	wire w1726;
	wire w1727;
	wire w1728;
	wire w1729;
	wire w1730;
	wire w1731;
	wire w1732;
	wire w1733;
	wire w1734;
	wire w1735;
	wire w1736;
	wire w1737;
	wire w1738;
	wire w1739;
	wire w1740;
	wire w1741;
	wire w1742;
	wire w1743;
	wire w1744;
	wire w1745;
	wire w1746;
	wire w1747;
	wire w1748;
	wire w1749;
	wire w1750;
	wire w1751;
	wire w1752;
	wire w1753;
	wire w1754;
	wire w1755;
	wire w1756;
	wire w1757;
	wire w1758;
	wire w1759;
	wire w1760;
	wire w1761;
	wire w1762;
	wire w1763;
	wire w1764;
	wire w1765;
	wire w1766;
	wire w1767;
	wire w1768;
	wire w1769;
	wire w1770;
	wire w1771;
	wire w1772;
	wire w1773;
	wire w1774;
	wire w1775;
	wire w1776;
	wire w1777;
	wire w1778;
	wire w1779;
	wire w1780;
	wire w1781;
	wire w1782;
	wire w1783;
	wire w1784;
	wire w1785;
	wire w1786;
	wire w1787;
	wire w1788;
	wire w1789;
	wire w1790;
	wire w1791;
	wire w1792;
	wire w1793;
	wire w1794;
	wire w1795;
	wire w1796;
	wire w1797;
	wire w1798;
	wire w1799;
	wire w1800;
	wire w1801;
	wire w1802;
	wire w1803;
	wire w1804;
	wire w1805;
	wire w1806;
	wire w1807;
	wire w1808;
	wire w1809;
	wire w1810;
	wire w1811;
	wire w1812;
	wire w1813;
	wire w1814;
	wire w1815;
	wire w1816;
	wire w1817;
	wire w1818;
	wire w1819;
	wire w1820;
	wire w1821;
	wire w1822;
	wire w1823;
	wire w1824;
	wire w1825;
	wire w1826;
	wire w1827;
	wire w1828;
	wire w1829;
	wire w1830;
	wire w1831;
	wire w1832;
	wire w1833;
	wire w1834;
	wire w1835;
	wire w1836;
	wire w1837;
	wire w1838;
	wire w1839;
	wire w1840;
	wire w1841;
	wire w1842;
	wire w1843;
	wire w1844;
	wire w1845;
	wire w1846;
	wire w1847;
	wire w1848;
	wire w1849;
	wire w1850;
	wire w1851;
	wire w1852;
	wire w1853;
	wire w1854;
	wire w1855;
	wire w1856;
	wire w1857;
	wire w1858;
	wire w1859;
	wire w1860;
	wire w1861;
	wire w1862;
	wire w1863;
	wire w1864;
	wire w1865;
	wire w1866;
	wire w1867;
	wire w1868;
	wire w1869;
	wire w1870;
	wire w1871;
	wire w1872;
	wire w1873;
	wire w1874;
	wire w1875;
	wire w1876;
	wire w1877;
	wire w1878;
	wire w1879;
	wire w1880;
	wire w1881;
	wire w1882;
	wire w1883;
	wire w1884;
	wire w1885;
	wire w1886;
	wire w1887;
	wire w1888;
	wire w1889;
	wire w1890;
	wire w1891;
	wire w1892;
	wire w1893;
	wire w1894;
	wire w1895;
	wire w1896;
	wire w1897;
	wire w1898;
	wire w1899;
	wire w1900;
	wire w1901;
	wire w1902;
	wire w1903;
	wire w1904;
	wire w1905;
	wire w1906;
	wire w1907;
	wire w1908;
	wire w1909;
	wire w1910;
	wire w1911;
	wire w1912;
	wire w1913;
	wire w1914;
	wire w1915;
	wire w1916;
	wire w1917;
	wire w1918;
	wire w1919;
	wire w1920;
	wire w1921;
	wire w1922;
	wire w1923;
	wire w1924;
	wire w1925;
	wire w1926;
	wire w1927;
	wire w1928;
	wire w1929;
	wire w1930;
	wire w1931;
	wire w1932;
	wire w1933;
	wire w1934;
	wire w1935;
	wire w1936;
	wire w1937;
	wire w1938;
	wire w1939;
	wire w1940;
	wire w1941;
	wire w1942;
	wire w1943;
	wire w1944;
	wire w1945;
	wire w1946;
	wire w1947;
	wire w1948;
	wire w1949;
	wire w1950;
	wire w1951;
	wire w1952;
	wire w1953;
	wire w1954;
	wire w1955;
	wire w1956;
	wire w1957;
	wire w1958;
	wire w1959;
	wire w1960;
	wire w1961;
	wire w1962;
	wire w1963;
	wire w1964;
	wire w1965;
	wire w1966;
	wire w1967;
	wire w1968;
	wire w1969;
	wire w1970;
	wire w1971;
	wire w1972;
	wire w1973;
	wire w1974;
	wire w1975;
	wire w1976;
	wire w1977;
	wire w1978;
	wire w1979;
	wire w1980;
	wire w1981;
	wire w1982;
	wire w1983;
	wire w1984;
	wire w1985;
	wire w1986;
	wire w1987;
	wire w1988;
	wire w1989;
	wire w1990;
	wire w1991;
	wire w1992;
	wire w1993;
	wire w1994;
	wire w1995;
	wire w1996;
	wire w1997;
	wire w1998;
	wire w1999;
	wire w2000;
	wire w2001;
	wire w2002;
	wire w2003;
	wire w2004;
	wire w2005;
	wire w2006;
	wire w2007;
	wire w2008;
	wire w2009;
	wire w2010;
	wire w2011;
	wire w2012;
	wire w2013;
	wire w2014;
	wire w2015;
	wire w2016;
	wire w2017;
	wire w2018;
	wire w2019;
	wire w2020;
	wire w2021;
	wire w2022;
	wire w2023;
	wire w2024;
	wire w2025;
	wire w2026;
	wire w2027;
	wire w2028;
	wire w2029;
	wire w2030;
	wire w2031;
	wire w2032;
	wire w2033;
	wire w2034;
	wire w2035;
	wire w2036;
	wire w2037;
	wire w2038;
	wire w2039;
	wire w2040;
	wire w2041;
	wire w2042;
	wire w2043;
	wire w2044;
	wire w2045;
	wire w2046;
	wire w2047;
	wire w2048;
	wire w2049;
	wire w2050;
	wire w2051;
	wire w2052;
	wire w2053;
	wire w2054;
	wire w2055;
	wire w2056;
	wire w2057;
	wire w2058;
	wire w2059;
	wire w2060;
	wire w2061;
	wire w2062;
	wire w2063;
	wire w2064;
	wire w2065;
	wire w2066;
	wire w2067;
	wire w2068;
	wire w2069;
	wire w2070;
	wire w2071;
	wire w2072;
	wire w2073;
	wire w2074;
	wire w2075;
	wire w2076;
	wire w2077;
	wire w2078;
	wire w2079;
	wire w2080;
	wire w2081;
	wire w2082;
	wire w2083;
	wire w2084;
	wire w2085;
	wire w2086;
	wire w2087;
	wire w2088;
	wire w2089;
	wire w2090;
	wire w2091;
	wire w2092;
	wire w2093;
	wire w2094;
	wire w2095;
	wire w2096;
	wire w2097;
	wire w2098;
	wire w2099;
	wire w2100;
	wire w2101;
	wire w2102;
	wire w2103;
	wire w2104;
	wire w2105;
	wire w2106;
	wire w2107;
	wire w2108;
	wire w2109;
	wire w2110;
	wire w2111;
	wire w2112;
	wire w2113;
	wire w2114;
	wire w2115;
	wire w2116;
	wire w2117;
	wire w2118;
	wire w2119;
	wire w2120;
	wire w2121;
	wire w2122;
	wire w2123;
	wire w2124;
	wire w2125;
	wire w2126;
	wire w2127;
	wire w2128;
	wire w2129;
	wire w2130;
	wire w2131;
	wire w2132;
	wire w2133;
	wire w2134;
	wire w2135;
	wire w2136;
	wire w2137;
	wire w2138;
	wire w2139;
	wire w2140;
	wire w2141;
	wire w2142;
	wire w2143;
	wire w2144;
	wire w2145;
	wire w2146;
	wire w2147;
	wire w2148;
	wire w2149;
	wire w2150;
	wire w2151;
	wire w2152;
	wire w2153;
	wire w2154;
	wire w2155;
	wire w2156;
	wire w2157;
	wire w2158;
	wire w2159;
	wire w2160;
	wire w2161;
	wire w2162;
	wire w2163;
	wire w2164;
	wire w2165;
	wire w2166;
	wire w2167;
	wire w2168;
	wire w2169;
	wire w2170;
	wire w2171;
	wire w2172;
	wire w2173;
	wire w2174;
	wire w2175;
	wire w2176;
	wire w2177;
	wire w2178;
	wire w2179;
	wire w2180;
	wire w2181;
	wire w2182;
	wire w2183;
	wire w2184;
	wire w2185;
	wire w2186;
	wire w2187;
	wire w2188;
	wire w2189;
	wire w2190;
	wire w2191;
	wire PSG_CLK2;
	wire PSG_CLK1;
	wire w2194;
	wire w2195;
	wire w2196;
	wire w2197;
	wire w2198;
	wire w2199;
	wire w2200;
	wire w2201;
	wire PSG_nCLK2;
	wire PSG_nCLK1;
	wire w2204;
	wire w2205;
	wire w2206;
	wire w2207;
	wire w2208;
	wire w2209;
	wire w2210;
	wire w2211;
	wire w2212;
	wire w2213;
	wire w2214;
	wire w2215;
	wire w2216;
	wire w2217;
	wire w2218;
	wire w2219;
	wire w2220;
	wire w2221;
	wire w2222;
	wire w2223;
	wire w2224;
	wire w2225;
	wire w2226;
	wire w2227;
	wire w2228;
	wire w2229;
	wire w2230;
	wire w2231;
	wire w2232;
	wire w2233;
	wire w2234;
	wire w2235;
	wire w2236;
	wire w2237;
	wire w2238;
	wire w2239;
	wire w2240;
	wire w2241;
	wire w2242;
	wire w2243;
	wire w2244;
	wire w2245;
	wire w2246;
	wire w2247;
	wire w2248;
	wire w2249;
	wire w2250;
	wire w2251;
	wire w2252;
	wire w2253;
	wire w2254;
	wire w2255;
	wire w2256;
	wire w2257;
	wire w2258;
	wire w2259;
	wire w2260;
	wire w2261;
	wire w2262;
	wire w2263;
	wire w2264;
	wire w2265;
	wire w2266;
	wire w2267;
	wire w2268;
	wire w2269;
	wire w2270;
	wire w2271;
	wire w2272;
	wire w2273;
	wire w2274;
	wire w2275;
	wire w2276;
	wire w2277;
	wire w2278;
	wire w2279;
	wire w2280;
	wire w2281;
	wire w2282;
	wire w2283;
	wire w2284;
	wire w2285;
	wire w2286;
	wire w2287;
	wire w2288;
	wire w2289;
	wire w2290;
	wire w2291;
	wire w2292;
	wire w2293;
	wire w2294;
	wire w2295;
	wire w2296;
	wire w2297;
	wire w2298;
	wire w2299;
	wire w2300;
	wire w2301;
	wire w2302;
	wire w2303;
	wire w2304;
	wire w2305;
	wire w2306;
	wire w2307;
	wire w2308;
	wire w2309;
	wire w2310;
	wire w2311;
	wire w2312;
	wire w2313;
	wire w2314;
	wire w2315;
	wire w2316;
	wire w2317;
	wire w2318;
	wire w2319;
	wire w2320;
	wire w2321;
	wire w2322;
	wire w2323;
	wire w2324;
	wire w2325;
	wire w2326;
	wire w2327;
	wire w2328;
	wire w2329;
	wire w2330;
	wire w2331;
	wire w2332;
	wire w2333;
	wire w2334;
	wire w2335;
	wire w2336;
	wire w2337;
	wire w2338;
	wire w2339;
	wire w2340;
	wire w2341;
	wire w2342;
	wire w2343;
	wire w2344;
	wire w2345;
	wire w2346;
	wire w2347;
	wire w2348;
	wire w2349;
	wire w2350;
	wire w2351;
	wire w2352;
	wire w2353;
	wire w2354;
	wire w2355;
	wire w2356;
	wire w2357;
	wire w2358;
	wire w2359;
	wire w2360;
	wire w2361;
	wire w2362;
	wire w2363;
	wire w2364;
	wire w2365;
	wire w2366;
	wire w2367;
	wire w2368;
	wire w2369;
	wire w2370;
	wire w2371;
	wire w2372;
	wire w2373;
	wire w2374;
	wire w2375;
	wire w2376;
	wire w2377;
	wire w2378;
	wire w2379;
	wire w2380;
	wire w2381;
	wire w2382;
	wire w2383;
	wire w2384;
	wire w2385;
	wire w2386;
	wire w2387;
	wire w2388;
	wire w2389;
	wire w2390;
	wire w2391;
	wire w2392;
	wire w2393;
	wire w2394;
	wire w2395;
	wire w2396;
	wire w2397;
	wire w2398;
	wire w2399;
	wire w2400;
	wire w2401;
	wire w2402;
	wire w2403;
	wire w2404;
	wire w2405;
	wire w2406;
	wire w2407;
	wire w2408;
	wire w2409;
	wire w2410;
	wire w2411;
	wire w2412;
	wire w2413;
	wire w2414;
	wire w2415;
	wire w2416;
	wire w2417;
	wire w2418;
	wire w2419;
	wire w2420;
	wire w2421;
	wire w2422;
	wire w2423;
	wire w2424;
	wire w2425;
	wire w2426;
	wire w2427;
	wire w2428;
	wire w2429;
	wire w2430;
	wire w2431;
	wire w2432;
	wire w2433;
	wire w2434;
	wire w2435;
	wire w2436;
	wire w2437;
	wire w2438;
	wire w2439;
	wire w2440;
	wire w2441;
	wire w2442;
	wire w2443;
	wire w2444;
	wire w2445;
	wire w2446;
	wire w2447;
	wire w2448;
	wire w2449;
	wire w2450;
	wire w2451;
	wire w2452;
	wire w2453;
	wire w2454;
	wire w2455;
	wire w2456;
	wire w2457;
	wire w2458;
	wire w2459;
	wire w2460;
	wire w2461;
	wire w2462;
	wire w2463;
	wire w2464;
	wire w2465;
	wire w2466;
	wire w2467;
	wire w2468;
	wire w2469;
	wire w2470;
	wire w2471;
	wire w2472;
	wire w2473;
	wire w2474;
	wire w2475;
	wire w2476;
	wire w2477;
	wire w2478;
	wire w2479;
	wire w2480;
	wire w2481;
	wire w2482;
	wire w2483;
	wire w2484;
	wire w2485;
	wire w2486;
	wire w2487;
	wire w2488;
	wire w2489;
	wire w2490;
	wire w2491;
	wire w2492;
	wire w2493;
	wire w2494;
	wire w2495;
	wire w2496;
	wire w2497;
	wire w2498;
	wire w2499;
	wire w2500;
	wire w2501;
	wire w2502;
	wire w2503;
	wire w2504;
	wire w2505;
	wire w2506;
	wire w2507;
	wire w2508;
	wire w2509;
	wire w2510;
	wire w2511;
	wire w2512;
	wire w2513;
	wire w2514;
	wire w2515;
	wire w2516;
	wire w2517;
	wire w2518;
	wire w2519;
	wire w2520;
	wire w2521;
	wire w2522;
	wire w2523;
	wire w2524;
	wire w2525;
	wire w2526;
	wire w2527;
	wire w2528;
	wire w2529;
	wire w2530;
	wire w2531;
	wire w2532;
	wire w2533;
	wire w2534;
	wire w2535;
	wire w2536;
	wire w2537;
	wire w2538;
	wire w2539;
	wire w2540;
	wire w2541;
	wire w2542;
	wire w2543;
	wire w2544;
	wire w2545;
	wire w2546;
	wire w2547;
	wire w2548;
	wire w2549;
	wire w2550;
	wire w2551;
	wire w2552;
	wire w2553;
	wire w2554;
	wire w2555;
	wire w2556;
	wire w2557;
	wire w2558;
	wire w2559;
	wire w2560;
	wire w2561;
	wire w2562;
	wire w2563;
	wire w2564;
	wire w2565;
	wire w2566;
	wire w2567;
	wire w2568;
	wire w2569;
	wire w2570;
	wire w2571;
	wire w2572;
	wire w2573;
	wire w2574;
	wire w2575;
	wire w2576;
	wire w2577;
	wire w2578;
	wire w2579;
	wire w2580;
	wire w2581;
	wire w2582;
	wire w2583;
	wire w2584;
	wire w2585;
	wire w2586;
	wire w2587;
	wire w2588;
	wire w2589;
	wire w2590;
	wire w2591;
	wire w2592;
	wire w2593;
	wire w2594;
	wire w2595;
	wire w2596;
	wire w2597;
	wire w2598;
	wire w2599;
	wire w2600;
	wire w2601;
	wire w2602;
	wire w2603;
	wire w2604;
	wire w2605;
	wire w2606;
	wire w2607;
	wire w2608;
	wire w2609;
	wire w2610;
	wire w2611;
	wire w2612;
	wire w2613;
	wire w2614;
	wire w2615;
	wire w2616;
	wire w2617;
	wire w2618;
	wire w2619;
	wire w2620;
	wire w2621;
	wire w2622;
	wire w2623;
	wire w2624;
	wire RES;
	wire w2626;
	wire w2627;
	wire w2628;
	wire w2629;
	wire EDCLK_O;
	wire nYS;
	wire w2632;
	wire w2633;
	wire w2634;
	wire w2635;
	wire w2636;
	wire w2637;
	wire w2638;
	wire w2639;
	wire w2640;
	wire w2641;
	wire w2642;
	wire w2643;
	wire w2644;
	wire w2645;
	wire w2646;
	wire w2647;
	wire w2648;
	wire w2649;
	wire w2650;
	wire w2651;
	wire w2652;
	wire w2653;
	wire w2654;
	wire w2655;
	wire w2656;
	wire w2657;
	wire w2658;
	wire w2659;
	wire w2660;
	wire w2661;
	wire w2662;
	wire w2663;
	wire w2664;
	wire w2665;
	wire w2666;
	wire w2667;
	wire w2668;
	wire w2669;
	wire w2670;
	wire w2671;
	wire w2672;
	wire w2673;
	wire w2674;
	wire w2675;
	wire w2676;
	wire w2677;
	wire w2678;
	wire w2679;
	wire w2680;
	wire w2681;
	wire w2682;
	wire w2683;
	wire w2684;
	wire w2685;
	wire w2686;
	wire w2687;
	wire w2688;
	wire w2689;
	wire w2690;
	wire w2691;
	wire w2692;
	wire w2693;
	wire w2694;
	wire w2695;
	wire w2696;
	wire SPR_PRIO;
	wire w2698;
	wire w2699;
	wire w2700;
	wire w2701;
	wire w2702;
	wire w2703;
	wire w2704;
	wire w2705;
	wire w2706;
	wire w2707;
	wire w2708;
	wire w2709;
	wire w2710;
	wire w2711;
	wire w2712;
	wire w2713;
	wire w2714;
	wire w2715;
	wire w2716;
	wire w2717;
	wire w2718;
	wire w2719;
	wire w2720;
	wire w2721;
	wire w2722;
	wire w2723;
	wire w2724;
	wire w2725;
	wire w2726;
	wire w2727;
	wire w2728;
	wire w2729;
	wire w2730;
	wire w2731;
	wire w2732;
	wire w2733;
	wire w2734;
	wire w2735;
	wire w2736;
	wire w2737;
	wire w2738;
	wire w2739;
	wire w2740;
	wire w2741;
	wire w2742;
	wire w2743;
	wire w2744;
	wire w2745;
	wire w2746;
	wire w2747;
	wire w2748;
	wire w2749;
	wire w2750;
	wire w2751;
	wire w2752;
	wire w2753;
	wire w2754;
	wire w2755;
	wire w2756;
	wire w2757;
	wire w2758;
	wire w2759;
	wire w2760;
	wire w2761;
	wire w2762;
	wire w2763;
	wire w2764;
	wire w2765;
	wire PLANE_A_PRIO;
	wire PLANE_B_PRIO;
	wire w2768;
	wire w2769;
	wire w2770;
	wire w2771;
	wire w2772;
	wire w2773;
	wire w2774;
	wire w2775;
	wire w2776;
	wire w2777;
	wire w2778;
	wire w2779;
	wire w2780;
	wire w2781;
	wire w2782;
	wire w2783;
	wire w2784;
	wire w2785;
	wire w2786;
	wire w2787;
	wire w2788;
	wire w2789;
	wire w2790;
	wire w2791;
	wire w2792;
	wire w2793;
	wire w2794;
	wire w2795;
	wire w2796;
	wire w2797;
	wire w2798;
	wire w2799;
	wire w2800;
	wire w2801;
	wire w2802;
	wire w2803;
	wire w2804;
	wire w2805;
	wire w2806;
	wire w2807;
	wire w2808;
	wire w2809;
	wire w2810;
	wire w2811;
	wire w2812;
	wire w2813;
	wire w2814;
	wire w2815;
	wire w2816;
	wire w2817;
	wire w2818;
	wire w2819;
	wire w2820;
	wire w2821;
	wire w2822;
	wire w2823;
	wire w2824;
	wire w2825;
	wire w2826;
	wire w2827;
	wire w2828;
	wire w2829;
	wire w2830;
	wire w2831;
	wire w2832;
	wire w2833;
	wire w2834;
	wire w2835;
	wire w2836;
	wire w2837;
	wire w2838;
	wire w2839;
	wire w2840;
	wire w2841;
	wire w2842;
	wire w2843;
	wire w2844;
	wire w2845;
	wire w2846;
	wire w2847;
	wire w2848;
	wire w2849;
	wire w2850;
	wire w2851;
	wire w2852;
	wire w2853;
	wire w2854;
	wire w2855;
	wire w2856;
	wire w2857;
	wire w2858;
	wire w2859;
	wire w2860;
	wire w2861;
	wire w2862;
	wire w2863;
	wire w2864;
	wire w2865;
	wire w2866;
	wire w2867;
	wire w2868;
	wire w2869;
	wire w2870;
	wire w2871;
	wire w2872;
	wire w2873;
	wire w2874;
	wire w2875;
	wire w2876;
	wire w2877;
	wire w2878;
	wire w2879;
	wire w2880;
	wire w2881;
	wire w2882;
	wire w2883;
	wire w2884;
	wire w2885;
	wire w2886;
	wire w2887;
	wire w2888;
	wire w2889;
	wire w2890;
	wire w2891;
	wire w2892;
	wire w2893;
	wire w2894;
	wire w2895;
	wire w2896;
	wire w2897;
	wire w2898;
	wire w2899;
	wire w2900;
	wire w2901;
	wire w2902;
	wire w2903;
	wire w2904;
	wire w2905;
	wire w2906;
	wire w2907;
	wire w2908;
	wire w2909;
	wire w2910;
	wire w2911;
	wire w2912;
	wire w2913;
	wire w2914;
	wire w2915;
	wire w2916;
	wire w2917;
	wire w2918;
	wire w2919;
	wire w2920;
	wire w2921;
	wire w2922;
	wire w2923;
	wire w2924;
	wire w2925;
	wire w2926;
	wire w2927;
	wire w2928;
	wire w2929;
	wire w2930;
	wire w2931;
	wire w2932;
	wire w2933;
	wire w2934;
	wire w2935;
	wire w2936;
	wire w2937;
	wire w2938;
	wire w2939;
	wire w2940;
	wire w2941;
	wire w2942;
	wire w2943;
	wire w2944;
	wire w2945;
	wire w2946;
	wire w2947;
	wire w2948;
	wire w2949;
	wire w2950;
	wire w2951;
	wire w2952;
	wire w2953;
	wire w2954;
	wire w2955;
	wire w2956;
	wire w2957;
	wire w2958;
	wire w2959;
	wire w2960;
	wire w2961;
	wire w2962;
	wire w2963;
	wire w2964;
	wire w2965;
	wire w2966;
	wire w2967;
	wire w2968;
	wire w2969;
	wire w2970;
	wire w2971;
	wire w2972;
	wire w2973;
	wire w2974;
	wire w2975;
	wire w2976;
	wire w2977;
	wire w2978;
	wire w2979;
	wire w2980;
	wire w2981;
	wire w2982;
	wire w2983;
	wire w2984;
	wire w2985;
	wire w2986;
	wire w2987;
	wire w2988;
	wire w2989;
	wire w2990;
	wire w2991;
	wire w2992;
	wire w2993;
	wire w2994;
	wire w2995;
	wire w2996;
	wire w2997;
	wire w2998;
	wire w2999;
	wire w3000;
	wire w3001;
	wire w3002;
	wire w3003;
	wire w3004;
	wire w3005;
	wire w3006;
	wire w3007;
	wire w3008;
	wire w3009;
	wire w3010;
	wire w3011;
	wire w3012;
	wire w3013;
	wire w3014;
	wire w3015;
	wire w3016;
	wire w3017;
	wire w3018;
	wire w3019;
	wire w3020;
	wire w3021;
	wire w3022;
	wire w3023;
	wire w3024;
	wire w3025;
	wire w3026;
	wire w3027;
	wire w3028;
	wire w3029;
	wire w3030;
	wire w3031;
	wire w3032;
	wire w3033;
	wire w3034;
	wire w3035;
	wire w3036;
	wire w3037;
	wire w3038;
	wire w3039;
	wire w3040;
	wire w3041;
	wire w3042;
	wire w3043;
	wire w3044;
	wire w3045;
	wire w3046;
	wire w3047;
	wire w3048;
	wire w3049;
	wire S[3];
	wire w3051;
	wire w3052;
	wire S[7];
	wire S[2];
	wire w3055;
	wire w3056;
	wire w3057;
	wire w3058;
	wire w3059;
	wire w3060;
	wire S[6];
	wire S[1];
	wire S[5];
	wire S[0];
	wire S[4];
	wire w3066;
	wire w3067;
	wire w3068;
	wire w3069;
	wire w3070;
	wire w3071;
	wire w3072;
	wire w3073;
	wire w3074;
	wire w3075;
	wire w3076;
	wire w3077;
	wire w3078;
	wire w3079;
	wire w3080;
	wire w3081;
	wire w3082;
	wire w3083;
	wire w3084;
	wire w3085;
	wire w3086;
	wire w3087;
	wire w3088;
	wire w3089;
	wire w3090;
	wire w3091;
	wire w3092;
	wire w3093;
	wire w3094;
	wire w3095;
	wire w3096;
	wire w3097;
	wire w3098;
	wire w3099;
	wire w3100;
	wire w3101;
	wire w3102;
	wire w3103;
	wire w3104;
	wire w3105;
	wire w3106;
	wire w3107;
	wire w3108;
	wire w3109;
	wire w3110;
	wire w3111;
	wire w3112;
	wire w3113;
	wire w3114;
	wire w3115;
	wire w3116;
	wire w3117;
	wire w3118;
	wire w3119;
	wire w3120;
	wire w3121;
	wire w3122;
	wire w3123;
	wire w3124;
	wire w3125;
	wire w3126;
	wire w3127;
	wire w3128;
	wire w3129;
	wire w3130;
	wire w3131;
	wire w3132;
	wire w3133;
	wire w3134;
	wire w3135;
	wire w3136;
	wire w3137;
	wire w3138;
	wire w3139;
	wire w3140;
	wire w3141;
	wire w3142;
	wire w3143;
	wire w3144;
	wire w3145;
	wire w3146;
	wire w3147;
	wire w3148;
	wire w3149;
	wire w3150;
	wire w3151;
	wire w3152;
	wire w3153;
	wire w3154;
	wire w3155;
	wire w3156;
	wire w3157;
	wire w3158;
	wire w3159;
	wire w3160;
	wire w3161;
	wire w3162;
	wire w3163;
	wire w3164;
	wire w3165;
	wire w3166;
	wire w3167;
	wire w3168;
	wire w3169;
	wire w3170;
	wire w3171;
	wire w3172;
	wire w3173;
	wire w3174;
	wire w3175;
	wire w3176;
	wire w3177;
	wire w3178;
	wire w3179;
	wire w3180;
	wire w3181;
	wire w3182;
	wire w3183;
	wire w3184;
	wire w3185;
	wire w3186;
	wire w3187;
	wire w3188;
	wire w3189;
	wire w3190;
	wire w3191;
	wire w3192;
	wire w3193;
	wire w3194;
	wire w3195;
	wire w3196;
	wire w3197;
	wire w3198;
	wire w3199;
	wire w3200;
	wire w3201;
	wire w3202;
	wire w3203;
	wire w3204;
	wire w3205;
	wire w3206;
	wire w3207;
	wire w3208;
	wire w3209;
	wire w3210;
	wire w3211;
	wire w3212;
	wire w3213;
	wire w3214;
	wire w3215;
	wire w3216;
	wire w3217;
	wire w3218;
	wire w3219;
	wire w3220;
	wire w3221;
	wire w3222;
	wire w3223;
	wire w3224;
	wire w3225;
	wire w3226;
	wire w3227;
	wire w3228;
	wire w3229;
	wire w3230;
	wire w3231;
	wire w3232;
	wire w3233;
	wire w3234;
	wire w3235;
	wire w3236;
	wire w3237;
	wire w3238;
	wire w3239;
	wire w3240;
	wire w3241;
	wire w3242;
	wire w3243;
	wire w3244;
	wire w3245;
	wire w3246;
	wire w3247;
	wire w3248;
	wire w3249;
	wire w3250;
	wire w3251;
	wire w3252;
	wire w3253;
	wire w3254;
	wire w3255;
	wire w3256;
	wire w3257;
	wire w3258;
	wire w3259;
	wire w3260;
	wire w3261;
	wire w3262;
	wire w3263;
	wire w3264;
	wire w3265;
	wire w3266;
	wire w3267;
	wire w3268;
	wire w3269;
	wire w3270;
	wire w3271;
	wire w3272;
	wire w3273;
	wire w3274;
	wire w3275;
	wire w3276;
	wire w3277;
	wire w3278;
	wire w3279;
	wire w3280;
	wire w3281;
	wire w3282;
	wire w3283;
	wire w3284;
	wire w3285;
	wire w3286;
	wire w3287;
	wire w3288;
	wire w3289;
	wire w3290;
	wire w3291;
	wire w3292;
	wire w3293;
	wire w3294;
	wire w3295;
	wire w3296;
	wire w3297;
	wire w3298;
	wire w3299;
	wire w3300;
	wire w3301;
	wire w3302;
	wire w3303;
	wire w3304;
	wire w3305;
	wire w3306;
	wire w3307;
	wire w3308;
	wire w3309;
	wire w3310;
	wire w3311;
	wire w3312;
	wire w3313;
	wire w3314;
	wire w3315;
	wire w3316;
	wire w3317;
	wire w3318;
	wire w3319;
	wire w3320;
	wire w3321;
	wire w3322;
	wire w3323;
	wire w3324;
	wire w3325;
	wire w3326;
	wire w3327;
	wire w3328;
	wire w3329;
	wire w3330;
	wire w3331;
	wire w3332;
	wire w3333;
	wire w3334;
	wire w3335;
	wire w3336;
	wire w3337;
	wire w3338;
	wire w3339;
	wire w3340;
	wire w3341;
	wire w3342;
	wire w3343;
	wire w3344;
	wire w3345;
	wire w3346;
	wire w3347;
	wire w3348;
	wire w3349;
	wire w3350;
	wire w3351;
	wire w3352;
	wire w3353;
	wire w3354;
	wire w3355;
	wire w3356;
	wire w3357;
	wire w3358;
	wire w3359;
	wire w3360;
	wire w3361;
	wire w3362;
	wire w3363;
	wire w3364;
	wire w3365;
	wire w3366;
	wire w3367;
	wire w3368;
	wire w3369;
	wire w3370;
	wire w3371;
	wire w3372;
	wire w3373;
	wire w3374;
	wire w3375;
	wire w3376;
	wire w3377;
	wire w3378;
	wire w3379;
	wire w3380;
	wire w3381;
	wire w3382;
	wire w3383;
	wire w3384;
	wire w3385;
	wire w3386;
	wire w3387;
	wire w3388;
	wire w3389;
	wire w3390;
	wire w3391;
	wire w3392;
	wire w3393;
	wire w3394;
	wire w3395;
	wire w3396;
	wire w3397;
	wire w3398;
	wire w3399;
	wire w3400;
	wire w3401;
	wire w3402;
	wire w3403;
	wire w3404;
	wire w3405;
	wire w3406;
	wire w3407;
	wire w3408;
	wire w3409;
	wire w3410;
	wire w3411;
	wire w3412;
	wire w3413;
	wire w3414;
	wire w3415;
	wire w3416;
	wire w3417;
	wire w3418;
	wire w3419;
	wire w3420;
	wire w3421;
	wire w3422;
	wire w3423;
	wire w3424;
	wire w3425;
	wire w3426;
	wire w3427;
	wire w3428;
	wire w3429;
	wire w3430;
	wire w3431;
	wire w3432;
	wire w3433;
	wire w3434;
	wire w3435;
	wire w3436;
	wire w3437;
	wire w3438;
	wire w3439;
	wire w3440;
	wire w3441;
	wire w3442;
	wire w3443;
	wire w3444;
	wire w3445;
	wire w3446;
	wire w3447;
	wire w3448;
	wire w3449;
	wire w3450;
	wire w3451;
	wire w3452;
	wire w3453;
	wire w3454;
	wire w3455;
	wire w3456;
	wire w3457;
	wire w3458;
	wire w3459;
	wire w3460;
	wire w3461;
	wire w3462;
	wire w3463;
	wire w3464;
	wire w3465;
	wire w3466;
	wire w3467;
	wire w3468;
	wire w3469;
	wire w3470;
	wire w3471;
	wire w3472;
	wire w3473;
	wire w3474;
	wire w3475;
	wire w3476;
	wire w3477;
	wire w3478;
	wire w3479;
	wire w3480;
	wire w3481;
	wire w3482;
	wire w3483;
	wire w3484;
	wire w3485;
	wire w3486;
	wire w3487;
	wire w3488;
	wire w3489;
	wire w3490;
	wire w3491;
	wire w3492;
	wire w3493;
	wire w3494;
	wire w3495;
	wire w3496;
	wire w3497;
	wire w3498;
	wire w3499;
	wire w3500;
	wire w3501;
	wire w3502;
	wire w3503;
	wire w3504;
	wire w3505;
	wire w3506;
	wire w3507;
	wire w3508;
	wire w3509;
	wire w3510;
	wire w3511;
	wire w3512;
	wire w3513;
	wire w3514;
	wire w3515;
	wire w3516;
	wire w3517;
	wire w3518;
	wire w3519;
	wire w3520;
	wire w3521;
	wire w3522;
	wire w3523;
	wire w3524;
	wire w3525;
	wire w3526;
	wire w3527;
	wire w3528;
	wire w3529;
	wire w3530;
	wire w3531;
	wire w3532;
	wire w3533;
	wire w3534;
	wire w3535;
	wire w3536;
	wire w3537;
	wire w3538;
	wire w3539;
	wire w3540;
	wire w3541;
	wire w3542;
	wire w3543;
	wire w3544;
	wire w3545;
	wire w3546;
	wire w3547;
	wire w3548;
	wire w3549;
	wire w3550;
	wire w3551;
	wire w3552;
	wire w3553;
	wire w3554;
	wire w3555;
	wire w3556;
	wire w3557;
	wire w3558;
	wire w3559;
	wire w3560;
	wire w3561;
	wire w3562;
	wire w3563;
	wire w3564;
	wire w3565;
	wire w3566;
	wire w3567;
	wire w3568;
	wire w3569;
	wire w3570;
	wire w3571;
	wire w3572;
	wire w3573;
	wire w3574;
	wire w3575;
	wire w3576;
	wire w3577;
	wire w3578;
	wire w3579;
	wire w3580;
	wire w3581;
	wire w3582;
	wire w3583;
	wire w3584;
	wire w3585;
	wire w3586;
	wire w3587;
	wire w3588;
	wire w3589;
	wire w3590;
	wire w3591;
	wire w3592;
	wire w3593;
	wire w3594;
	wire w3595;
	wire w3596;
	wire w3597;
	wire w3598;
	wire w3599;
	wire w3600;
	wire w3601;
	wire w3602;
	wire w3603;
	wire w3604;
	wire w3605;
	wire w3606;
	wire w3607;
	wire w3608;
	wire w3609;
	wire w3610;
	wire w3611;
	wire w3612;
	wire w3613;
	wire w3614;
	wire w3615;
	wire w3616;
	wire w3617;
	wire w3618;
	wire w3619;
	wire w3620;
	wire w3621;
	wire w3622;
	wire w3623;
	wire w3624;
	wire w3625;
	wire w3626;
	wire w3627;
	wire w3628;
	wire w3629;
	wire w3630;
	wire w3631;
	wire w3632;
	wire w3633;
	wire w3634;
	wire w3635;
	wire w3636;
	wire w3637;
	wire w3638;
	wire w3639;
	wire w3640;
	wire w3641;
	wire w3642;
	wire w3643;
	wire w3644;
	wire w3645;
	wire w3646;
	wire w3647;
	wire w3648;
	wire w3649;
	wire w3650;
	wire w3651;
	wire w3652;
	wire w3653;
	wire w3654;
	wire w3655;
	wire w3656;
	wire w3657;
	wire w3658;
	wire w3659;
	wire w3660;
	wire w3661;
	wire w3662;
	wire w3663;
	wire w3664;
	wire w3665;
	wire w3666;
	wire w3667;
	wire w3668;
	wire w3669;
	wire w3670;
	wire w3671;
	wire w3672;
	wire w3673;
	wire w3674;
	wire w3675;
	wire w3676;
	wire w3677;
	wire w3678;
	wire w3679;
	wire w3680;
	wire w3681;
	wire w3682;
	wire w3683;
	wire w3684;
	wire w3685;
	wire w3686;
	wire w3687;
	wire w3688;
	wire w3689;
	wire w3690;
	wire w3691;
	wire w3692;
	wire w3693;
	wire w3694;
	wire w3695;
	wire w3696;
	wire w3697;
	wire w3698;
	wire w3699;
	wire w3700;
	wire w3701;
	wire w3702;
	wire w3703;
	wire w3704;
	wire w3705;
	wire w3706;
	wire w3707;
	wire w3708;
	wire w3709;
	wire w3710;
	wire w3711;
	wire w3712;
	wire w3713;
	wire w3714;
	wire w3715;
	wire w3716;
	wire w3717;
	wire w3718;
	wire w3719;
	wire w3720;
	wire w3721;
	wire w3722;
	wire w3723;
	wire w3724;
	wire w3725;
	wire w3726;
	wire w3727;
	wire w3728;
	wire w3729;
	wire w3730;
	wire w3731;
	wire w3732;
	wire w3733;
	wire w3734;
	wire w3735;
	wire w3736;
	wire w3737;
	wire w3738;
	wire w3739;
	wire w3740;
	wire w3741;
	wire w3742;
	wire w3743;
	wire w3744;
	wire w3745;
	wire w3746;
	wire w3747;
	wire w3748;
	wire w3749;
	wire w3750;
	wire w3751;
	wire w3752;
	wire w3753;
	wire w3754;
	wire w3755;
	wire w3756;
	wire w3757;
	wire w3758;
	wire w3759;
	wire w3760;
	wire w3761;
	wire w3762;
	wire w3763;
	wire w3764;
	wire w3765;
	wire w3766;
	wire w3767;
	wire w3768;
	wire w3769;
	wire w3770;
	wire w3771;
	wire w3772;
	wire w3773;
	wire w3774;
	wire w3775;
	wire w3776;
	wire w3777;
	wire w3778;
	wire w3779;
	wire w3780;
	wire w3781;
	wire w3782;
	wire w3783;
	wire w3784;
	wire w3785;
	wire w3786;
	wire w3787;
	wire w3788;
	wire w3789;
	wire w3790;
	wire w3791;
	wire w3792;
	wire w3793;
	wire w3794;
	wire w3795;
	wire w3796;
	wire w3797;
	wire w3798;
	wire w3799;
	wire w3800;
	wire w3801;
	wire w3802;
	wire w3803;
	wire w3804;
	wire w3805;
	wire w3806;
	wire w3807;
	wire w3808;
	wire w3809;
	wire w3810;
	wire w3811;
	wire w3812;
	wire w3813;
	wire w3814;
	wire w3815;
	wire w3816;
	wire w3817;
	wire w3818;
	wire w3819;
	wire w3820;
	wire w3821;
	wire w3822;
	wire w3823;
	wire w3824;
	wire w3825;
	wire w3826;
	wire w3827;
	wire w3828;
	wire w3829;
	wire w3830;
	wire w3831;
	wire w3832;
	wire w3833;
	wire w3834;
	wire w3835;
	wire w3836;
	wire w3837;
	wire w3838;
	wire w3839;
	wire w3840;
	wire w3841;
	wire w3842;
	wire w3843;
	wire w3844;
	wire w3845;
	wire w3846;
	wire w3847;
	wire w3848;
	wire w3849;
	wire w3850;
	wire w3851;
	wire w3852;
	wire w3853;
	wire w3854;
	wire w3855;
	wire w3856;
	wire w3857;
	wire w3858;
	wire w3859;
	wire w3860;
	wire w3861;
	wire w3862;
	wire w3863;
	wire w3864;
	wire w3865;
	wire w3866;
	wire w3867;
	wire w3868;
	wire w3869;
	wire w3870;
	wire w3871;
	wire w3872;
	wire w3873;
	wire w3874;
	wire w3875;
	wire w3876;
	wire w3877;
	wire w3878;
	wire w3879;
	wire w3880;
	wire w3881;
	wire w3882;
	wire w3883;
	wire w3884;
	wire w3885;
	wire w3886;
	wire w3887;
	wire w3888;
	wire w3889;
	wire w3890;
	wire w3891;
	wire w3892;
	wire w3893;
	wire w3894;
	wire w3895;
	wire w3896;
	wire w3897;
	wire w3898;
	wire w3899;
	wire w3900;
	wire w3901;
	wire w3902;
	wire w3903;
	wire w3904;
	wire w3905;
	wire w3906;
	wire w3907;
	wire w3908;
	wire w3909;
	wire w3910;
	wire w3911;
	wire w3912;
	wire w3913;
	wire w3914;
	wire w3915;
	wire w3916;
	wire w3917;
	wire w3918;
	wire w3919;
	wire w3920;
	wire w3921;
	wire w3922;
	wire w3923;
	wire w3924;
	wire w3925;
	wire w3926;
	wire w3927;
	wire w3928;
	wire w3929;
	wire w3930;
	wire w3931;
	wire w3932;
	wire w3933;
	wire w3934;
	wire w3935;
	wire w3936;
	wire w3937;
	wire w3938;
	wire w3939;
	wire w3940;
	wire w3941;
	wire w3942;
	wire w3943;
	wire w3944;
	wire w3945;
	wire w3946;
	wire w3947;
	wire w3948;
	wire w3949;
	wire w3950;
	wire w3951;
	wire w3952;
	wire w3953;
	wire w3954;
	wire w3955;
	wire w3956;
	wire w3957;
	wire w3958;
	wire w3959;
	wire w3960;
	wire w3961;
	wire w3962;
	wire w3963;
	wire w3964;
	wire w3965;
	wire w3966;
	wire w3967;
	wire w3968;
	wire w3969;
	wire w3970;
	wire w3971;
	wire w3972;
	wire w3973;
	wire w3974;
	wire w3975;
	wire w3976;
	wire w3977;
	wire w3978;
	wire w3979;
	wire w3980;
	wire w3981;
	wire w3982;
	wire w3983;
	wire w3984;
	wire w3985;
	wire w3986;
	wire w3987;
	wire w3988;
	wire w3989;
	wire w3990;
	wire w3991;
	wire w3992;
	wire w3993;
	wire w3994;
	wire w3995;
	wire w3996;
	wire w3997;
	wire w3998;
	wire w3999;
	wire w4000;
	wire w4001;
	wire w4002;
	wire w4003;
	wire w4004;
	wire w4005;
	wire w4006;
	wire w4007;
	wire w4008;
	wire w4009;
	wire w4010;
	wire w4011;
	wire w4012;
	wire w4013;
	wire w4014;
	wire w4015;
	wire w4016;
	wire w4017;
	wire w4018;
	wire w4019;
	wire w4020;
	wire w4021;
	wire w4022;
	wire w4023;
	wire w4024;
	wire w4025;
	wire w4026;
	wire w4027;
	wire w4028;
	wire w4029;
	wire w4030;
	wire w4031;
	wire w4032;
	wire w4033;
	wire w4034;
	wire w4035;
	wire w4036;
	wire w4037;
	wire w4038;
	wire w4039;
	wire w4040;
	wire w4041;
	wire w4042;
	wire w4043;
	wire w4044;
	wire w4045;
	wire w4046;
	wire w4047;
	wire w4048;
	wire w4049;
	wire w4050;
	wire w4051;
	wire w4052;
	wire w4053;
	wire w4054;
	wire w4055;
	wire w4056;
	wire w4057;
	wire w4058;
	wire w4059;
	wire w4060;
	wire w4061;
	wire w4062;
	wire w4063;
	wire w4064;
	wire w4065;
	wire w4066;
	wire w4067;
	wire w4068;
	wire w4069;
	wire w4070;
	wire w4071;
	wire w4072;
	wire w4073;
	wire w4074;
	wire w4075;
	wire w4076;
	wire w4077;
	wire w4078;
	wire w4079;
	wire w4080;
	wire w4081;
	wire w4082;
	wire w4083;
	wire w4084;
	wire w4085;
	wire w4086;
	wire w4087;
	wire w4088;
	wire w4089;
	wire w4090;
	wire w4091;
	wire w4092;
	wire w4093;
	wire w4094;
	wire w4095;
	wire w4096;
	wire w4097;
	wire w4098;
	wire w4099;
	wire w4100;
	wire w4101;
	wire w4102;
	wire w4103;
	wire w4104;
	wire w4105;
	wire w4106;
	wire w4107;
	wire w4108;
	wire w4109;
	wire w4110;
	wire w4111;
	wire w4112;
	wire w4113;
	wire w4114;
	wire w4115;
	wire w4116;
	wire w4117;
	wire w4118;
	wire w4119;
	wire w4120;
	wire w4121;
	wire w4122;
	wire w4123;
	wire w4124;
	wire w4125;
	wire w4126;
	wire w4127;
	wire w4128;
	wire w4129;
	wire w4130;
	wire w4131;
	wire w4132;
	wire w4133;
	wire w4134;
	wire w4135;
	wire w4136;
	wire w4137;
	wire w4138;
	wire w4139;
	wire w4140;
	wire w4141;
	wire w4142;
	wire w4143;
	wire w4144;
	wire w4145;
	wire w4146;
	wire w4147;
	wire w4148;
	wire w4149;
	wire w4150;
	wire w4151;
	wire w4152;
	wire w4153;
	wire w4154;
	wire w4155;
	wire w4156;
	wire w4157;
	wire w4158;
	wire w4159;
	wire w4160;
	wire w4161;
	wire w4162;
	wire w4163;
	wire w4164;
	wire w4165;
	wire w4166;
	wire w4167;
	wire w4168;
	wire w4169;
	wire w4170;
	wire w4171;
	wire w4172;
	wire w4173;
	wire w4174;
	wire w4175;
	wire w4176;
	wire w4177;
	wire w4178;
	wire w4179;
	wire w4180;
	wire w4181;
	wire w4182;
	wire w4183;
	wire w4184;
	wire w4185;
	wire w4186;
	wire w4187;
	wire w4188;
	wire w4189;
	wire w4190;
	wire w4191;
	wire w4192;
	wire w4193;
	wire w4194;
	wire w4195;
	wire w4196;
	wire w4197;
	wire w4198;
	wire w4199;
	wire w4200;
	wire w4201;
	wire w4202;
	wire w4203;
	wire w4204;
	wire w4205;
	wire w4206;
	wire w4207;
	wire w4208;
	wire w4209;
	wire w4210;
	wire w4211;
	wire w4212;
	wire w4213;
	wire w4214;
	wire w4215;
	wire w4216;
	wire w4217;
	wire w4218;
	wire w4219;
	wire w4220;
	wire w4221;
	wire w4222;
	wire w4223;
	wire w4224;
	wire w4225;
	wire w4226;
	wire w4227;
	wire w4228;
	wire w4229;
	wire w4230;
	wire w4231;
	wire w4232;
	wire w4233;
	wire w4234;
	wire w4235;
	wire w4236;
	wire w4237;
	wire w4238;
	wire w4239;
	wire w4240;
	wire w4241;
	wire w4242;
	wire w4243;
	wire w4244;
	wire w4245;
	wire w4246;
	wire w4247;
	wire w4248;
	wire w4249;
	wire w4250;
	wire w4251;
	wire w4252;
	wire w4253;
	wire w4254;
	wire w4255;
	wire w4256;
	wire w4257;
	wire w4258;
	wire w4259;
	wire w4260;
	wire w4261;
	wire w4262;
	wire w4263;
	wire w4264;
	wire w4265;
	wire w4266;
	wire w4267;
	wire w4268;
	wire w4269;
	wire w4270;
	wire w4271;
	wire w4272;
	wire w4273;
	wire w4274;
	wire w4275;
	wire w4276;
	wire w4277;
	wire w4278;
	wire w4279;
	wire w4280;
	wire w4281;
	wire w4282;
	wire w4283;
	wire w4284;
	wire w4285;
	wire w4286;
	wire w4287;
	wire w4288;
	wire w4289;
	wire w4290;
	wire w4291;
	wire w4292;
	wire w4293;
	wire w4294;
	wire w4295;
	wire w4296;
	wire w4297;
	wire w4298;
	wire w4299;
	wire w4300;
	wire w4301;
	wire w4302;
	wire w4303;
	wire w4304;
	wire w4305;
	wire w4306;
	wire w4307;
	wire w4308;
	wire w4309;
	wire w4310;
	wire w4311;
	wire w4312;
	wire w4313;
	wire w4314;
	wire w4315;
	wire w4316;
	wire w4317;
	wire w4318;
	wire w4319;
	wire w4320;
	wire w4321;
	wire w4322;
	wire w4323;
	wire w4324;
	wire w4325;
	wire w4326;
	wire w4327;
	wire w4328;
	wire w4329;
	wire w4330;
	wire w4331;
	wire w4332;
	wire w4333;
	wire w4334;
	wire w4335;
	wire w4336;
	wire w4337;
	wire w4338;
	wire w4339;
	wire w4340;
	wire w4341;
	wire w4342;
	wire w4343;
	wire w4344;
	wire w4345;
	wire w4346;
	wire w4347;
	wire w4348;
	wire w4349;
	wire w4350;
	wire w4351;
	wire w4352;
	wire w4353;
	wire w4354;
	wire w4355;
	wire w4356;
	wire w4357;
	wire w4358;
	wire w4359;
	wire w4360;
	wire w4361;
	wire w4362;
	wire w4363;
	wire w4364;
	wire w4365;
	wire w4366;
	wire w4367;
	wire w4368;
	wire w4369;
	wire w4370;
	wire w4371;
	wire w4372;
	wire w4373;
	wire w4374;
	wire w4375;
	wire w4376;
	wire w4377;
	wire w4378;
	wire w4379;
	wire w4380;
	wire w4381;
	wire w4382;
	wire w4383;
	wire w4384;
	wire w4385;
	wire w4386;
	wire w4387;
	wire w4388;
	wire w4389;
	wire w4390;
	wire w4391;
	wire w4392;
	wire w4393;
	wire w4394;
	wire w4395;
	wire w4396;
	wire w4397;
	wire w4398;
	wire w4399;
	wire w4400;
	wire w4401;
	wire w4402;
	wire w4403;
	wire w4404;
	wire w4405;
	wire w4406;
	wire w4407;
	wire w4408;
	wire w4409;
	wire w4410;
	wire w4411;
	wire w4412;
	wire w4413;
	wire w4414;
	wire w4415;
	wire w4416;
	wire w4417;
	wire w4418;
	wire w4419;
	wire w4420;
	wire w4421;
	wire w4422;
	wire w4423;
	wire w4424;
	wire w4425;
	wire w4426;
	wire w4427;
	wire w4428;
	wire w4429;
	wire w4430;
	wire w4431;
	wire w4432;
	wire w4433;
	wire w4434;
	wire w4435;
	wire w4436;
	wire w4437;
	wire w4438;
	wire w4439;
	wire w4440;
	wire w4441;
	wire w4442;
	wire w4443;
	wire 68K CPU CLOCK;
	wire w4445;
	wire w4446;
	wire w4447;
	wire w4448;
	wire w4449;
	wire w4450;
	wire w4451;
	wire w4452;
	wire w4453;
	wire w4454;
	wire w4455;
	wire w4456;
	wire w4457;
	wire w4458;
	wire w4459;
	wire w4460;
	wire w4461;
	wire w4462;
	wire w4463;
	wire w4464;
	wire w4465;
	wire w4466;
	wire w4467;
	wire w4468;
	wire w4469;
	wire w4470;
	wire w4471;
	wire w4472;
	wire w4473;
	wire w4474;
	wire w4475;
	wire w4476;
	wire w4477;
	wire w4478;
	wire w4479;
	wire w4480;
	wire w4481;
	wire w4482;
	wire w4483;
	wire w4484;
	wire w4485;
	wire w4486;
	wire w4487;
	wire w4488;
	wire nRAS1;
	wire nCAS1;
	wire nWE1;
	wire nWE0;
	wire nOE1;
	wire AD_RD_DIR;
	wire w4495;
	wire w4496;
	wire w4497;
	wire w4498;
	wire w4499;
	wire w4500;
	wire w4501;
	wire w4502;
	wire w4503;
	wire w4504;
	wire w4505;
	wire w4506;
	wire w4507;
	wire w4508;
	wire w4509;
	wire w4510;
	wire w4511;
	wire w4512;
	wire w4513;
	wire w4514;
	wire w4515;
	wire w4516;
	wire w4517;
	wire w4518;
	wire w4519;
	wire w4520;
	wire w4521;
	wire w4522;
	wire w4523;
	wire w4524;
	wire w4525;
	wire w4526;
	wire w4527;
	wire w4528;
	wire w4529;
	wire w4530;
	wire w4531;
	wire w4532;
	wire w4533;
	wire w4534;
	wire w4535;
	wire w4536;
	wire w4537;
	wire w4538;
	wire w4539;
	wire w4540;
	wire w4541;
	wire w4542;
	wire w4543;
	wire w4544;
	wire w4545;
	wire w4546;
	wire w4547;
	wire w4548;
	wire w4549;
	wire w4550;
	wire w4551;
	wire w4552;
	wire w4553;
	wire w4554;
	wire w4555;
	wire w4556;
	wire w4557;
	wire w4558;
	wire w4559;
	wire w4560;
	wire w4561;
	wire w4562;
	wire w4563;
	wire w4564;
	wire w4565;
	wire w4566;
	wire w4567;
	wire w4568;
	wire w4569;
	wire w4570;
	wire w4571;
	wire w4572;
	wire w4573;
	wire w4574;
	wire w4575;
	wire w4576;
	wire w4577;
	wire w4578;
	wire w4579;
	wire w4580;
	wire w4581;
	wire w4582;
	wire w4583;
	wire w4584;
	wire w4585;
	wire w4586;
	wire w4587;
	wire w4588;
	wire w4589;
	wire w4590;
	wire w4591;
	wire w4592;
	wire w4593;
	wire w4594;
	wire w4595;
	wire w4596;
	wire w4597;
	wire w4598;
	wire w4599;
	wire w4600;
	wire w4601;
	wire w4602;
	wire w4603;
	wire w4604;
	wire w4605;
	wire w4606;
	wire w4607;
	wire w4608;
	wire w4609;
	wire w4610;
	wire w4611;
	wire w4612;
	wire w4613;
	wire w4614;
	wire w4615;
	wire w4616;
	wire w4617;
	wire w4618;
	wire w4619;
	wire w4620;
	wire w4621;
	wire w4622;
	wire w4623;
	wire w4624;
	wire w4625;
	wire w4626;
	wire w4627;
	wire w4628;
	wire w4629;
	wire w4630;
	wire w4631;
	wire w4632;
	wire w4633;
	wire w4634;
	wire w4635;
	wire w4636;
	wire w4637;
	wire w4638;
	wire w4639;
	wire w4640;
	wire w4641;
	wire w4642;
	wire w4643;
	wire w4644;
	wire w4645;
	wire w4646;
	wire w4647;
	wire w4648;
	wire w4649;
	wire w4650;
	wire w4651;
	wire w4652;
	wire w4653;
	wire w4654;
	wire w4655;
	wire w4656;
	wire w4657;
	wire w4658;
	wire w4659;
	wire w4660;
	wire w4661;
	wire w4662;
	wire w4663;
	wire w4664;
	wire w4665;
	wire w4666;
	wire w4667;
	wire w4668;
	wire w4669;
	wire w4670;
	wire w4671;
	wire w4672;
	wire w4673;
	wire w4674;
	wire w4675;
	wire w4676;
	wire w4677;
	wire w4678;
	wire w4679;
	wire w4680;
	wire w4681;
	wire w4682;
	wire w4683;
	wire w4684;
	wire w4685;
	wire w4686;
	wire w4687;
	wire w4688;
	wire w4689;
	wire w4690;
	wire w4691;
	wire w4692;
	wire w4693;
	wire w4694;
	wire w4695;
	wire w4696;
	wire w4697;
	wire w4698;
	wire w4699;
	wire w4700;
	wire w4701;
	wire w4702;
	wire w4703;
	wire w4704;
	wire w4705;
	wire w4706;
	wire w4707;
	wire w4708;
	wire w4709;
	wire w4710;
	wire w4711;
	wire w4712;
	wire w4713;
	wire w4714;
	wire w4715;
	wire w4716;
	wire w4717;
	wire w4718;
	wire w4719;
	wire w4720;
	wire w4721;
	wire w4722;
	wire w4723;
	wire w4724;
	wire w4725;
	wire w4726;
	wire w4727;
	wire w4728;
	wire w4729;
	wire w4730;
	wire w4731;
	wire w4732;
	wire w4733;
	wire w4734;
	wire w4735;
	wire w4736;
	wire w4737;
	wire w4738;
	wire w4739;
	wire w4740;
	wire w4741;
	wire w4742;
	wire w4743;
	wire w4744;
	wire w4745;
	wire w4746;
	wire w4747;
	wire w4748;
	wire w4749;
	wire w4750;
	wire w4751;
	wire w4752;
	wire w4753;
	wire w4754;
	wire w4755;
	wire w4756;
	wire w4757;
	wire w4758;
	wire w4759;
	wire w4760;
	wire w4761;
	wire w4762;
	wire w4763;
	wire w4764;
	wire w4765;
	wire w4766;
	wire w4767;
	wire w4768;
	wire w4769;
	wire w4770;
	wire w4771;
	wire w4772;
	wire w4773;
	wire w4774;
	wire w4775;
	wire w4776;
	wire w4777;
	wire w4778;
	wire w4779;
	wire w4780;
	wire w4781;
	wire w4782;
	wire w4783;
	wire w4784;
	wire w4785;
	wire w4786;
	wire w4787;
	wire w4788;
	wire w4789;
	wire w4790;
	wire w4791;
	wire w4792;
	wire w4793;
	wire w4794;
	wire w4795;
	wire w4796;
	wire w4797;
	wire w4798;
	wire w4799;
	wire w4800;
	wire w4801;
	wire w4802;
	wire w4803;
	wire w4804;
	wire w4805;
	wire w4806;
	wire w4807;
	wire w4808;
	wire w4809;
	wire w4810;
	wire w4811;
	wire w4812;
	wire w4813;
	wire w4814;
	wire w4815;
	wire w4816;
	wire w4817;
	wire w4818;
	wire w4819;
	wire w4820;
	wire w4821;
	wire w4822;
	wire w4823;
	wire w4824;
	wire w4825;
	wire w4826;
	wire w4827;
	wire w4828;
	wire w4829;
	wire w4830;
	wire w4831;
	wire w4832;
	wire w4833;
	wire w4834;
	wire w4835;
	wire w4836;
	wire w4837;
	wire w4838;
	wire w4839;
	wire w4840;
	wire w4841;
	wire w4842;
	wire w4843;
	wire w4844;
	wire w4845;
	wire w4846;
	wire w4847;
	wire w4848;
	wire w4849;
	wire w4850;
	wire w4851;
	wire w4852;
	wire w4853;
	wire w4854;
	wire w4855;
	wire w4856;
	wire w4857;
	wire w4858;
	wire w4859;
	wire w4860;
	wire w4861;
	wire w4862;
	wire w4863;
	wire w4864;
	wire w4865;
	wire w4866;
	wire w4867;
	wire w4868;
	wire w4869;
	wire w4870;
	wire w4871;
	wire w4872;
	wire w4873;
	wire w4874;
	wire w4875;
	wire w4876;
	wire w4877;
	wire w4878;
	wire w4879;
	wire w4880;
	wire w4881;
	wire w4882;
	wire w4883;
	wire w4884;
	wire w4885;
	wire w4886;
	wire w4887;
	wire w4888;
	wire w4889;
	wire w4890;
	wire w4891;
	wire w4892;
	wire w4893;
	wire w4894;
	wire w4895;
	wire w4896;
	wire w4897;
	wire w4898;
	wire w4899;
	wire w4900;
	wire w4901;
	wire w4902;
	wire w4903;
	wire w4904;
	wire w4905;
	wire w4906;
	wire w4907;
	wire w4908;
	wire w4909;
	wire w4910;
	wire w4911;
	wire w4912;
	wire w4913;
	wire w4914;
	wire w4915;
	wire w4916;
	wire w4917;
	wire w4918;
	wire w4919;
	wire w4920;
	wire w4921;
	wire w4922;
	wire w4923;
	wire w4924;
	wire w4925;
	wire w4926;
	wire w4927;
	wire w4928;
	wire w4929;
	wire w4930;
	wire w4931;
	wire w4932;
	wire w4933;
	wire w4934;
	wire w4935;
	wire w4936;
	wire w4937;
	wire w4938;
	wire w4939;
	wire w4940;
	wire w4941;
	wire w4942;
	wire w4943;
	wire w4944;
	wire w4945;
	wire w4946;
	wire w4947;
	wire w4948;
	wire w4949;
	wire w4950;
	wire w4951;
	wire w4952;
	wire w4953;
	wire w4954;
	wire w4955;
	wire w4956;
	wire w4957;
	wire w4958;
	wire w4959;
	wire w4960;
	wire w4961;
	wire w4962;
	wire w4963;
	wire w4964;
	wire w4965;
	wire w4966;
	wire w4967;
	wire w4968;
	wire w4969;
	wire w4970;
	wire w4971;
	wire w4972;
	wire w4973;
	wire w4974;
	wire w4975;
	wire w4976;
	wire w4977;
	wire w4978;
	wire w4979;
	wire w4980;
	wire w4981;
	wire w4982;
	wire w4983;
	wire w4984;
	wire w4985;
	wire w4986;
	wire w4987;
	wire w4988;
	wire w4989;
	wire w4990;
	wire w4991;
	wire w4992;
	wire w4993;
	wire w4994;
	wire w4995;
	wire w4996;
	wire w4997;
	wire w4998;
	wire w4999;
	wire w5000;
	wire w5001;
	wire w5002;
	wire w5003;
	wire w5004;
	wire w5005;
	wire w5006;
	wire w5007;
	wire w5008;
	wire w5009;
	wire w5010;
	wire w5011;
	wire w5012;
	wire w5013;
	wire w5014;
	wire w5015;
	wire w5016;
	wire w5017;
	wire w5018;
	wire w5019;
	wire w5020;
	wire w5021;
	wire w5022;
	wire w5023;
	wire w5024;
	wire w5025;
	wire w5026;
	wire w5027;
	wire w5028;
	wire w5029;
	wire w5030;
	wire w5031;
	wire w5032;
	wire w5033;
	wire w5034;
	wire w5035;
	wire w5036;
	wire w5037;
	wire w5038;
	wire w5039;
	wire w5040;
	wire w5041;
	wire w5042;
	wire w5043;
	wire w5044;
	wire w5045;
	wire w5046;
	wire w5047;
	wire w5048;
	wire w5049;
	wire w5050;
	wire w5051;
	wire w5052;
	wire w5053;
	wire w5054;
	wire w5055;
	wire w5056;
	wire w5057;
	wire w5058;
	wire w5059;
	wire w5060;
	wire w5061;
	wire w5062;
	wire w5063;
	wire w5064;
	wire w5065;
	wire w5066;
	wire w5067;
	wire w5068;
	wire w5069;
	wire w5070;
	wire w5071;
	wire w5072;
	wire w5073;
	wire w5074;
	wire w5075;
	wire w5076;
	wire w5077;
	wire w5078;
	wire w5079;
	wire w5080;
	wire w5081;
	wire w5082;
	wire w5083;
	wire w5084;
	wire w5085;
	wire w5086;
	wire w5087;
	wire w5088;
	wire w5089;
	wire w5090;
	wire w5091;
	wire w5092;
	wire w5093;
	wire w5094;
	wire w5095;
	wire w5096;
	wire w5097;
	wire w5098;
	wire w5099;
	wire w5100;
	wire w5101;
	wire w5102;
	wire w5103;
	wire w5104;
	wire w5105;
	wire w5106;
	wire w5107;
	wire w5108;
	wire w5109;
	wire w5110;
	wire w5111;
	wire w5112;
	wire w5113;
	wire w5114;
	wire w5115;
	wire w5116;
	wire w5117;
	wire w5118;
	wire w5119;
	wire w5120;
	wire w5121;
	wire w5122;
	wire w5123;
	wire w5124;
	wire w5125;
	wire w5126;
	wire w5127;
	wire w5128;
	wire w5129;
	wire w5130;
	wire w5131;
	wire w5132;
	wire w5133;
	wire w5134;
	wire w5135;
	wire w5136;
	wire w5137;
	wire w5138;
	wire w5139;
	wire w5140;
	wire w5141;
	wire w5142;
	wire w5143;
	wire w5144;
	wire w5145;
	wire w5146;
	wire w5147;
	wire w5148;
	wire w5149;
	wire w5150;
	wire w5151;
	wire w5152;
	wire w5153;
	wire w5154;
	wire w5155;
	wire w5156;
	wire w5157;
	wire w5158;
	wire w5159;
	wire w5160;
	wire w5161;
	wire w5162;
	wire w5163;
	wire w5164;
	wire w5165;
	wire w5166;
	wire w5167;
	wire w5168;
	wire w5169;
	wire w5170;
	wire w5171;
	wire w5172;
	wire w5173;
	wire w5174;
	wire w5175;
	wire w5176;
	wire w5177;
	wire w5178;
	wire w5179;
	wire w5180;
	wire w5181;
	wire w5182;
	wire w5183;
	wire w5184;
	wire w5185;
	wire w5186;
	wire w5187;
	wire w5188;
	wire w5189;
	wire w5190;
	wire w5191;
	wire w5192;
	wire w5193;
	wire w5194;
	wire w5195;
	wire w5196;
	wire w5197;
	wire w5198;
	wire w5199;
	wire w5200;
	wire w5201;
	wire w5202;
	wire w5203;
	wire w5204;
	wire w5205;
	wire w5206;
	wire w5207;
	wire w5208;
	wire w5209;
	wire w5210;
	wire w5211;
	wire w5212;
	wire w5213;
	wire w5214;
	wire w5215;
	wire w5216;
	wire w5217;
	wire w5218;
	wire w5219;
	wire w5220;
	wire w5221;
	wire w5222;
	wire w5223;
	wire w5224;
	wire w5225;
	wire w5226;
	wire w5227;
	wire w5228;
	wire w5229;
	wire w5230;
	wire w5231;
	wire w5232;
	wire w5233;
	wire w5234;
	wire w5235;
	wire w5236;
	wire w5237;
	wire w5238;
	wire w5239;
	wire w5240;
	wire w5241;
	wire w5242;
	wire w5243;
	wire w5244;
	wire w5245;
	wire w5246;
	wire w5247;
	wire w5248;
	wire w5249;
	wire w5250;
	wire w5251;
	wire w5252;
	wire w5253;
	wire w5254;
	wire w5255;
	wire w5256;
	wire w5257;
	wire w5258;
	wire w5259;
	wire w5260;
	wire w5261;
	wire w5262;
	wire w5263;
	wire w5264;
	wire w5265;
	wire w5266;
	wire w5267;
	wire w5268;
	wire w5269;
	wire w5270;
	wire w5271;
	wire w5272;
	wire w5273;
	wire w5274;
	wire w5275;
	wire w5276;
	wire w5277;
	wire w5278;
	wire w5279;
	wire w5280;
	wire w5281;
	wire w5282;
	wire w5283;
	wire w5284;
	wire w5285;
	wire w5286;
	wire w5287;
	wire w5288;
	wire w5289;
	wire w5290;
	wire w5291;
	wire w5292;
	wire w5293;
	wire w5294;
	wire w5295;
	wire w5296;
	wire w5297;
	wire w5298;
	wire w5299;
	wire w5300;
	wire w5301;
	wire w5302;
	wire w5303;
	wire w5304;
	wire w5305;
	wire w5306;
	wire w5307;
	wire w5308;
	wire w5309;
	wire w5310;
	wire w5311;
	wire w5312;
	wire w5313;
	wire w5314;
	wire w5315;
	wire w5316;
	wire w5317;
	wire w5318;
	wire w5319;
	wire w5320;
	wire w5321;
	wire w5322;
	wire w5323;
	wire w5324;
	wire w5325;
	wire w5326;
	wire w5327;
	wire w5328;
	wire w5329;
	wire w5330;
	wire w5331;
	wire w5332;
	wire w5333;
	wire w5334;
	wire w5335;
	wire w5336;
	wire w5337;
	wire w5338;
	wire w5339;
	wire w5340;
	wire w5341;
	wire w5342;
	wire w5343;
	wire w5344;
	wire w5345;
	wire w5346;
	wire w5347;
	wire w5348;
	wire w5349;
	wire w5350;
	wire w5351;
	wire w5352;
	wire w5353;
	wire w5354;
	wire w5355;
	wire w5356;
	wire w5357;
	wire w5358;
	wire w5359;
	wire w5360;
	wire w5361;
	wire w5362;
	wire w5363;
	wire w5364;
	wire w5365;
	wire w5366;
	wire w5367;
	wire w5368;
	wire w5369;
	wire w5370;
	wire w5371;
	wire w5372;
	wire w5373;
	wire w5374;
	wire w5375;
	wire w5376;
	wire w5377;
	wire w5378;
	wire w5379;
	wire w5380;
	wire w5381;
	wire w5382;
	wire w5383;
	wire w5384;
	wire w5385;
	wire w5386;
	wire w5387;
	wire w5388;
	wire w5389;
	wire w5390;
	wire w5391;
	wire w5392;
	wire w5393;
	wire w5394;
	wire w5395;
	wire w5396;
	wire w5397;
	wire w5398;
	wire w5399;
	wire w5400;
	wire w5401;
	wire w5402;
	wire w5403;
	wire w5404;
	wire w5405;
	wire w5406;
	wire w5407;
	wire w5408;
	wire w5409;
	wire w5410;
	wire w5411;
	wire w5412;
	wire w5413;
	wire w5414;
	wire w5415;
	wire w5416;
	wire w5417;
	wire w5418;
	wire w5419;
	wire w5420;
	wire w5421;
	wire w5422;
	wire w5423;
	wire w5424;
	wire w5425;
	wire w5426;
	wire w5427;
	wire w5428;
	wire w5429;
	wire w5430;
	wire w5431;
	wire w5432;
	wire w5433;
	wire w5434;
	wire w5435;
	wire w5436;
	wire w5437;
	wire w5438;
	wire w5439;
	wire w5440;
	wire w5441;
	wire w5442;
	wire w5443;
	wire w5444;
	wire w5445;
	wire w5446;
	wire w5447;
	wire w5448;
	wire w5449;
	wire w5450;
	wire w5451;
	wire w5452;
	wire w5453;
	wire w5454;
	wire w5455;
	wire w5456;
	wire w5457;
	wire w5458;
	wire w5459;
	wire w5460;
	wire w5461;
	wire w5462;
	wire w5463;
	wire w5464;
	wire w5465;
	wire w5466;
	wire w5467;
	wire w5468;
	wire w5469;
	wire w5470;
	wire w5471;
	wire w5472;
	wire w5473;
	wire w5474;
	wire w5475;
	wire w5476;
	wire w5477;
	wire w5478;
	wire w5479;
	wire w5480;
	wire w5481;
	wire w5482;
	wire w5483;
	wire w5484;
	wire w5485;
	wire w5486;
	wire w5487;
	wire w5488;
	wire w5489;
	wire w5490;
	wire w5491;
	wire w5492;
	wire w5493;
	wire w5494;
	wire w5495;
	wire w5496;
	wire w5497;
	wire w5498;
	wire w5499;
	wire w5500;
	wire w5501;
	wire w5502;
	wire w5503;
	wire w5504;
	wire w5505;
	wire w5506;
	wire w5507;
	wire w5508;
	wire w5509;
	wire w5510;
	wire w5511;
	wire w5512;
	wire w5513;
	wire w5514;
	wire w5515;
	wire w5516;
	wire w5517;
	wire w5518;
	wire w5519;
	wire w5520;
	wire w5521;
	wire w5522;
	wire w5523;
	wire w5524;
	wire w5525;
	wire w5526;
	wire w5527;
	wire w5528;
	wire w5529;
	wire w5530;
	wire w5531;
	wire w5532;
	wire w5533;
	wire w5534;
	wire w5535;
	wire w5536;
	wire w5537;
	wire w5538;
	wire w5539;
	wire w5540;
	wire w5541;
	wire w5542;
	wire w5543;
	wire w5544;
	wire w5545;
	wire w5546;
	wire w5547;
	wire w5548;
	wire w5549;
	wire w5550;
	wire w5551;
	wire w5552;
	wire w5553;
	wire w5554;
	wire w5555;
	wire w5556;
	wire w5557;
	wire w5558;
	wire w5559;
	wire w5560;
	wire w5561;
	wire w5562;
	wire w5563;
	wire w5564;
	wire w5565;
	wire w5566;
	wire w5567;
	wire w5568;
	wire w5569;
	wire w5570;
	wire w5571;
	wire w5572;
	wire w5573;
	wire w5574;
	wire w5575;
	wire w5576;
	wire w5577;
	wire w5578;
	wire w5579;
	wire w5580;
	wire w5581;
	wire w5582;
	wire w5583;
	wire w5584;
	wire w5585;
	wire w5586;
	wire w5587;
	wire w5588;
	wire w5589;
	wire w5590;
	wire w5591;
	wire w5592;
	wire w5593;
	wire w5594;
	wire w5595;
	wire w5596;
	wire w5597;
	wire w5598;
	wire w5599;
	wire w5600;
	wire w5601;
	wire w5602;
	wire w5603;
	wire w5604;
	wire w5605;
	wire w5606;
	wire w5607;
	wire w5608;
	wire w5609;
	wire w5610;
	wire w5611;
	wire w5612;
	wire w5613;
	wire w5614;
	wire w5615;
	wire w5616;
	wire w5617;
	wire w5618;
	wire w5619;
	wire w5620;
	wire w5621;
	wire w5622;
	wire w5623;
	wire w5624;
	wire w5625;
	wire w5626;
	wire w5627;
	wire w5628;
	wire w5629;
	wire w5630;
	wire w5631;
	wire w5632;
	wire w5633;
	wire w5634;
	wire w5635;
	wire w5636;
	wire w5637;
	wire w5638;
	wire w5639;
	wire w5640;
	wire w5641;
	wire w5642;
	wire w5643;
	wire w5644;
	wire w5645;
	wire w5646;
	wire w5647;
	wire w5648;
	wire w5649;
	wire w5650;
	wire w5651;
	wire w5652;
	wire w5653;
	wire w5654;
	wire w5655;
	wire w5656;
	wire w5657;
	wire w5658;
	wire w5659;
	wire w5660;
	wire w5661;
	wire w5662;
	wire w5663;
	wire w5664;
	wire w5665;
	wire w5666;
	wire w5667;
	wire w5668;
	wire w5669;
	wire w5670;
	wire w5671;
	wire w5672;
	wire w5673;
	wire w5674;
	wire w5675;
	wire w5676;
	wire w5677;
	wire w5678;
	wire w5679;
	wire w5680;
	wire w5681;
	wire w5682;
	wire w5683;
	wire w5684;
	wire w5685;
	wire w5686;
	wire w5687;
	wire w5688;
	wire w5689;
	wire w5690;
	wire w5691;
	wire w5692;
	wire w5693;
	wire w5694;
	wire w5695;
	wire w5696;
	wire w5697;
	wire w5698;
	wire w5699;
	wire w5700;
	wire w5701;
	wire w5702;
	wire w5703;
	wire w5704;
	wire w5705;
	wire w5706;
	wire w5707;
	wire w5708;
	wire w5709;
	wire w5710;
	wire w5711;
	wire w5712;
	wire w5713;
	wire w5714;
	wire w5715;
	wire w5716;
	wire w5717;
	wire w5718;
	wire w5719;
	wire w5720;
	wire w5721;
	wire w5722;
	wire w5723;
	wire w5724;
	wire w5725;
	wire w5726;
	wire w5727;
	wire w5728;
	wire w5729;
	wire w5730;
	wire w5731;
	wire w5732;
	wire w5733;
	wire w5734;
	wire w5735;
	wire w5736;
	wire w5737;
	wire w5738;
	wire w5739;
	wire w5740;
	wire w5741;
	wire w5742;
	wire w5743;
	wire w5744;
	wire w5745;
	wire w5746;
	wire w5747;
	wire w5748;
	wire w5749;
	wire w5750;
	wire w5751;
	wire w5752;
	wire w5753;
	wire w5754;
	wire w5755;
	wire w5756;
	wire w5757;
	wire w5758;
	wire w5759;
	wire w5760;
	wire w5761;
	wire w5762;
	wire w5763;
	wire w5764;
	wire w5765;
	wire w5766;
	wire w5767;
	wire w5768;
	wire w5769;
	wire w5770;
	wire w5771;
	wire w5772;
	wire w5773;
	wire w5774;
	wire w5775;
	wire w5776;
	wire w5777;
	wire w5778;
	wire w5779;
	wire w5780;
	wire w5781;
	wire w5782;
	wire w5783;
	wire w5784;
	wire w5785;
	wire w5786;
	wire w5787;
	wire w5788;
	wire w5789;
	wire w5790;
	wire w5791;
	wire w5792;
	wire w5793;
	wire w5794;
	wire w5795;
	wire w5796;
	wire w5797;
	wire w5798;
	wire w5799;
	wire w5800;
	wire w5801;
	wire w5802;
	wire w5803;
	wire w5804;
	wire w5805;
	wire w5806;
	wire w5807;
	wire w5808;
	wire w5809;
	wire w5810;
	wire w5811;
	wire w5812;
	wire w5813;
	wire w5814;
	wire w5815;
	wire w5816;
	wire w5817;
	wire w5818;
	wire w5819;
	wire w5820;
	wire w5821;
	wire w5822;
	wire w5823;
	wire w5824;
	wire w5825;
	wire w5826;
	wire w5827;
	wire w5828;
	wire w5829;
	wire w5830;
	wire w5831;
	wire w5832;
	wire w5833;
	wire w5834;
	wire w5835;
	wire w5836;
	wire w5837;
	wire w5838;
	wire w5839;
	wire w5840;
	wire w5841;
	wire w5842;
	wire w5843;
	wire w5844;
	wire w5845;
	wire w5846;
	wire w5847;
	wire w5848;
	wire w5849;
	wire w5850;
	wire w5851;
	wire w5852;
	wire w5853;
	wire w5854;
	wire w5855;
	wire w5856;
	wire w5857;
	wire w5858;
	wire w5859;
	wire w5860;
	wire w5861;
	wire w5862;
	wire w5863;
	wire w5864;
	wire w5865;
	wire w5866;
	wire w5867;
	wire w5868;
	wire w5869;
	wire w5870;
	wire w5871;
	wire w5872;
	wire w5873;
	wire w5874;
	wire w5875;
	wire w5876;
	wire w5877;
	wire w5878;
	wire w5879;
	wire w5880;
	wire w5881;
	wire w5882;
	wire w5883;
	wire w5884;
	wire w5885;
	wire w5886;
	wire w5887;
	wire w5888;
	wire w5889;
	wire w5890;
	wire w5891;
	wire w5892;
	wire w5893;
	wire w5894;
	wire w5895;
	wire w5896;
	wire w5897;
	wire w5898;
	wire w5899;
	wire w5900;
	wire w5901;
	wire w5902;
	wire w5903;
	wire w5904;
	wire w5905;
	wire w5906;
	wire w5907;
	wire w5908;
	wire w5909;
	wire w5910;
	wire w5911;
	wire w5912;
	wire w5913;
	wire w5914;
	wire w5915;
	wire w5916;
	wire w5917;
	wire w5918;
	wire w5919;
	wire w5920;
	wire w5921;
	wire w5922;
	wire w5923;
	wire w5924;
	wire w5925;
	wire w5926;
	wire w5927;
	wire w5928;
	wire w5929;
	wire w5930;
	wire w5931;
	wire w5932;
	wire w5933;
	wire w5934;
	wire w5935;
	wire w5936;
	wire w5937;
	wire w5938;
	wire w5939;
	wire w5940;
	wire w5941;
	wire w5942;
	wire w5943;
	wire w5944;
	wire w5945;
	wire w5946;
	wire w5947;
	wire w5948;
	wire w5949;
	wire w5950;
	wire w5951;
	wire w5952;
	wire w5953;
	wire w5954;
	wire w5955;
	wire w5956;
	wire w5957;
	wire w5958;
	wire w5959;
	wire w5960;
	wire w5961;
	wire w5962;
	wire w5963;
	wire w5964;
	wire w5965;
	wire w5966;
	wire w5967;
	wire w5968;
	wire w5969;
	wire w5970;
	wire w5971;
	wire w5972;
	wire w5973;
	wire w5974;
	wire w5975;
	wire w5976;
	wire w5977;
	wire w5978;
	wire w5979;
	wire w5980;
	wire w5981;
	wire w5982;
	wire w5983;
	wire w5984;
	wire w5985;
	wire w5986;
	wire w5987;
	wire w5988;
	wire w5989;
	wire w5990;
	wire w5991;
	wire w5992;
	wire w5993;
	wire w5994;
	wire w5995;
	wire w5996;
	wire w5997;
	wire w5998;
	wire w5999;
	wire w6000;
	wire w6001;
	wire w6002;
	wire w6003;
	wire w6004;
	wire w6005;
	wire w6006;
	wire w6007;
	wire w6008;
	wire w6009;
	wire w6010;
	wire w6011;
	wire w6012;
	wire w6013;
	wire w6014;
	wire w6015;
	wire w6016;
	wire w6017;
	wire w6018;
	wire w6019;
	wire w6020;
	wire w6021;
	wire w6022;
	wire w6023;
	wire w6024;
	wire w6025;
	wire w6026;
	wire w6027;
	wire w6028;
	wire w6029;
	wire w6030;
	wire w6031;
	wire w6032;
	wire w6033;
	wire w6034;
	wire w6035;
	wire w6036;
	wire w6037;
	wire w6038;
	wire w6039;
	wire w6040;
	wire w6041;
	wire w6042;
	wire w6043;
	wire w6044;
	wire w6045;
	wire w6046;
	wire w6047;
	wire w6048;
	wire w6049;
	wire w6050;
	wire w6051;
	wire w6052;
	wire w6053;
	wire w6054;
	wire w6055;
	wire w6056;
	wire w6057;
	wire w6058;
	wire w6059;
	wire w6060;
	wire w6061;
	wire w6062;
	wire w6063;
	wire w6064;
	wire w6065;
	wire w6066;
	wire w6067;
	wire w6068;
	wire w6069;
	wire w6070;
	wire w6071;
	wire w6072;
	wire w6073;
	wire w6074;
	wire w6075;
	wire w6076;
	wire w6077;
	wire w6078;
	wire w6079;
	wire w6080;
	wire w6081;
	wire w6082;
	wire w6083;
	wire w6084;
	wire w6085;
	wire w6086;
	wire w6087;
	wire w6088;
	wire w6089;
	wire w6090;
	wire w6091;
	wire w6092;
	wire w6093;
	wire w6094;
	wire w6095;
	wire w6096;
	wire w6097;
	wire w6098;
	wire w6099;
	wire w6100;
	wire w6101;
	wire w6102;
	wire w6103;
	wire w6104;
	wire w6105;
	wire w6106;
	wire w6107;
	wire w6108;
	wire w6109;
	wire w6110;
	wire w6111;
	wire w6112;
	wire w6113;
	wire w6114;
	wire w6115;
	wire w6116;
	wire w6117;
	wire w6118;
	wire w6119;
	wire w6120;
	wire w6121;
	wire w6122;
	wire w6123;
	wire w6124;
	wire w6125;
	wire w6126;
	wire w6127;
	wire w6128;
	wire w6129;
	wire w6130;
	wire w6131;
	wire w6132;
	wire w6133;
	wire w6134;
	wire w6135;
	wire w6136;
	wire w6137;
	wire w6138;
	wire w6139;
	wire w6140;
	wire w6141;
	wire w6142;
	wire w6143;
	wire w6144;
	wire w6145;
	wire w6146;
	wire w6147;
	wire w6148;
	wire w6149;
	wire w6150;
	wire w6151;
	wire w6152;
	wire w6153;
	wire w6154;
	wire w6155;
	wire w6156;
	wire w6157;
	wire w6158;
	wire w6159;
	wire w6160;
	wire w6161;
	wire w6162;
	wire w6163;
	wire w6164;
	wire w6165;
	wire w6166;
	wire w6167;
	wire w6168;
	wire w6169;
	wire w6170;
	wire w6171;
	wire w6172;
	wire w6173;
	wire w6174;
	wire w6175;
	wire w6176;
	wire w6177;
	wire w6178;
	wire w6179;
	wire w6180;
	wire w6181;
	wire w6182;
	wire w6183;
	wire w6184;
	wire w6185;
	wire w6186;
	wire w6187;
	wire w6188;
	wire w6189;
	wire w6190;
	wire w6191;
	wire w6192;
	wire w6193;
	wire w6194;
	wire w6195;
	wire w6196;
	wire w6197;
	wire w6198;
	wire w6199;
	wire w6200;
	wire w6201;
	wire w6202;
	wire w6203;
	wire w6204;
	wire w6205;
	wire w6206;
	wire w6207;
	wire w6208;
	wire w6209;
	wire w6210;
	wire w6211;
	wire w6212;
	wire w6213;
	wire w6214;
	wire w6215;
	wire w6216;
	wire w6217;
	wire w6218;
	wire w6219;
	wire w6220;
	wire w6221;
	wire w6222;
	wire w6223;
	wire w6224;
	wire w6225;
	wire w6226;
	wire w6227;
	wire w6228;
	wire w6229;
	wire w6230;
	wire w6231;
	wire w6232;
	wire w6233;
	wire w6234;
	wire w6235;
	wire w6236;
	wire w6237;
	wire w6238;
	wire w6239;
	wire w6240;
	wire w6241;
	wire w6242;
	wire w6243;
	wire w6244;
	wire w6245;
	wire w6246;
	wire w6247;
	wire w6248;
	wire w6249;
	wire w6250;
	wire w6251;
	wire w6252;
	wire w6253;
	wire w6254;
	wire w6255;
	wire w6256;
	wire w6257;
	wire w6258;
	wire w6259;
	wire w6260;
	wire w6261;
	wire w6262;
	wire w6263;
	wire w6264;
	wire w6265;
	wire w6266;
	wire w6267;
	wire w6268;
	wire w6269;
	wire w6270;
	wire w6271;
	wire w6272;
	wire w6273;
	wire w6274;
	wire w6275;
	wire w6276;
	wire w6277;
	wire w6278;
	wire w6279;
	wire w6280;
	wire w6281;
	wire w6282;
	wire w6283;
	wire w6284;
	wire w6285;
	wire w6286;
	wire w6287;
	wire w6288;
	wire w6289;
	wire w6290;
	wire w6291;
	wire w6292;
	wire w6293;
	wire w6294;
	wire w6295;
	wire w6296;
	wire w6297;
	wire w6298;
	wire w6299;
	wire w6300;
	wire w6301;
	wire w6302;
	wire w6303;
	wire w6304;
	wire w6305;
	wire w6306;
	wire w6307;
	wire w6308;
	wire w6309;
	wire w6310;
	wire w6311;
	wire w6312;
	wire w6313;
	wire w6314;
	wire w6315;
	wire w6316;
	wire w6317;
	wire w6318;
	wire w6319;
	wire w6320;
	wire w6321;
	wire w6322;
	wire w6323;
	wire w6324;
	wire w6325;
	wire w6326;
	wire w6327;
	wire w6328;
	wire w6329;
	wire w6330;
	wire w6331;
	wire w6332;
	wire w6333;
	wire w6334;
	wire w6335;
	wire w6336;
	wire w6337;
	wire w6338;
	wire w6339;
	wire w6340;
	wire w6341;
	wire w6342;
	wire w6343;
	wire w6344;
	wire w6345;
	wire w6346;
	wire w6347;
	wire w6348;
	wire w6349;
	wire w6350;
	wire w6351;
	wire w6352;
	wire w6353;
	wire w6354;
	wire w6355;
	wire w6356;
	wire w6357;
	wire w6358;
	wire w6359;
	wire w6360;
	wire w6361;
	wire w6362;
	wire w6363;
	wire w6364;
	wire w6365;
	wire w6366;
	wire w6367;
	wire w6368;
	wire w6369;
	wire w6370;
	wire w6371;
	wire w6372;
	wire w6373;
	wire w6374;
	wire w6375;
	wire w6376;
	wire w6377;
	wire w6378;
	wire w6379;
	wire w6380;
	wire w6381;
	wire w6382;
	wire w6383;
	wire w6384;
	wire w6385;
	wire w6386;
	wire w6387;
	wire w6388;
	wire w6389;
	wire w6390;
	wire w6391;
	wire w6392;
	wire w6393;
	wire w6394;
	wire w6395;
	wire w6396;
	wire w6397;
	wire w6398;
	wire w6399;
	wire w6400;
	wire w6401;
	wire w6402;
	wire w6403;
	wire w6404;
	wire w6405;
	wire w6406;
	wire w6407;
	wire w6408;
	wire w6409;
	wire w6410;
	wire w6411;
	wire w6412;
	wire w6413;
	wire w6414;
	wire w6415;
	wire w6416;
	wire w6417;
	wire w6418;
	wire w6419;
	wire w6420;
	wire w6421;
	wire w6422;
	wire w6423;
	wire w6424;
	wire w6425;
	wire w6426;
	wire w6427;
	wire w6428;
	wire w6429;
	wire w6430;
	wire w6431;
	wire w6432;
	wire w6433;
	wire w6434;
	wire w6435;
	wire w6436;
	wire w6437;
	wire w6438;
	wire w6439;
	wire w6440;
	wire w6441;
	wire w6442;
	wire w6443;
	wire w6444;
	wire w6445;
	wire w6446;
	wire w6447;
	wire w6448;
	wire w6449;
	wire w6450;
	wire w6451;
	wire w6452;
	wire w6453;
	wire w6454;
	wire w6455;
	wire w6456;
	wire w6457;
	wire w6458;
	wire w6459;
	wire w6460;
	wire w6461;
	wire w6462;
	wire w6463;
	wire w6464;
	wire w6465;
	wire w6466;
	wire w6467;
	wire w6468;
	wire w6469;
	wire w6470;
	wire w6471;
	wire w6472;
	wire w6473;
	wire w6474;
	wire w6475;
	wire w6476;
	wire w6477;
	wire w6478;
	wire w6479;
	wire w6480;
	wire w6481;
	wire w6482;
	wire w6483;
	wire w6484;
	wire w6485;
	wire w6486;
	wire w6487;
	wire w6488;
	wire w6489;
	wire w6490;
	wire w6491;
	wire w6492;
	wire w6493;
	wire w6494;
	wire w6495;
	wire w6496;
	wire w6497;
	wire w6498;
	wire w6499;
	wire w6500;
	wire w6501;
	wire w6502;
	wire w6503;
	wire w6504;
	wire w6505;
	wire w6506;
	wire w6507;
	wire w6508;
	wire w6509;
	wire w6510;
	wire w6511;
	wire w6512;
	wire w6513;
	wire w6514;
	wire w6515;
	wire w6516;
	wire w6517;
	wire w6518;
	wire w6519;
	wire w6520;
	wire w6521;
	wire w6522;
	wire w6523;
	wire w6524;
	wire w6525;
	wire w6526;
	wire w6527;
	wire w6528;
	wire w6529;
	wire w6530;
	wire w6531;
	wire w6532;
	wire w6533;
	wire w6534;
	wire w6535;
	wire w6536;
	wire w6537;
	wire w6538;
	wire w6539;
	wire w6540;
	wire w6541;
	wire w6542;
	wire w6543;
	wire w6544;
	wire w6545;
	wire w6546;
	wire w6547;
	wire w6548;
	wire w6549;
	wire w6550;
	wire w6551;
	wire w6552;
	wire w6553;
	wire w6554;
	wire w6555;
	wire w6556;
	wire w6557;
	wire w6558;
	wire w6559;
	wire w6560;
	wire w6561;
	wire w6562;
	wire w6563;
	wire w6564;
	wire w6565;
	wire w6566;
	wire w6567;
	wire w6568;
	wire w6569;
	wire w6570;
	wire w6571;
	wire w6572;
	wire w6573;
	wire w6574;
	wire w6575;
	wire w6576;
	wire w6577;
	wire w6578;
	wire w6579;
	wire w6580;
	wire w6581;
	wire w6582;
	wire w6583;
	wire w6584;
	wire w6585;
	wire w6586;
	wire w6587;
	wire w6588;
	wire w6589;
	wire w6590;
	wire w6591;
	wire w6592;
	wire w6593;
	wire w6594;
	wire w6595;
	wire w6596;
	wire w6597;
	wire w6598;
	wire w6599;
	wire w6600;
	wire w6601;
	wire w6602;
	wire w6603;
	wire w6604;
	wire w6605;
	wire w6606;
	wire w6607;
	wire w6608;
	wire w6609;
	wire w6610;
	wire w6611;
	wire w6612;
	wire w6613;
	wire w6614;
	wire w6615;
	wire w6616;
	wire w6617;
	wire w6618;
	wire w6619;
	wire w6620;
	wire w6621;
	wire w6622;
	wire w6623;
	wire w6624;
	wire w6625;
	wire w6626;
	wire w6627;
	wire w6628;
	wire w6629;
	wire w6630;
	wire w6631;
	wire w6632;
	wire w6633;
	wire w6634;
	wire w6635;
	wire w6636;
	wire w6637;
	wire w6638;
	wire w6639;
	wire w6640;
	wire w6641;
	wire w6642;
	wire w6643;
	wire w6644;
	wire w6645;
	wire w6646;
	wire w6647;
	wire w6648;
	wire w6649;
	wire w6650;
	wire w6651;
	wire w6652;
	wire w6653;
	wire w6654;
	wire w6655;
	wire w6656;
	wire w6657;
	wire w6658;
	wire w6659;
	wire w6660;
	wire w6661;
	wire w6662;
	wire w6663;
	wire w6664;
	wire w6665;
	wire w6666;
	wire w6667;
	wire w6668;
	wire w6669;
	wire w6670;
	wire w6671;
	wire w6672;
	wire w6673;
	wire w6674;
	wire w6675;
	wire w6676;
	wire w6677;
	wire w6678;
	wire w6679;
	wire w6680;
	wire w6681;
	wire w6682;
	wire w6683;
	wire w6684;
	wire w6685;
	wire w6686;
	wire w6687;
	wire w6688;
	wire w6689;
	wire w6690;
	wire w6691;
	wire w6692;
	wire w6693;
	wire w6694;
	wire w6695;
	wire w6696;
	wire w6697;
	wire w6698;
	wire w6699;
	wire w6700;
	wire w6701;
	wire w6702;
	wire w6703;
	wire w6704;
	wire w6705;
	wire w6706;
	wire w6707;
	wire w6708;
	wire w6709;
	wire w6710;
	wire w6711;
	wire w6712;
	wire w6713;
	wire w6714;
	wire w6715;
	wire w6716;
	wire w6717;
	wire w6718;
	wire w6719;
	wire w6720;
	wire w6721;
	wire w6722;
	wire w6723;
	wire w6724;
	wire w6725;
	wire w6726;
	wire w6727;
	wire w6728;
	wire w6729;
	wire w6730;
	wire w6731;
	wire w6732;
	wire w6733;
	wire w6734;
	wire w6735;
	wire w6736;
	wire w6737;
	wire w6738;
	wire w6739;
	wire w6740;
	wire w6741;
	wire w6742;
	wire w6743;
	wire w6744;
	wire w6745;
	wire w6746;
	wire w6747;
	wire w6748;
	wire w6749;
	wire w6750;
	wire w6751;
	wire w6752;
	wire w6753;
	wire w6754;
	wire w6755;
	wire w6756;
	wire w6757;
	wire w6758;
	wire w6759;
	wire w6760;
	wire w6761;
	wire w6762;
	wire w6763;
	wire w6764;
	wire w6765;
	wire w6766;
	wire w6767;
	wire w6768;
	wire w6769;
	wire w6770;
	wire w6771;
	wire w6772;
	wire w6773;
	wire w6774;
	wire w6775;
	wire w6776;
	wire w6777;
	wire w6778;
	wire w6779;
	wire w6780;
	wire w6781;
	wire w6782;
	wire w6783;
	wire w6784;
	wire w6785;
	wire w6786;
	wire w6787;
	wire w6788;
	wire w6789;
	wire w6790;
	wire w6791;
	wire w6792;
	wire w6793;
	wire w6794;
	wire w6795;
	wire w6796;
	wire w6797;
	wire w6798;
	wire w6799;
	wire w6800;
	wire w6801;
	wire w6802;
	wire w6803;
	wire w6804;
	wire w6805;
	wire w6806;

	assign CH0_EN = w2009;
	assign CH0VOL[0] = w2012;
	assign CH0VOL[1] = w2013;
	assign CH1_EN = w2010;
	assign CH1VOL[0] = w2072;
	assign CH1VOL[1] = w2073;
	assign CH2_EN = w2007;
	assign CH2VOL[0] = w2092;
	assign CH2VOL[1] = w2091;
	assign CH3_EN = w2008;
	assign CH3VOL[0] = w2114;
	assign CH3VOL[1] = w2113;
	assign PSGDAC0[0] = w2014;
	assign PSGDAC0[1] = w2015;
	assign PSGDAC0[2] = w2016;
	assign PSGDAC0[3] = w2017;
	assign PSGDAC0[4] = w2018;
	assign PSGDAC0[5] = w2019;
	assign PSGDAC0[6] = w2020;
	assign PSGDAC0[7] = w2021;
	assign PSGDAC1[0] = w2074;
	assign PSGDAC1[1] = w2075;
	assign PSGDAC1[2] = w2076;
	assign PSGDAC1[3] = w2077;
	assign PSGDAC1[4] = w2078;
	assign PSGDAC1[5] = w2079;
	assign PSGDAC1[6] = w2080;
	assign PSGDAC1[7] = w2081;
	assign PSGDAC2[0] = w2103;
	assign PSGDAC2[1] = w2104;
	assign PSGDAC2[2] = w2105;
	assign PSGDAC2[3] = w2106;
	assign PSGDAC2[4] = w2107;
	assign PSGDAC2[5] = w2108;
	assign PSGDAC2[6] = w2109;
	assign PSGDAC2[7] = w2110;
	assign PSGDAC3[0] = w2112;
	assign PSGDAC3[1] = w2111;
	assign PSGDAC3[2] = w2119;
	assign PSGDAC3[3] = w2118;
	assign PSGDAC3[4] = w2117;
	assign PSGDAC3[5] = w2116;
	assign PSGDAC3[6] = w2115;
	assign PSGDAC3[7] = w2120;
	assign w1201 = CAi[22];
	assign CAo[22] = w1358;
	assign CA[19] = CA[19];
	assign DTACK_OUT = w1051;
	assign Z80_INT = w1052;
	assign RA[7] = w1109;
	assign RA[6] = w1108;
	assign RA[5] = w1107;
	assign RA[4] = w1106;
	assign RA[2] = w1104;
	assign RA[1] = w1103;
	assign RA[0] = w1102;
	assign nRAS0 = w1334;
	assign RA[3] = w1105;
	assign nCAS0 = w1407;
	assign nOE0 = w1398;
	assign nLWR = w1399;
	assign nUWR = w1309;
	assign w1386 = DTACK_IN;
	assign w996 = RnW;
	assign w1378 = nLDS;
	assign w1369 = nUDS;
	assign w1252 = nAS;
	assign w1367 = nM1;
	assign w1368 = nWR;
	assign w1365 = nRD;
	assign w1366 = nIORQ;
	assign nILP2 = w1371;
	assign nILP1 = w1370;
	assign w1233 = nINTAK;
	assign w1364 = nMREQ;
	assign w1235 = nBG;
	assign BGACK_OUT = w1250;
	assign w1385 = BGACK_IN;
	assign nBR = w1428;
	assign VSYNC = w1696;
	assign nCSYNC = w1995;
	assign w1690 = nCSYNC_IN;
	assign nHSYNC = w1753;
	assign w1965 = nHSYNC_IN;
	assign DB[15] = DB[15];
	assign DB[14] = DB[14];
	assign DB[13] = DB[13];
	assign DB[12] = DB[12];
	assign DB[11] = DB[11];
	assign DB[10] = DB[10];
	assign DB[9] = DB[9];
	assign DB[8] = DB[8];
	assign DB[7] = DB[7];
	assign DB[6] = DB[6];
	assign DB[5] = DB[5];
	assign DB[4] = DB[4];
	assign DB[3] = DB[3];
	assign DB[2] = DB[2];
	assign DB[1] = DB[1];
	assign DB[0] = DB[0];
	assign CA[0] = CA[0];
	assign CA[1] = CA[1];
	assign CA[2] = CA[2];
	assign CA[3] = CA[3];
	assign CA[4] = CA[4];
	assign CA[5] = CA[5];
	assign CA[6] = CA[6];
	assign CA[7] = CA[7];
	assign CA[8] = CA[8];
	assign CA[9] = CA[9];
	assign CA[10] = CA[10];
	assign CA[11] = CA[11];
	assign CA[12] = CA[12];
	assign CA[13] = CA[13];
	assign CA[14] = CA[14];
	assign CA[15] = CA[15];
	assign CA[17] = CA[17];
	assign CA[18] = CA[18];
	assign CA[20] = CA[20];
	assign CA[21] = CA[21];
	assign R_DAC[0] = w2946;
	assign R_DAC[1] = w2911;
	assign R_DAC[2] = w2945;
	assign R_DAC[3] = w2910;
	assign R_DAC[4] = w2944;
	assign R_DAC[5] = w2943;
	assign R_DAC[6] = w2942;
	assign R_DAC[7] = w2941;
	assign R_DAC[8] = w2907;
	assign G_DAC[0] = w2939;
	assign G_DAC[1] = w2938;
	assign G_DAC[2] = w2901;
	assign G_DAC[3] = w2900;
	assign G_DAC[4] = w2899;
	assign G_DAC[5] = w2898;
	assign G_DAC[6] = w2897;
	assign G_DAC[7] = w2896;
	assign G_DAC[8] = w2895;
	assign R_DAC[9] = w2908;
	assign R_DAC[10] = w2905;
	assign R_DAC[11] = w2909;
	assign R_DAC[12] = w2904;
	assign R_DAC[13] = w2906;
	assign R_DAC[14] = w2903;
	assign R_DAC[15] = w2902;
	assign R_DAC[16] = w2940;
	assign B_DAC[0] = w2887;
	assign B_DAC[1] = w2937;
	assign B_DAC[2] = w2933;
	assign B_DAC[3] = w2934;
	assign B_DAC[4] = w2935;
	assign B_DAC[5] = w2932;
	assign B_DAC[6] = w2936;
	assign B_DAC[7] = w2994;
	assign B_DAC[8] = w2888;
	assign G_DAC[9] = w2889;
	assign G_DAC[10] = w2894;
	assign G_DAC[11] = w2893;
	assign G_DAC[12] = w2992;
	assign G_DAC[13] = w2892;
	assign G_DAC[14] = w2891;
	assign G_DAC[15] = w2890;
	assign G_DAC[16] = w2993;
	assign B_DAC[9] = w2885;
	assign B_DAC[10] = w2886;
	assign B_DAC[11] = w2931;
	assign B_DAC[12] = w2930;
	assign B_DAC[13] = w2929;
	assign B_DAC[14] = w2928;
	assign B_DAC[15] = w2926;
	assign B_DAC[16] = w2927;
	assign nOE1 = nOE1;
	assign nWE0 = nWE0;
	assign nWE1 = nWE1;
	assign nCAS1 = nCAS1;
	assign nRAS1 = nRAS1;
	assign AD_RD_DIR = AD_RD_DIR;
	assign nYS = nYS;
	assign nSC = w2594;
	assign nSE0_1 = w2487;
	assign ADo[7] = w2447;
	assign ADo[6] = w2455;
	assign ADo[5] = w2632;
	assign ADo[4] = w2462;
	assign ADo[3] = w2572;
	assign ADo[2] = w2571;
	assign ADo[1] = w2523;
	assign ADo[0] = w2686;
	assign RDo[6] = w2633;
	assign RDo[5] = w2663;
	assign RDo[4] = w2638;
	assign RDo[3] = w2637;
	assign RDo[2] = w2665;
	assign RDo[1] = w2687;
	assign RDo[0] = w2494;
	assign w2534 = RDi[6];
	assign w2448 = RDi[7];
	assign w2461 = RDi[4];
	assign w2676 = RDi[5];
	assign w2528 = RDi[2];
	assign w2536 = RDi[3];
	assign w2666 = RDi[0];
	assign w2570 = RDi[1];
	assign w2535 = ADi[6];
	assign w2636 = ADi[7];
	assign w2480 = ADi[4];
	assign w2664 = ADi[5];
	assign w2522 = ADi[2];
	assign w2527 = ADi[3];
	assign w2495 = ADi[0];
	assign w2514 = ADi[1];
	assign RDo[7] = w2635;
	assign w5260 = SD[7];
	assign w5261 = SD[6];
	assign w6661 = SD[5];
	assign w6663 = SD[4];
	assign w5262 = SD[3];
	assign w5259 = SD[2];
	assign w6662 = SD[1];
	assign w5258 = SD[0];
	assign CLK1 = 68K CPU CLOCK;
	assign CLK0 = w1401;
	assign w4467 = EDCLKi;
	assign EDCLKo = EDCLK_O;
	assign w4443 = MCLK;
	assign SUB_CLK = w4432;
	assign w4485 = nRES_PAD;
	assign w1429 = 68kCLKi;
	assign EDCLKd = w1485;
	assign CA_PAD_DIR = w2444;
	assign DB_PAD_DIR = w2445;
	assign w403 = SEL0_M3;
	assign w6667 = nPAL;
	assign w436 = nHL;
	assign SPA/Bo = w2811;
	assign w2788 = SPA/Bi;

	// Instances

	vdp_slatch g1 (.nQ(w351), .D(VPOS[7]), .C(w1556), .nC(w1557) );
	vdp_slatch g2 (.nQ(w1519), .D(HPOS[8]), .C(w372), .nC(w373) );
	vdp_slatch g3 (.nQ(w356), .D(w298), .C(w1458), .nC(w374) );
	vdp_slatch g4 (.D(w299), .C(w1554), .nC(w1555), .nQ(w6769) );
	vdp_slatch g5 (.nQ(w357), .D(w358), .C(w1552), .nC(w1553) );
	vdp_slatch g6 (.nQ(w301), .D(w302), .C(w1550), .nC(w1551) );
	vdp_slatch g7 (.nQ(w359), .D(w358), .C(w375), .nC(w376) );
	vdp_slatch g8 (.nQ(w362), .D(w302), .C(w377), .nC(w378) );
	vdp_slatch g9 (.nQ(w360), .D(w358), .C(w425), .nC(w1455) );
	vdp_slatch g10 (.nQ(w363), .D(w302), .C(w1454), .nC(w383) );
	vdp_slatch g11 (.nQ(w361), .D(w358), .C(w381), .nC(w380) );
	vdp_slatch g12 (.nQ(w304), .D(w302), .C(w379), .nC(w1453) );
	vdp_slatch g13 (.Q(w302), .D(DB[7]), .C(w365), .nC(w364) );
	vdp_slatch g14 (.Q(w358), .D(w926), .C(w368), .nC(w367) );
	vdp_sr_bit g15 (.D(w305), .C2(HCLK2), .C1(HCLK1), .Q(FIFOo[7]), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g16 (.A(1'b1), .nZ(DB[7]), .nE(w1452) );
	vdp_notif0 g17 (.A(w304), .nZ(w305), .nE(w2011) );
	vdp_notif0 g18 (.A(w361), .nZ(w355), .nE(w382) );
	vdp_notif0 g19 (.A(w303), .nZ(AD_DATA[7]), .nE(w1598) );
	vdp_notif0 g20 (.A(w363), .nZ(w305), .nE(w1549) );
	vdp_notif0 g21 (.A(w360), .nZ(w355), .nE(w1597) );
	vdp_notif0 g22 (.A(w1525), .nZ(AD_DATA[7]), .nE(w400) );
	vdp_notif0 g23 (.A(w362), .nZ(w305), .nE(w399) );
	vdp_notif0 g24 (.A(w359), .nZ(w355), .nE(w1456) );
	vdp_notif0 g25 (.A(w1524), .nZ(AD_DATA[7]), .nE(w414) );
	vdp_notif0 g26 (.A(w301), .nZ(w305), .nE(w392) );
	vdp_notif0 g27 (.A(w300), .nZ(AD_DATA[7]), .nE(w412) );
	vdp_notif0 g28 (.A(w356), .nZ(DB[7]), .nE(w1595) );
	vdp_notif0 g29 (.nZ(DB[15]), .nE(w393), .A(w6769) );
	vdp_notif0 g30 (.A(w357), .nZ(w355), .nE(w1596) );
	vdp_notif0 g31 (.A(w351), .nZ(DB[15]), .nE(w1594) );
	vdp_notif0 g32 (.A(w428), .nZ(DB[7]), .nE(w394) );
	vdp_aon22 g33 (.Z(w428), .A1(w1519), .A2(w1558), .B1(w398), .B2(w351) );
	vdp_aon22 g34 (.A2(w396), .B1(w397), .B2(AD_DATA[7]), .A1(w355), .Z(w298) );
	vdp_aon22 g35 (.A2(w6675), .B1(w6676), .B2(w355), .A1(AD_DATA[7]), .Z(w299) );
	vdp_aon22 g36 (.Z(w300), .A2(w395), .B1(w1559), .B2(w301), .A1(w357) );
	vdp_aon22 g37 (.Z(w1524), .A2(w419), .B1(w418), .B2(w359), .A1(w362) );
	vdp_aon22 g38 (.Z(w1525), .A2(w426), .B1(w427), .B2(w360), .A1(w363) );
	vdp_aon22 g39 (.Z(w303), .A2(w6671), .B1(w6672), .B2(w304), .A1(w361) );
	vdp_aon22 g40 (.Z(w926), .A1(DB[15]), .A2(w366), .B1(w370), .B2(DB[7]) );
	vdp_slatch g41 (.nQ(w220), .D(VPOS[6]), .C(w1556), .nC(w1557) );
	vdp_slatch g42 (.nQ(w223), .D(HPOS[7]), .C(w372), .nC(w373) );
	vdp_slatch g43 (.nQ(w225), .D(w261), .C(w1458), .nC(w374) );
	vdp_slatch g44 (.nQ(w263), .D(w1425), .C(w1554), .nC(w1555) );
	vdp_slatch g45 (.nQ(w226), .D(w227), .C(w1552), .nC(w1553) );
	vdp_slatch g46 (.nQ(w265), .D(w266), .C(w1550), .nC(w1551) );
	vdp_slatch g47 (.nQ(w228), .D(w227), .C(w375), .nC(w376) );
	vdp_slatch g48 (.nQ(w230), .D(w266), .C(w377), .nC(w378) );
	vdp_slatch g49 (.nQ(w231), .D(w227), .C(w425), .nC(w1455) );
	vdp_slatch g50 (.nQ(w233), .D(w266), .C(w1454), .nC(w383) );
	vdp_slatch g51 (.nQ(w234), .D(w227), .C(w381), .nC(w380) );
	vdp_slatch g52 (.nQ(w268), .D(w266), .C(w379), .nC(w1453) );
	vdp_slatch g53 (.Q(w266), .D(DB[6]), .C(w365), .nC(w364) );
	vdp_slatch g54 (.Q(w227), .D(w269), .C(w368), .nC(w367) );
	vdp_sr_bit g55 (.D(w262), .Q(FIFOo[6]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g56 (.A(1'b1), .nZ(DB[6]), .nE(w1452) );
	vdp_notif0 g57 (.A(w268), .nZ(w262), .nE(w2011) );
	vdp_notif0 g58 (.A(w234), .nZ(RD_DATA[6]), .nE(w382) );
	vdp_notif0 g59 (.A(w267), .nZ(AD_DATA[6]), .nE(w1598) );
	vdp_notif0 g60 (.A(w233), .nZ(w262), .nE(w1549) );
	vdp_notif0 g61 (.A(w231), .nZ(RD_DATA[6]), .nE(w1597) );
	vdp_notif0 g62 (.A(w232), .nZ(AD_DATA[6]), .nE(w400) );
	vdp_notif0 g63 (.A(w230), .nZ(w262), .nE(w399) );
	vdp_notif0 g64 (.A(w228), .nZ(RD_DATA[6]), .nE(w1456) );
	vdp_notif0 g65 (.A(w229), .nZ(AD_DATA[6]), .nE(w414) );
	vdp_notif0 g66 (.A(w265), .nZ(w262), .nE(w392) );
	vdp_notif0 g67 (.A(w264), .nZ(AD_DATA[6]), .nE(w412) );
	vdp_notif0 g68 (.A(w225), .nZ(DB[6]), .nE(w1595) );
	vdp_notif0 g69 (.A(w263), .nZ(DB[14]), .nE(w393) );
	vdp_notif0 g70 (.A(w226), .nZ(RD_DATA[6]), .nE(w1596) );
	vdp_notif0 g71 (.A(w220), .nZ(DB[14]), .nE(w1594) );
	vdp_notif0 g72 (.A(w224), .nZ(DB[6]), .nE(w394) );
	vdp_aon22 g73 (.A2(w1558), .B1(w398), .B2(w220), .A1(w223), .Z(w224) );
	vdp_aon22 g74 (.Z(w261), .A2(w396), .B1(w397), .B2(AD_DATA[6]), .A1(RD_DATA[6]) );
	vdp_aon22 g75 (.Z(w1425), .A2(w6675), .B1(w6676), .B2(RD_DATA[6]), .A1(AD_DATA[6]) );
	vdp_aon22 g76 (.Z(w264), .A2(w395), .B1(w1559), .B2(w265), .A1(w226) );
	vdp_aon22 g77 (.Z(w229), .A2(w419), .B1(w418), .B2(w230), .A1(w228) );
	vdp_aon22 g78 (.Z(w232), .A2(w426), .B1(w427), .B2(w233), .A1(w231) );
	vdp_aon22 g79 (.Z(w267), .A2(w6671), .B1(w6672), .B2(w268), .A1(w234) );
	vdp_aon22 g80 (.Z(w269), .A1(DB[14]), .A2(w366), .B1(w370), .B2(DB[6]) );
	vdp_slatch g81 (.nQ(w335), .D(VPOS[5]), .C(w1556), .nC(w1557) );
	vdp_slatch g82 (.nQ(w1520), .D(HPOS[6]), .C(w372), .nC(w373) );
	vdp_slatch g83 (.nQ(w340), .D(w289), .C(w1458), .nC(w374) );
	vdp_slatch g84 (.D(w290), .C(w1554), .nC(w1555), .nQ(w6770) );
	vdp_slatch g85 (.nQ(w341), .D(w347), .C(w1552), .nC(w1553) );
	vdp_slatch g86 (.nQ(w292), .D(w293), .C(w1550), .nC(w1551) );
	vdp_slatch g87 (.nQ(w343), .D(w347), .C(w375), .nC(w376) );
	vdp_slatch g88 (.nQ(w342), .D(w293), .C(w377), .nC(w378) );
	vdp_slatch g89 (.nQ(w345), .D(w347), .C(w425), .nC(w1455) );
	vdp_slatch g90 (.nQ(w348), .D(w293), .C(w1454), .nC(w383) );
	vdp_slatch g91 (.nQ(w349), .D(w347), .C(w381), .nC(w380) );
	vdp_slatch g92 (.nQ(w295), .D(w293), .C(w379), .nC(w1453) );
	vdp_slatch g93 (.Q(w293), .D(DB[5]), .C(w365), .nC(w364) );
	vdp_slatch g94 (.Q(w347), .D(w296), .C(w368), .nC(w367) );
	vdp_sr_bit g95 (.D(w297), .Q(FIFOo[5]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g96 (.A(1'b1), .nZ(DB[5]), .nE(w1452) );
	vdp_notif0 g97 (.A(w295), .nZ(w297), .nE(w2011) );
	vdp_notif0 g98 (.A(w349), .nZ(RD_DATA[5]), .nE(w382) );
	vdp_notif0 g99 (.A(w294), .nZ(AD_DATA[5]), .nE(w1598) );
	vdp_notif0 g100 (.A(w348), .nZ(w297), .nE(w1549) );
	vdp_notif0 g101 (.A(w345), .nZ(RD_DATA[5]), .nE(w1597) );
	vdp_notif0 g102 (.A(w346), .nZ(AD_DATA[5]), .nE(w400) );
	vdp_notif0 g103 (.A(w342), .nZ(w297), .nE(w399) );
	vdp_notif0 g104 (.A(w343), .nZ(RD_DATA[5]), .nE(w1456) );
	vdp_notif0 g105 (.A(w344), .nZ(AD_DATA[5]), .nE(w414) );
	vdp_notif0 g106 (.A(w292), .nZ(w297), .nE(w392) );
	vdp_notif0 g107 (.A(w291), .nZ(AD_DATA[5]), .nE(w412) );
	vdp_notif0 g108 (.A(w340), .nZ(DB[5]), .nE(w1595) );
	vdp_notif0 g109 (.nZ(DB[13]), .nE(w393), .A(w6770) );
	vdp_notif0 g110 (.A(w341), .nZ(RD_DATA[5]), .nE(w1596) );
	vdp_notif0 g111 (.A(w335), .nZ(DB[13]), .nE(w1594) );
	vdp_notif0 g112 (.A(w339), .nZ(DB[5]), .nE(w394) );
	vdp_aon22 g113 (.Z(w339), .A1(w1520), .A2(w1558), .B1(w398), .B2(w335) );
	vdp_aon22 g114 (.A2(w396), .B1(w397), .B2(AD_DATA[5]), .A1(RD_DATA[5]), .Z(w289) );
	vdp_aon22 g115 (.A2(w6675), .B1(w6676), .B2(RD_DATA[5]), .A1(AD_DATA[5]), .Z(w290) );
	vdp_aon22 g116 (.Z(w291), .A2(w395), .B1(w1559), .B2(w292), .A1(w341) );
	vdp_aon22 g117 (.Z(w344), .A2(w419), .B1(w418), .B2(w343), .A1(w342) );
	vdp_aon22 g118 (.Z(w346), .A2(w426), .B1(w427), .B2(w345), .A1(w348) );
	vdp_aon22 g119 (.Z(w294), .A2(w6671), .B1(w6672), .B2(w295), .A1(w349) );
	vdp_aon22 g120 (.Z(w296), .A1(DB[13]), .A2(w366), .B1(w370), .B2(DB[5]) );
	vdp_slatch g121 (.nQ(w205), .D(VPOS[4]), .C(w1556), .nC(w1557) );
	vdp_slatch g122 (.nQ(w208), .D(HPOS[5]), .C(w372), .nC(w373) );
	vdp_slatch g123 (.nQ(w1560), .D(w253), .C(w1458), .nC(w374) );
	vdp_slatch g124 (.D(w1523), .C(w1554), .nC(w1555), .nQ(w6771) );
	vdp_slatch g125 (.nQ(w210), .D(w211), .C(w1552), .nC(w1553) );
	vdp_slatch g126 (.nQ(w256), .D(w257), .C(w1550), .nC(w1551) );
	vdp_slatch g127 (.nQ(w212), .D(w211), .C(w375), .nC(w376) );
	vdp_slatch g128 (.nQ(w214), .D(w257), .C(w377), .nC(w378) );
	vdp_slatch g129 (.nQ(w215), .D(w211), .C(w425), .nC(w1455) );
	vdp_slatch g130 (.nQ(w217), .D(w257), .C(w1454), .nC(w383) );
	vdp_slatch g131 (.nQ(w218), .D(w211), .C(w381), .nC(w380) );
	vdp_slatch g132 (.nQ(w259), .D(w257), .C(w379), .nC(w1453) );
	vdp_slatch g133 (.Q(w257), .D(DB[4]), .C(w365), .nC(w364) );
	vdp_slatch g134 (.Q(w211), .D(w260), .C(w368), .nC(w367) );
	vdp_sr_bit g135 (.D(w254), .Q(FIFOo[4]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g136 (.A(1'b1), .nZ(DB[4]), .nE(w1452) );
	vdp_notif0 g137 (.A(w259), .nZ(w254), .nE(w2011) );
	vdp_notif0 g138 (.A(w218), .nZ(RD_DATA[4]), .nE(w382) );
	vdp_notif0 g139 (.A(w258), .nZ(AD_DATA[4]), .nE(w1598) );
	vdp_notif0 g140 (.A(w217), .nZ(w254), .nE(w1549) );
	vdp_notif0 g141 (.A(w215), .nZ(RD_DATA[4]), .nE(w1597) );
	vdp_notif0 g142 (.A(w216), .nZ(AD_DATA[4]), .nE(w400) );
	vdp_notif0 g143 (.A(w214), .nZ(w254), .nE(w399) );
	vdp_notif0 g144 (.A(w212), .nZ(RD_DATA[4]), .nE(w1456) );
	vdp_notif0 g145 (.A(w213), .nZ(AD_DATA[4]), .nE(w414) );
	vdp_notif0 g146 (.A(w256), .nZ(w254), .nE(w392) );
	vdp_notif0 g147 (.A(w255), .nZ(AD_DATA[4]), .nE(w412) );
	vdp_notif0 g148 (.A(w1560), .nZ(DB[4]), .nE(w1595) );
	vdp_notif0 g149 (.nZ(DB[12]), .nE(w393), .A(w6771) );
	vdp_notif0 g150 (.A(w210), .nZ(RD_DATA[4]), .nE(w1596) );
	vdp_notif0 g151 (.A(w205), .nZ(DB[12]), .nE(w1594) );
	vdp_notif0 g152 (.A(w209), .nZ(DB[4]), .nE(w394) );
	vdp_aon22 g153 (.A2(w1558), .B1(w398), .B2(w205), .A1(w208), .Z(w209) );
	vdp_aon22 g154 (.Z(w253), .A2(w396), .B1(w397), .B2(AD_DATA[4]), .A1(RD_DATA[4]) );
	vdp_aon22 g155 (.Z(w1523), .A2(w6675), .B1(w6676), .B2(RD_DATA[4]), .A1(AD_DATA[4]) );
	vdp_aon22 g156 (.Z(w255), .A2(w395), .B1(w1559), .B2(w256), .A1(w210) );
	vdp_aon22 g157 (.Z(w213), .A2(w419), .B1(w418), .B2(w214), .A1(w212) );
	vdp_aon22 g158 (.Z(w216), .A2(w426), .B1(w427), .B2(w217), .A1(w215) );
	vdp_aon22 g159 (.Z(w258), .A2(w6671), .B1(w6672), .B2(w259), .A1(w218) );
	vdp_aon22 g160 (.Z(w260), .A1(DB[12]), .A2(w366), .B1(w370), .B2(DB[4]) );
	vdp_slatch g161 (.nQ(w319), .D(VPOS[3]), .C(w1556), .nC(w1557) );
	vdp_slatch g162 (.nQ(w1521), .D(HPOS[4]), .C(w372), .nC(w373) );
	vdp_slatch g163 (.nQ(w324), .D(w280), .C(w1458), .nC(w374) );
	vdp_slatch g164 (.D(w281), .C(w1554), .nC(w1555), .nQ(w6772) );
	vdp_slatch g165 (.nQ(w325), .D(w328), .C(w1552), .nC(w1553) );
	vdp_slatch g166 (.nQ(w283), .D(w284), .C(w1550), .nC(w1551) );
	vdp_slatch g167 (.nQ(w326), .D(w328), .C(w375), .nC(w376) );
	vdp_slatch g168 (.nQ(w327), .D(w284), .C(w377), .nC(w378) );
	vdp_slatch g169 (.nQ(w330), .D(w328), .C(w425), .nC(w1455) );
	vdp_slatch g170 (.nQ(w332), .D(w284), .C(w1454), .nC(w383) );
	vdp_slatch g171 (.nQ(w333), .D(w328), .C(w381), .nC(w380) );
	vdp_slatch g172 (.nQ(w286), .D(w284), .C(w379), .nC(w1453) );
	vdp_slatch g173 (.Q(w284), .D(DB[3]), .C(w365), .nC(w364) );
	vdp_slatch g174 (.Q(w328), .D(w287), .C(w368), .nC(w367) );
	vdp_sr_bit g175 (.D(w288), .Q(FIFOo[3]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g176 (.A(1'b1), .nZ(DB[3]), .nE(w1452) );
	vdp_notif0 g177 (.A(w286), .nZ(w288), .nE(w2011) );
	vdp_notif0 g178 (.A(w333), .nZ(w321), .nE(w382) );
	vdp_notif0 g179 (.A(w285), .nZ(AD_DATA[3]), .nE(w1598) );
	vdp_notif0 g180 (.A(w332), .nZ(w288), .nE(w1549) );
	vdp_notif0 g181 (.A(w330), .nZ(w321), .nE(w1597) );
	vdp_notif0 g182 (.A(w331), .nZ(AD_DATA[3]), .nE(w400) );
	vdp_notif0 g183 (.A(w327), .nZ(w288), .nE(w399) );
	vdp_notif0 g184 (.A(w326), .nZ(w321), .nE(w1456) );
	vdp_notif0 g185 (.A(w329), .nZ(AD_DATA[3]), .nE(w414) );
	vdp_notif0 g186 (.A(w283), .nZ(w288), .nE(w392) );
	vdp_notif0 g187 (.A(w282), .nZ(AD_DATA[3]), .nE(w412) );
	vdp_notif0 g188 (.A(w324), .nZ(DB[3]), .nE(w1595) );
	vdp_notif0 g189 (.nZ(DB[11]), .nE(w393), .A(w6772) );
	vdp_notif0 g190 (.A(w325), .nZ(w321), .nE(w1596) );
	vdp_notif0 g191 (.A(w319), .nZ(DB[11]), .nE(w1594) );
	vdp_notif0 g192 (.A(w323), .nZ(DB[3]), .nE(w394) );
	vdp_aon22 g193 (.Z(w323), .A1(w1521), .A2(w1558), .B1(w398), .B2(w319) );
	vdp_aon22 g194 (.A2(w396), .B1(w397), .B2(AD_DATA[3]), .A1(w321), .Z(w280) );
	vdp_aon22 g195 (.A2(w6675), .B1(w6676), .B2(w321), .A1(AD_DATA[3]), .Z(w281) );
	vdp_aon22 g196 (.Z(w282), .A2(w395), .B1(w1559), .B2(w283), .A1(w325) );
	vdp_aon22 g197 (.Z(w329), .A2(w419), .B1(w418), .B2(w326), .A1(w327) );
	vdp_aon22 g198 (.Z(w331), .A2(w426), .B1(w427), .B2(w330), .A1(w332) );
	vdp_aon22 g199 (.Z(w285), .A2(w6671), .B1(w6672), .B2(w286), .A1(w333) );
	vdp_aon22 g200 (.Z(w287), .A1(DB[11]), .A2(w366), .B1(w370), .B2(DB[3]) );
	vdp_slatch g201 (.nQ(w191), .D(VPOS[2]), .C(w1556), .nC(w1557) );
	vdp_slatch g202 (.nQ(w1561), .D(HPOS[3]), .C(w372), .nC(w373) );
	vdp_slatch g203 (.nQ(w193), .D(w244), .C(w1458), .nC(w374) );
	vdp_slatch g204 (.D(w1459), .C(w1554), .nC(w1555), .nQ(w6773) );
	vdp_slatch g205 (.nQ(w194), .D(w197), .C(w1552), .nC(w1553) );
	vdp_slatch g206 (.nQ(w247), .D(w248), .C(w1550), .nC(w1551) );
	vdp_slatch g207 (.nQ(w195), .D(w197), .C(w375), .nC(w376) );
	vdp_slatch g208 (.nQ(w198), .D(w248), .C(w377), .nC(w378) );
	vdp_slatch g209 (.nQ(w199), .D(w197), .C(w425), .nC(w1455) );
	vdp_slatch g210 (.nQ(w201), .D(w248), .C(w1454), .nC(w383) );
	vdp_slatch g211 (.nQ(w202), .D(w197), .C(w381), .nC(w380) );
	vdp_slatch g212 (.nQ(w250), .D(w248), .C(w379), .nC(w1453) );
	vdp_slatch g213 (.Q(w248), .D(DB[2]), .C(w365), .nC(w364) );
	vdp_slatch g214 (.Q(w197), .D(w251), .C(w368), .nC(w367) );
	vdp_sr_bit g215 (.D(w245), .Q(FIFOo[2]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g216 (.A(w203), .nZ(DB[2]), .nE(w1452) );
	vdp_notif0 g217 (.A(w250), .nZ(w245), .nE(w2011) );
	vdp_notif0 g218 (.A(w202), .nZ(RD_DATA[2]), .nE(w382) );
	vdp_notif0 g219 (.A(w249), .nZ(AD_DATA[2]), .nE(w1598) );
	vdp_notif0 g220 (.A(w201), .nZ(w245), .nE(w1549) );
	vdp_notif0 g221 (.A(w199), .nZ(RD_DATA[2]), .nE(w1597) );
	vdp_notif0 g222 (.A(w200), .nZ(AD_DATA[2]), .nE(w400) );
	vdp_notif0 g223 (.A(w198), .nZ(w245), .nE(w399) );
	vdp_notif0 g224 (.A(w195), .nZ(RD_DATA[2]), .nE(w1456) );
	vdp_notif0 g225 (.A(w196), .nZ(AD_DATA[2]), .nE(w414) );
	vdp_notif0 g226 (.A(w247), .nZ(w245), .nE(w392) );
	vdp_notif0 g227 (.A(w246), .nZ(AD_DATA[2]), .nE(w412) );
	vdp_notif0 g228 (.A(w193), .nZ(DB[2]), .nE(w1595) );
	vdp_notif0 g229 (.nZ(DB[10]), .nE(w393), .A(w6773) );
	vdp_notif0 g230 (.A(w194), .nZ(RD_DATA[2]), .nE(w1596) );
	vdp_notif0 g231 (.A(w191), .nZ(DB[10]), .nE(w1594) );
	vdp_notif0 g232 (.A(w192), .nZ(DB[2]), .nE(w394) );
	vdp_aon22 g233 (.A2(w1558), .B1(w398), .B2(w191), .A1(w1561), .Z(w192) );
	vdp_aon22 g234 (.Z(w244), .A2(w396), .B1(w397), .B2(AD_DATA[2]), .A1(RD_DATA[2]) );
	vdp_aon22 g235 (.Z(w1459), .A2(w6675), .B1(w6676), .B2(RD_DATA[2]), .A1(AD_DATA[2]) );
	vdp_aon22 g236 (.Z(w246), .A2(w395), .B1(w1559), .B2(w247), .A1(w194) );
	vdp_aon22 g237 (.Z(w196), .A2(w419), .B1(w418), .B2(w198), .A1(w195) );
	vdp_aon22 g238 (.Z(w200), .A2(w426), .B1(w427), .B2(w201), .A1(w199) );
	vdp_aon22 g239 (.Z(w249), .A2(w6671), .B1(w6672), .B2(w250), .A1(w202) );
	vdp_aon22 g240 (.Z(w251), .A1(DB[10]), .A2(w366), .B1(w370), .B2(DB[2]) );
	vdp_slatch g241 (.nQ(w306), .D(VPOS[1]), .C(w1556), .nC(w1557) );
	vdp_slatch g242 (.nQ(w1522), .D(HPOS[2]), .C(w372), .nC(w373) );
	vdp_slatch g243 (.nQ(w309), .D(w270), .C(w1458), .nC(w374) );
	vdp_slatch g244 (.D(w271), .C(w1554), .nC(w1555), .nQ(w6774) );
	vdp_slatch g245 (.nQ(w310), .D(w313), .C(w1552), .nC(w1553) );
	vdp_slatch g246 (.nQ(w273), .D(w274), .C(w1550), .nC(w1551) );
	vdp_slatch g247 (.nQ(w312), .D(w313), .C(w375), .nC(w376) );
	vdp_slatch g248 (.nQ(w311), .D(w274), .C(w377), .nC(w378) );
	vdp_slatch g249 (.nQ(w315), .D(w313), .C(w425), .nC(w1455) );
	vdp_slatch g250 (.nQ(w317), .D(w274), .C(w1454), .nC(w383) );
	vdp_slatch g251 (.nQ(w318), .D(w313), .C(w381), .nC(w380) );
	vdp_slatch g252 (.nQ(w276), .D(w274), .C(w379), .nC(w1453) );
	vdp_slatch g253 (.Q(w274), .D(DB[1]), .C(w365), .nC(w364) );
	vdp_slatch g254 (.Q(w313), .D(w278), .C(w368), .nC(w367) );
	vdp_sr_bit g255 (.D(w279), .Q(FIFOo[1]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g256 (.A(w1599), .nZ(DB[1]), .nE(w1452) );
	vdp_notif0 g257 (.A(w276), .nZ(w279), .nE(w2011) );
	vdp_notif0 g258 (.A(w318), .nZ(RD_DATA[1]), .nE(w382) );
	vdp_notif0 g259 (.A(w275), .nZ(AD_DATA[1]), .nE(w1598) );
	vdp_notif0 g260 (.A(w317), .nZ(w279), .nE(w1549) );
	vdp_notif0 g261 (.A(w315), .nZ(RD_DATA[1]), .nE(w1597) );
	vdp_notif0 g262 (.A(w316), .nZ(AD_DATA[1]), .nE(w400) );
	vdp_notif0 g263 (.A(w311), .nZ(w279), .nE(w399) );
	vdp_notif0 g264 (.A(w312), .nZ(RD_DATA[1]), .nE(w1456) );
	vdp_notif0 g265 (.A(w314), .nZ(AD_DATA[1]), .nE(w414) );
	vdp_notif0 g266 (.A(w273), .nZ(w279), .nE(w392) );
	vdp_notif0 g267 (.A(w272), .nZ(AD_DATA[1]), .nE(w412) );
	vdp_notif0 g268 (.A(w309), .nZ(DB[1]), .nE(w1595) );
	vdp_notif0 g269 (.nZ(DB[9]), .nE(w393), .A(w6774) );
	vdp_notif0 g270 (.A(w310), .nZ(RD_DATA[1]), .nE(w1596) );
	vdp_notif0 g271 (.A(w306), .nZ(DB[9]), .nE(w1594) );
	vdp_notif0 g272 (.A(w1457), .nZ(DB[1]), .nE(w394) );
	vdp_aon22 g273 (.Z(w1457), .A1(w1522), .A2(w1558), .B1(w398), .B2(w306) );
	vdp_aon22 g274 (.A2(w396), .B1(w397), .B2(AD_DATA[1]), .A1(RD_DATA[1]), .Z(w270) );
	vdp_aon22 g275 (.A2(w6675), .B1(w6676), .B2(RD_DATA[1]), .A1(AD_DATA[1]), .Z(w271) );
	vdp_aon22 g276 (.Z(w272), .A2(w395), .B1(w1559), .B2(w273), .A1(w310) );
	vdp_aon22 g277 (.Z(w314), .A2(w419), .B1(w418), .B2(w312), .A1(w311) );
	vdp_aon22 g278 (.Z(w316), .A2(w426), .B1(w427), .B2(w315), .A1(w317) );
	vdp_aon22 g279 (.Z(w275), .A2(w6671), .B1(w6672), .B2(w276), .A1(w318) );
	vdp_aon22 g280 (.Z(w278), .A1(DB[9]), .A2(w366), .B1(w370), .B2(DB[1]) );
	vdp_slatch g281 (.nQ(w176), .D(w174), .C(w1556), .nC(w1557) );
	vdp_slatch g282 (.D(HPOS[1]), .nQ(w1451), .C(w372), .nC(w373) );
	vdp_slatch g283 (.nQ(w178), .D(w236), .C(w1458), .nC(w374) );
	vdp_slatch g284 (.D(w1426), .C(w1554), .nC(w1555), .nQ(w6775) );
	vdp_slatch g285 (.nQ(w179), .D(w183), .C(w1552), .nC(w1553) );
	vdp_slatch g286 (.nQ(w239), .D(w240), .C(w1550), .nC(w1551) );
	vdp_slatch g287 (.nQ(w180), .D(w183), .C(w375), .nC(w376) );
	vdp_slatch g288 (.nQ(w182), .D(w240), .C(w377), .nC(w378) );
	vdp_slatch g289 (.nQ(w184), .D(w183), .C(w425), .nC(w1455) );
	vdp_slatch g290 (.nQ(w186), .D(w240), .C(w1454), .nC(w383) );
	vdp_slatch g291 (.nQ(w187), .D(w183), .C(w381), .nC(w380) );
	vdp_slatch g292 (.nQ(w242), .D(w240), .C(w379), .nC(w1453) );
	vdp_slatch g293 (.Q(w240), .D(DB[0]), .C(w365), .nC(w364) );
	vdp_slatch g294 (.D(w243), .Q(w183), .C(w368), .nC(w367) );
	vdp_sr_bit g295 (.D(w237), .C2(HCLK2), .C1(HCLK1), .Q(FIFOo[0]), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g296 (.A(1'b1), .nZ(DB[0]), .nE(w1452) );
	vdp_notif0 g297 (.A(w242), .nZ(w237), .nE(w2011) );
	vdp_notif0 g298 (.A(w187), .nZ(RD_DATA[0]), .nE(w382) );
	vdp_notif0 g299 (.A(w241), .nZ(AD_DATA[0]), .nE(w1598) );
	vdp_notif0 g300 (.A(w186), .nZ(w237), .nE(w1549) );
	vdp_notif0 g301 (.A(w184), .nZ(RD_DATA[0]), .nE(w1597) );
	vdp_notif0 g302 (.A(w185), .nZ(AD_DATA[0]), .nE(w400) );
	vdp_notif0 g303 (.A(w182), .nZ(w237), .nE(w399) );
	vdp_notif0 g304 (.A(w180), .nZ(RD_DATA[0]), .nE(w1456) );
	vdp_notif0 g305 (.A(w181), .nZ(AD_DATA[0]), .nE(w414) );
	vdp_notif0 g306 (.A(w239), .nZ(w237), .nE(w392) );
	vdp_notif0 g307 (.A(w238), .nZ(AD_DATA[0]), .nE(w412) );
	vdp_notif0 g308 (.A(w178), .nZ(DB[0]), .nE(w1595) );
	vdp_notif0 g309 (.nZ(DB[8]), .nE(w393), .A(w6775) );
	vdp_notif0 g310 (.A(w179), .nZ(RD_DATA[0]), .nE(w1596) );
	vdp_notif0 g311 (.A(w176), .nZ(DB[8]), .nE(w1594) );
	vdp_notif0 g312 (.A(w177), .nZ(DB[0]), .nE(w394) );
	vdp_aon22 g313 (.A2(w1558), .B1(w398), .B2(w176), .A1(w1451), .Z(w177) );
	vdp_aon22 g314 (.Z(w236), .A2(w396), .B1(w397), .B2(AD_DATA[0]), .A1(RD_DATA[0]) );
	vdp_aon22 g315 (.Z(w1426), .A2(w6675), .B1(w6676), .B2(RD_DATA[0]), .A1(AD_DATA[0]) );
	vdp_aon22 g316 (.Z(w238), .A2(w395), .B1(w1559), .B2(w239), .A1(w179) );
	vdp_aon22 g317 (.Z(w181), .A2(w419), .B1(w418), .B2(w182), .A1(w180) );
	vdp_aon22 g318 (.Z(w185), .A2(w426), .B1(w427), .B2(w186), .A1(w184) );
	vdp_aon22 g319 (.Z(w241), .A2(w6671), .B1(w6672), .B2(w242), .A1(w187) );
	vdp_aon22 g320 (.Z(w243), .A1(DB[8]), .A2(w366), .B1(w370), .B2(DB[0]) );
	vdp_not g321 (.A(w277), .nZ(w1599) );
	vdp_not g322 (.A(w252), .nZ(w203) );
	vdp_not g323 (.A(w402), .nZ(w1594) );
	vdp_not g324 (.A(w406), .nZ(w394) );
	vdp_not g325 (.A(w411), .nZ(w1595) );
	vdp_not g326 (.A(w411), .nZ(w393) );
	vdp_sr_bit g327 (.D(w410), .C2(HCLK2), .C1(HCLK1), .Q(w942), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g328 (.D(w455), .Q(w424), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g329 (.D(w424), .Q(w422), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g330 (.D(w422), .Q(w416), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g331 (.D(w420), .Q(w461), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g332 (.D(w461), .Q(w417), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g333 (.D(w462), .Q(w410), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g334 (.D(w413), .Q(w407), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g335 (.A(w444), .nZ(w1596) );
	vdp_not g336 (.A(w444), .nZ(w412) );
	vdp_not g337 (.A(w444), .nZ(w392) );
	vdp_not g338 (.A(w446), .nZ(w1456) );
	vdp_not g339 (.A(w446), .nZ(w414) );
	vdp_not g340 (.A(w446), .nZ(w399) );
	vdp_not g341 (.A(w458), .nZ(w1597) );
	vdp_not g342 (.A(w458), .nZ(w400) );
	vdp_not g343 (.A(w458), .nZ(w1549) );
	vdp_not g344 (.A(w447), .nZ(w382) );
	vdp_not g345 (.A(w447), .nZ(w1598) );
	vdp_not g346 (.A(w447), .nZ(w2011) );
	vdp_not g347 (.A(w1016), .nZ(w1452) );
	vdp_not g348 (.A(w422), .nZ(w401) );
	vdp_not g349 (.A(w403), .nZ(w404) );
	vdp_comp_str g350 (.A(w437), .Z(w1556), .nZ(w1557) );
	vdp_comp_str g351 (.A(w438), .Z(w372), .nZ(w373) );
	vdp_comp_str g352 (.A(w408), .Z(w1458), .nZ(w374) );
	vdp_comp_str g353 (.A(w409), .Z(w1554), .nZ(w1555) );
	vdp_comp_str g354 (.A(w463), .Z(w1552), .nZ(w1553) );
	vdp_comp_str g355 (.A(w463), .Z(w1550), .nZ(w1551) );
	vdp_comp_str g356 (.A(w460), .Z(w375), .nZ(w376) );
	vdp_comp_str g357 (.A(w460), .Z(w377), .nZ(w378) );
	vdp_comp_str g358 (.A(w504), .Z(w425), .nZ(w1455) );
	vdp_comp_str g359 (.A(w504), .Z(w1454), .nZ(w383) );
	vdp_comp_str g360 (.A(w454), .Z(w381), .nZ(w380) );
	vdp_comp_str g361 (.A(w454), .Z(w379), .nZ(w1453) );
	vdp_comp_str g362 (.A(w465), .Z(w365), .nZ(w364) );
	vdp_comp_str g363 (.A(w465), .Z(w368), .nZ(w367) );
	vdp_comp_we g364 (.A(w403), .Z(w366), .nZ(w370) );
	vdp_comp_we g365 (.A(w443), .Z(w6671), .nZ(w6672) );
	vdp_comp_we g366 (.A(w443), .Z(w426), .nZ(w427) );
	vdp_comp_we g367 (.A(w443), .Z(w419), .nZ(w418) );
	vdp_comp_we g368 (.A(w443), .Z(w395), .nZ(w1559) );
	vdp_comp_we g369 (.A(w448), .Z(w6675), .nZ(w6676) );
	vdp_comp_we g370 (.A(w405), .Z(w396), .nZ(w397) );
	vdp_comp_we g371 (.A(w441), .Z(w1558), .nZ(w398) );
	vdp_and g372 (.Z(w408), .B(HCLK1), .A(w407) );
	vdp_and g373 (.Z(w409), .B(HCLK1), .A(w410) );
	vdp_and g374 (.Z(w413), .B(w417), .A(w415) );
	vdp_and g375 (.Z(w462), .B(w417), .A(w421) );
	vdp_nand g376 (.Z(w421), .B(w448), .A(w401) );
	vdp_nand g377 (.Z(w415), .B(w448), .A(w422) );
	vdp_and3 g378 (.Z(w448), .B(w434), .A(w403), .C(w435) );
	vdp_and3 g379 (.Z(w405), .B(w404), .A(w416), .C(128k) );
	vdp_not g380 (.A(128k), .nZ(w435) );
	vdp_sr_bit g381 (.D(w432), .C2(HCLK2), .C1(HCLK1), .Q(w431), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g382 (.D(w1435), .Q(w469), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g383 (.D(w1514), .C2(HCLK2), .C1(HCLK1), .Q(w495), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g384 (.A(w496), .nZ(w423) );
	vdp_fa g385 (.SUM(w456), .A(w495), .B(1'b0), .CI(w497) );
	vdp_not g386 (.A(w432), .nZ(w430) );
	vdp_not g387 (.A(M5), .nZ(w468) );
	vdp_not g388 (.A(w440), .nZ(w438) );
	vdp_not g389 (.A(w450), .nZ(w451) );
	vdp_not g390 (.A(w502), .nZ(w453) );
	vdp_not g391 (.A(w495), .nZ(w452) );
	vdp_slatch g392 (.Q(w489), .D(w493), .C(w475), .nC(w429) );
	vdp_slatch g393 (.Q(w1502), .D(w493), .C(w487), .nC(w459) );
	vdp_slatch g394 (.Q(w490), .D(w493), .C(w473), .nC(w445) );
	vdp_slatch g395 (.Q(w491), .D(w493), .C(w471), .nC(w442) );
	vdp_slatch g396 (.Q(w492), .D(w466), .C(w475), .nC(w429) );
	vdp_slatch g397 (.Q(w494), .D(w466), .C(w487), .nC(w459) );
	vdp_slatch g398 (.Q(w1501), .D(w466), .E(w473), .nE(w445) );
	vdp_slatch g399 (.Q(w488), .D(w466), .C(w471), .nC(w442) );
	vdp_slatch g400 (.Q(w480), .D(w467), .C(w475), .nC(w429) );
	vdp_slatch g401 (.Q(w474), .D(w467), .C(w487), .nC(w459) );
	vdp_slatch g402 (.Q(w478), .D(w467), .C(w473), .nC(w445) );
	vdp_slatch g403 (.Q(w481), .D(w467), .C(w471), .nC(w442) );
	vdp_comp_dff g404 (.D(w436), .C2(HCLK2), .C1(HCLK1), .Q(w432), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and g405 (.Z(w1435), .B(w430), .A(w431) );
	vdp_or g406 (.Z(w437), .B(w468), .A(w438) );
	vdp_or g407 (.Z(w441), .B(CA[0]), .A(w403) );
	vdp_and3 g408 (.Z(w444), .B(w496), .A(w452), .C(w502) );
	vdp_and3 g409 (.Z(w446), .B(w496), .A(w453), .C(w495) );
	vdp_and3 g410 (.Z(w447), .B(w452), .A(w453), .C(w496) );
	vdp_xor g411 (.Z(w449), .B(w500), .A(w499) );
	vdp_aon22 g412 (.Z(w443), .A1(w451), .A2(w500), .B1(w519), .B2(w450) );
	vdp_and3 g413 (.Z(w458), .B(w495), .A(w502), .C(w496) );
	vdp_comp_str g414 (.A(w504), .Z(w475), .nZ(w429) );
	vdp_comp_str g415 (.A(w454), .Z(w471), .nZ(w442) );
	vdp_comp_str g416 (.A(w463), .Z(w473), .nZ(w445) );
	vdp_comp_str g417 (.A(w460), .Z(w487), .nZ(w459) );
	vdp_nand g418 (.Z(w450), .B(w501), .A(w449) );
	vdp_and g419 (.Z(w1514), .B(w498), .A(w456) );
	vdp_aoi21 g420 (.Z(w440), .B(w439), .A1(HCLK1), .A2(w469) );
	vdp_nor g421 (.Z(w439), .B(w472), .A(w468) );
	vdp_nor g422 (.Z(w434), .B(w466), .A(w467) );
	vdp_not g423 (.A(w483), .nZ(w545) );
	vdp_not g424 (.A(w482), .nZ(w549) );
	vdp_nor g425 (.Z(w609), .A(w530), .B(w483) );
	vdp_or g426 (.A(w1434), .Z(w484), .B(w485) );
	vdp_comp_we g427 (.A(w583), .nZ(w476), .Z(w524) );
	vdp_aon22 g428 (.Z(w482), .A1(w524), .A2(w467), .B1(w476), .B2(w486) );
	vdp_aon22 g429 (.Z(w548), .A1(w524), .A2(w509), .B1(w476), .B2(w484) );
	vdp_aon22 g430 (.Z(w539), .A1(w524), .A2(w535), .B1(w476), .B2(w499) );
	vdp_aon22 g431 (.Z(w483), .A1(w524), .A2(w466), .B1(w476), .B2(w531) );
	vdp_aon22 g432 (.Z(w544), .A1(w524), .A2(w529), .B1(w476), .B2(w500) );
	vdp_aon22 g433 (.Z(w530), .A1(w524), .A2(w493), .B1(w476), .B2(w523) );
	vdp_and g434 (.Z(w543), .A(w522), .B(w521) );
	vdp_and g435 (.Z(w479), .A(w522), .B(w502) );
	vdp_and g436 (.Z(w1503), .A(w495), .B(w521) );
	vdp_and g437 (.Z(w477), .A(w495), .B(w502) );
	vdp_and g438 (.Z(w1436), .A(w498), .B(w517) );
	vdp_fa g439 (.SUM(w517), .A(w502), .B(w503), .CO(w497), .CI(w518) );
	vdp_sr_bit g440 (.D(w1436), .C2(HCLK2), .C1(HCLK1), .Q(w502), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g441 (.A(w520), .nZ(w1438) );
	vdp_not g442 (.A(w510), .nZ(w513) );
	vdp_and g443 (.Z(w503), .A(w578), .B(w1438) );
	vdp_and3 g444 (.Z(w460), .B(w511), .A(w510), .C(w514) );
	vdp_and3 g445 (.Z(w504), .B(w511), .A(w510), .C(w512) );
	vdp_xor g446 (.Z(w516), .A(w495), .B(w510) );
	vdp_not g447 (.A(w502), .nZ(w521) );
	vdp_not g448 (.A(w495), .nZ(w522) );
	vdp_not g449 (.A(w501), .nZ(w1437) );
	vdp_and5 g450 (.Z(w38), .A(w546), .B(w539), .C(w550), .D(w549), .E(w483) );
	vdp_and5 g451 (.Z(w37), .A(w546), .B(w544), .C(w550), .D(w549), .E(w483) );
	vdp_aon2222 g452 (.C2(w540), .B2(w538), .A2(w537), .C1(w1503), .B1(w479), .A1(w543), .Z(w485), .D2(w541), .D1(w477) );
	vdp_aon2222 g453 (.C2(w474), .B2(w478), .A2(w481), .C1(w1503), .B1(w479), .A1(w543), .Z(w486), .D2(w480), .D1(w477) );
	vdp_aon2222 g454 (.C2(w1449), .B2(w534), .A2(w1450), .C1(w1503), .B1(w479), .A1(w543), .Z(w499), .D2(w532), .D1(w477) );
	vdp_aon2222 g455 (.C2(w494), .B2(w1501), .A2(w488), .C1(w1503), .B1(w479), .A1(w543), .Z(w531), .D2(w492), .D1(w477) );
	vdp_aon2222 g456 (.C2(w1504), .B2(w528), .A2(w525), .C1(w1503), .B1(w479), .A1(w543), .Z(w500), .D2(w542), .D1(w477) );
	vdp_aon2222 g457 (.C2(w1502), .B2(w490), .A2(w491), .C1(w1503), .B1(w479), .A1(w543), .Z(w523), .D2(w489), .D1(w477) );
	vdp_nor g458 (.Z(w520), .A(w1437), .B(w449) );
	vdp_or g459 (.Z(w465), .B(w507), .A(w969) );
	vdp_cnt_bit g460 (.R(SYSRES), .Q(w510), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2), .CI(w508) );
	vdp_cnt_bit g461 (.R(SYSRES), .Q(w512), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2), .CI(w571), .CO(w508) );
	vdp_not g462 (.A(w512), .nZ(w514) );
	vdp_not g463 (.A(w1439), .nZ(w511) );
	vdp_and3 g464 (.Z(w454), .B(w511), .A(w513), .C(w514) );
	vdp_and3 g465 (.Z(w463), .B(w511), .A(w513), .C(w512) );
	vdp_xor g466 (.Z(w515), .A(w502), .B(w512) );
	vdp_fa g467 (.SUM(w1563), .A(w579), .B(w519), .CO(w518), .CI(1'b0) );
	vdp_and g468 (.Z(w579), .A(w520), .B(w578) );
	vdp_and g469 (.Z(w1448), .A(w498), .B(w1563) );
	vdp_sr_bit g470 (.D(w1448), .C2(HCLK2), .C1(HCLK1), .Q(w519), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g471 (.A(w1446), .nZ(w564) );
	vdp_comp_str g472 (.A(w454), .Z(w558), .nZ(w536) );
	vdp_comp_str g473 (.A(w463), .Z(w566), .nZ(w526) );
	vdp_comp_str g474 (.A(w460), .Z(w565), .nZ(w533) );
	vdp_comp_str g475 (.A(w504), .Z(w567), .nZ(w527) );
	vdp_slatch g476 (.Q(w542), .D(w529), .C(w567), .nC(w527) );
	vdp_slatch g477 (.Q(w1504), .D(w529), .C(w565), .nC(w533) );
	vdp_slatch g478 (.Q(w528), .D(w529), .C(w566), .nC(w526) );
	vdp_slatch g479 (.Q(w525), .D(w529), .C(w558), .nC(w536) );
	vdp_slatch g480 (.Q(w532), .D(w535), .C(w567), .nC(w527) );
	vdp_slatch g481 (.Q(w1449), .D(w535), .C(w565), .nC(w533) );
	vdp_slatch g482 (.Q(w534), .D(w535), .C(w566), .nC(w526) );
	vdp_slatch g483 (.Q(w1450), .D(w535), .C(w558), .nC(w536) );
	vdp_slatch g484 (.Q(w541), .D(w509), .C(w567), .nC(w527) );
	vdp_slatch g485 (.Q(w540), .D(w509), .C(w565), .nC(w533) );
	vdp_slatch g486 (.Q(w538), .D(w509), .C(w566), .nC(w526) );
	vdp_slatch g487 (.Q(w537), .D(w509), .C(w558), .nC(w536) );
	vdp_and5 g488 (.Z(w173), .A(w546), .B(w539), .C(w549), .D(w530), .E(w545) );
	vdp_and5 g489 (.Z(w172), .A(w546), .B(w544), .C(w549), .D(w530), .E(w545) );
	vdp_not g490 (.A(M5), .nZ(w1434) );
	vdp_not g491 (.A(w530), .nZ(w550) );
	vdp_not g492 (.A(w547), .nZ(w546) );
	vdp_oai21 g493 (.A1(w583), .Z(w547), .A2(w578), .B(w548) );
	vdp_and3 g494 (.Z(w569), .B(w578), .A(w501), .C(w519) );
	vdp_nor g495 (.Z(w1447), .A(w568), .B(w519) );
	vdp_nor g496 (.Z(w576), .A(w516), .B(w515) );
	vdp_aoi21 g497 (.A1(DCLK1), .Z(w1439), .A2(w507), .B(w570) );
	vdp_comb1 g498 (.Z(w1446), .A1(w578), .B(w580), .A2(w1447), .C(HCLK1) );
	vdp_not g499 (.A(w556), .nZ(w35) );
	vdp_not g500 (.A(w1506), .nZ(w551) );
	vdp_not g501 (.A(128k), .nZ(w554) );
	vdp_not g502 (.A(w553), .nZ(w128) );
	vdp_not g503 (.A(w1507), .nZ(w129) );
	vdp_not g504 (.A(w1508), .nZ(w552) );
	vdp_not g505 (.A(VRAMA[0]), .nZ(w1509) );
	vdp_not g506 (.A(w560), .nZ(w559) );
	vdp_not g507 (.A(w495), .nZ(w605) );
	vdp_not g508 (.A(w502), .nZ(w607) );
	vdp_not g509 (.A(w581), .nZ(w604) );
	vdp_not g510 (.A(w403), .nZ(w603) );
	vdp_not g511 (.A(128k), .nZ(w1513) );
	vdp_not g512 (.A(w519), .nZ(w599) );
	vdp_not g513 (.A(SYSRES), .nZ(w498) );
	vdp_not g514 (.A(w587), .nZ(w1441) );
	vdp_not g515 (.A(w34), .nZ(w1440) );
	vdp_not g516 (.A(w577), .nZ(w595) );
	vdp_not g517 (.A(w570), .nZ(w574) );
	vdp_not g518 (.A(w574), .nZ(w575) );
	vdp_sr_bit g519 (.D(w1442), .C2(HCLK2), .C1(HCLK1), .Q(w578), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g520 (.D(w1445), .Q(w583), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_slatch g521 (.Q(w455), .D(VRAMA[0]), .C(w595), .nC(w577) );
	vdp_and g522 (.A(w32), .Z(w1442), .B(w1441) );
	vdp_and g523 (.A(w1440), .Z(w496), .B(w3) );
	vdp_and g524 (.A(w3), .Z(w577), .B(HCLK1) );
	vdp_and g525 (.A(w587), .Z(w34), .B(w585) );
	vdp_and g526 (.A(w586), .Z(w36), .B(w587) );
	vdp_and g527 (.A(w586), .B(w569) );
	vdp_or g528 (.A(w573), .Z(w571), .B(w507) );
	vdp_or g529 (.A(w575), .Z(w941), .B(1'b0) );
	vdp_or g530 (.A(SYSRES), .Z(w597), .B(w590) );
	vdp_and g531 (.A(w578), .Z(w1443), .B(DMA_BUSY) );
	vdp_and g532 (.A(w609), .Z(w501), .B(w1512) );
	vdp_and g533 (.A(w1513), .Z(w1512), .B(w403) );
	vdp_or g534 (.A(w569), .Z(w602), .B(w568) );
	vdp_or g535 (.A(DMA_BUSY), .Z(w1510), .B(w563) );
	vdp_or g536 (.A(DMA_BUSY), .Z(w1511), .B(w562) );
	vdp_and g537 (.A(M5), .Z(w581), .B(REG_BUS[0]) );
	vdp_or g538 (.A(w539), .Z(w555), .B(w554) );
	vdp_and g539 (.A(w544), .Z(w1505), .B(128k) );
	vdp_aon22 g540 (.Z(w529), .A2(w1510), .B1(w603), .B2(w581), .A1(w403) );
	vdp_aon22 g541 (.Z(w535), .A2(w1511), .B1(w604), .B2(w603), .A1(w403) );
	vdp_and3 g542 (.A(w32), .Z(w1445), .B(w36), .C(w1444) );
	vdp_rs_ff g543 (.Q(w1444), .R(w597), .S(w1443) );
	vdp_oai21 g544 (.A1(VRAMA[0]), .Z(w560), .A2(128k), .B(w589) );
	vdp_oai21 g545 (.A1(128k), .Z(w1508), .A2(w1509), .B(w589) );
	vdp_aoi21 g546 (.A1(w544), .Z(w1507), .A2(w557), .B(w559) );
	vdp_aoi21 g547 (.A1(w539), .Z(w553), .A2(w557), .B(w552) );
	vdp_aoi21 g548 (.A1(w557), .Z(w1506), .A2(w555), .B(w589) );
	vdp_aoi21 g549 (.A1(w557), .Z(w556), .A2(w1505), .B(w589) );
	vdp_and4 g550 (.A(w546), .Z(w557), .B(w550), .C(w545), .D(w549) );
	vdp_not g551 (.A(w634), .nZ(w1433) );
	vdp_not g552 (.A(w646), .nZ(w645) );
	vdp_and3 g553 (.A(w599), .Z(w600), .B(w636), .C(w645) );
	vdp_and3 g554 (.A(w607), .Z(w623), .B(w610), .C(w605) );
	vdp_and3 g555 (.A(w502), .Z(w627), .B(w610), .C(w605) );
	vdp_and3 g556 (.A(w607), .Z(w616), .B(w610), .C(w495) );
	vdp_and3 g557 (.A(w502), .Z(w620), .B(w610), .C(w495) );
	vdp_or g558 (.A(w601), .Z(w633), .B(w635) );
	vdp_or g559 (.A(w601), .Z(w639), .B(w643) );
	vdp_or g560 (.A(w669), .Z(w588), .B(w642) );
	vdp_and3 g561 (.Z(w586), .B(DMA_BUSY), .A(w668), .C(w641) );
	vdp_or3 g562 (.Z(w592), .B(w583), .A(w589), .C(w640) );
	vdp_and g563 (.A(w593), .Z(w507), .B(w594) );
	vdp_and g564 (.A(w578), .Z(w610), .B(w599) );
	vdp_bufif0 g565 (.A(w591), .Z(VRAMA[8]), .nE(w647) );
	vdp_aoi221 g566 (.Z(w634), .A2(w600), .B1(w587), .B2(w576), .A1(w576), .C(SYSRES) );
	vdp_aon33 g567 (.Z(w1033), .A2(w576), .B1(w1543), .B2(w576), .A1(w644), .A3(w1543), .B3(w596) );
	vdp_not g568 (.A(w602), .nZ(w1461) );
	vdp_comp_str g569 (.A(w564), .Z(w1462), .nZ(w630) );
	vdp_not g570 (.A(w627), .nZ(w629) );
	vdp_comp_str g571 (.A(w463), .Z(w1464), .nZ(w1463) );
	vdp_not g572 (.A(w602), .nZ(w847) );
	vdp_comp_str g573 (.A(w564), .Z(w631), .nZ(w632) );
	vdp_not g574 (.A(w580), .nZ(w647) );
	vdp_not g575 (.A(w627), .nZ(w1544) );
	vdp_comp_str g576 (.A(w463), .Z(w1465), .nZ(w628) );
	vdp_not g577 (.A(w623), .nZ(w622) );
	vdp_comp_str g578 (.A(w454), .Z(w1466), .nZ(w1548) );
	vdp_not g579 (.A(w623), .nZ(w624) );
	vdp_comp_str g580 (.A(w504), .Z(w1467), .nZ(w621) );
	vdp_comp_str g581 (.A(w454), .Z(w625), .nZ(w626) );
	vdp_not g582 (.A(w616), .nZ(w613) );
	vdp_comp_str g583 (.A(w460), .Z(w614), .nZ(w615) );
	vdp_not g584 (.A(w616), .nZ(w846) );
	vdp_comp_str g585 (.A(w460), .Z(w1546), .nZ(w1547) );
	vdp_not g586 (.A(w620), .nZ(w617) );
	vdp_comp_str g587 (.A(w504), .Z(w618), .nZ(w619) );
	vdp_not g588 (.A(w620), .nZ(w1545) );
	vdp_sr_bit g589 (.D(w1433), .Q(w587), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g590 (.D(w636), .Q(w646), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g591 (.D(w578), .Q(w636), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g592 (.D(w1033), .Q(w644), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g593 (.D(w571), .Q(w596), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_not g594 (.A(SYSRES), .nZ(w1543) );
	vdp_not g595 (.A(w1515), .nZ(w640) );
	vdp_sr_bit g596 (.D(w593), .Q(w594), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g597 (.D(w584), .C2(HCLK2), .C1(HCLK1), .Q(w590), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_dlatch_inv g598 (.D(w593), .C(HCLK2), .Q(w1515), .nC(nHCLK2) );
	vdp_slatch g599 (.D(w658), .C(w614), .nC(w615), .nQ(w6691) );
	vdp_slatch g600 (.D(REG_BUS[7]), .C(w1546), .nC(w1547), .nQ(w6692) );
	vdp_slatch g601 (.D(w658), .C(w618), .nC(w619), .nQ(w6711) );
	vdp_slatch g602 (.D(REG_BUS[7]), .C(w1467), .nC(w621), .nQ(w6709) );
	vdp_slatch g603 (.D(w658), .C(w1466), .nC(w1548), .nQ(w6725) );
	vdp_slatch g604 (.D(REG_BUS[7]), .C(w625), .nC(w626), .nQ(w6727) );
	vdp_slatch g605 (.D(w658), .C(w1465), .nC(w628), .nQ(w6745) );
	vdp_slatch g606 (.D(REG_BUS[7]), .C(w1464), .nC(w1463), .nQ(w6743) );
	vdp_slatch g607 (.D(VRAMA[9]), .C(w1462), .nC(w630), .nQ(w6759) );
	vdp_slatch g608 (.D(VRAMA[7]), .C(w631), .nC(w632), .nQ(w6760) );
	vdp_notif0 g609 (.nZ(VRAMA[7]), .nE(w847), .A(w6760) );
	vdp_notif0 g610 (.nZ(VRAMA[9]), .nE(w1461), .A(w6759) );
	vdp_notif0 g611 (.nZ(VRAMA[7]), .nE(w629), .A(w6743) );
	vdp_notif0 g612 (.nZ(VRAMA[9]), .nE(w1544), .A(w6745) );
	vdp_notif0 g613 (.nZ(VRAMA[7]), .nE(w624), .A(w6727) );
	vdp_notif0 g614 (.nZ(VRAMA[9]), .nE(w617), .A(w6711) );
	vdp_notif0 g615 (.nZ(VRAMA[7]), .nE(w1545), .A(w6709) );
	vdp_notif0 g616 (.nZ(VRAMA[9]), .nE(w622), .A(w6725) );
	vdp_notif0 g617 (.nZ(VRAMA[9]), .nE(w613), .A(w6691) );
	vdp_notif0 g618 (.nZ(VRAMA[7]), .nE(w846), .A(w6692) );
	vdp_bufif0 g619 (.A(w658), .Z(VRAMA[9]), .nE(w647) );
	vdp_bufif0 g620 (.A(REG_BUS[7]), .Z(VRAMA[7]), .nE(w647) );
	vdp_bufif0 g621 (.A(w651), .Z(VRAMA[8]), .nE(w1497) );
	vdp_bufif0 g622 (.A(w651), .Z(CA[8]), .nE(w849) );
	vdp_bufif0 g623 (.A(w650), .Z(VRAMA[7]), .nE(w1495) );
	vdp_bufif0 g624 (.A(w650), .Z(CA[7]), .nE(w848) );
	vdp_slatch g625 (.Q(w668), .D(REG_BUS[7]), .nQ(w665), .C(w1589), .nC(w1590) );
	vdp_not g626 (.A(REG_BUS[0]), .nZ(w663) );
	vdp_not g627 (.A(REG_BUS[7]), .nZ(w670) );
	vdp_and3 g628 (.Z(w669), .B(w641), .A(w665), .C(DMA_BUSY) );
	vdp_nand g629 (.A(w661), .Z(w690), .B(w662) );
	vdp_cnt_bit_load g630 (.D(REG_BUS[0]), .nL(w1592), .L(w1601), .R(1'b0), .Q(w651), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w633), .CO(w655) );
	vdp_cnt_bit_load g631 (.D(REG_BUS[7]), .nL(w1432), .L(w803), .R(1'b0), .Q(w650), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w653), .CO(w635) );
	vdp_cnt_bit_load g632 (.D(w663), .nL(w1591), .L(w812), .R(1'b0), .Q(w661), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w639), .CO(w660) );
	vdp_cnt_bit_load g633 (.D(w670), .nL(w793), .L(w794), .R(1'b0), .Q(w664), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w666), .CO(w643) );
	vdp_slatch g634 (.D(w678), .C(w614), .nC(w615), .nQ(w6690) );
	vdp_slatch g635 (.D(REG_BUS[6]), .C(w1546), .nC(w1547), .nQ(w6693) );
	vdp_slatch g636 (.D(w678), .C(w618), .nC(w619), .nQ(w6710) );
	vdp_slatch g637 (.D(REG_BUS[6]), .C(w1467), .nC(w621), .nQ(w6708) );
	vdp_slatch g638 (.D(w678), .C(w1466), .nC(w1548), .nQ(w6724) );
	vdp_slatch g639 (.D(REG_BUS[6]), .C(w625), .nC(w626), .nQ(w6726) );
	vdp_slatch g640 (.D(w678), .C(w1465), .nC(w628), .nQ(w6744) );
	vdp_slatch g641 (.D(REG_BUS[6]), .C(w1464), .nC(w1463), .nQ(w6742) );
	vdp_slatch g642 (.D(VRAMA[10]), .C(w1462), .nC(w630), .nQ(w6758) );
	vdp_slatch g643 (.D(VRAMA[6]), .C(w631), .nC(w632), .nQ(w6761) );
	vdp_notif0 g644 (.nZ(VRAMA[6]), .nE(w847), .A(w6761) );
	vdp_notif0 g645 (.nZ(VRAMA[10]), .nE(w1461), .A(w6758) );
	vdp_notif0 g646 (.nZ(VRAMA[6]), .nE(w629), .A(w6742) );
	vdp_notif0 g647 (.nZ(VRAMA[10]), .nE(w1544), .A(w6744) );
	vdp_notif0 g648 (.nZ(VRAMA[6]), .nE(w624), .A(w6726) );
	vdp_notif0 g649 (.nZ(VRAMA[10]), .nE(w617), .A(w6710) );
	vdp_notif0 g650 (.nZ(VRAMA[6]), .nE(w1545), .A(w6708) );
	vdp_notif0 g651 (.nZ(VRAMA[10]), .nE(w622), .A(w6724) );
	vdp_notif0 g652 (.nZ(VRAMA[10]), .nE(w613), .A(w6690) );
	vdp_notif0 g653 (.nZ(VRAMA[6]), .nE(w846), .A(w6693) );
	vdp_bufif0 g654 (.A(w678), .Z(VRAMA[10]), .nE(w647) );
	vdp_bufif0 g655 (.A(REG_BUS[6]), .Z(VRAMA[6]), .nE(w1498) );
	vdp_bufif0 g656 (.A(w649), .Z(VRAMA[9]), .nE(w1497) );
	vdp_bufif0 g657 (.A(w649), .Z(CA[9]), .nE(w849) );
	vdp_bufif0 g658 (.A(w672), .Z(VRAMA[6]), .nE(w1495) );
	vdp_bufif0 g659 (.A(w672), .Z(CA[6]), .nE(w848) );
	vdp_slatch g660 (.Q(w685), .D(REG_BUS[6]), .nQ(w641), .C(w1589), .nC(w1590) );
	vdp_not g661 (.A(REG_BUS[1]), .nZ(w681) );
	vdp_not g662 (.A(REG_BUS[6]), .nZ(w683) );
	vdp_and3 g663 (.Z(w642), .B(DMA_BUSY), .A(w685), .C(w665) );
	vdp_cnt_bit_load g664 (.D(REG_BUS[1]), .nL(w1592), .L(w1601), .R(1'b0), .Q(w649), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w655), .CO(w674) );
	vdp_cnt_bit_load g665 (.D(REG_BUS[6]), .nL(w1432), .L(w803), .R(1'b0), .Q(w672), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w673), .CO(w653) );
	vdp_cnt_bit_load g666 (.D(w681), .nL(w1591), .L(w812), .R(1'b0), .Q(w662), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w660), .CO(w680) );
	vdp_cnt_bit_load g667 (.D(w683), .nL(w793), .L(w794), .R(1'b0), .Q(w682), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w686), .CO(w666) );
	vdp_nand3 g668 (.Z(w689), .B(w682), .A(w688), .C(w664) );
	vdp_slatch g669 (.D(w702), .C(w614), .nC(w615), .nQ(w6689) );
	vdp_slatch g670 (.D(REG_BUS[5]), .C(w1546), .nC(w1547), .nQ(w6694) );
	vdp_slatch g671 (.D(w702), .C(w618), .nC(w619), .nQ(w6712) );
	vdp_slatch g672 (.D(REG_BUS[5]), .C(w1467), .nC(w621), .nQ(w6707) );
	vdp_slatch g673 (.D(w702), .C(w1466), .nC(w1548), .nQ(w6723) );
	vdp_slatch g674 (.D(w702), .C(w1465), .nC(w628), .nQ(w6746) );
	vdp_slatch g675 (.D(REG_BUS[5]), .C(w1464), .nC(w1463), .nQ(w6741) );
	vdp_slatch g676 (.D(VRAMA[11]), .C(w1462), .nC(w630), .nQ(w6757) );
	vdp_slatch g677 (.D(VRAMA[5]), .C(w631), .nC(w632), .nQ(w6762) );
	vdp_notif0 g678 (.nZ(VRAMA[5]), .nE(w847), .A(w6762) );
	vdp_notif0 g679 (.nZ(VRAMA[11]), .nE(w1461), .A(w6757) );
	vdp_notif0 g680 (.nZ(VRAMA[5]), .nE(w629), .A(w6741) );
	vdp_notif0 g681 (.nZ(VRAMA[11]), .nE(w1544), .A(w6746) );
	vdp_notif0 g682 (.nZ(VRAMA[5]), .nE(w624), .A(w6728) );
	vdp_notif0 g683 (.nZ(VRAMA[11]), .nE(w617), .A(w6712) );
	vdp_notif0 g684 (.nZ(VRAMA[5]), .nE(w1545), .A(w6707) );
	vdp_notif0 g685 (.nZ(VRAMA[11]), .nE(w622), .A(w6723) );
	vdp_notif0 g686 (.nZ(VRAMA[11]), .nE(w613), .A(w6689) );
	vdp_notif0 g687 (.nZ(VRAMA[5]), .nE(w846), .A(w6694) );
	vdp_bufif0 g688 (.A(w702), .Z(VRAMA[11]), .nE(w647) );
	vdp_bufif0 g689 (.A(REG_BUS[5]), .Z(VRAMA[5]), .nE(w1498) );
	vdp_bufif0 g690 (.A(w671), .Z(VRAMA[10]), .nE(w1497) );
	vdp_bufif0 g691 (.A(w671), .Z(CA[10]), .nE(w849) );
	vdp_bufif0 g692 (.A(w704), .Z(VRAMA[5]), .nE(w1495) );
	vdp_bufif0 g693 (.A(w704), .Z(CA[5]), .nE(w848) );
	vdp_slatch g694 (.Q(CA[18]), .D(REG_BUS[2]), .C(w1589), .nC(w1590) );
	vdp_not g695 (.A(REG_BUS[2]), .nZ(w697) );
	vdp_not g696 (.A(REG_BUS[5]), .nZ(w696) );
	vdp_and3 g697 (.Z(w585), .B(DMA_BUSY), .A(w685), .C(w668) );
	vdp_cnt_bit_load g698 (.D(REG_BUS[2]), .nL(w1592), .L(w1601), .R(1'b0), .Q(w671), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w674), .CO(w707) );
	vdp_cnt_bit_load g699 (.D(REG_BUS[5]), .nL(w1432), .L(w803), .R(1'b0), .Q(w704), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w703), .CO(w673) );
	vdp_cnt_bit_load g700 (.D(w697), .nL(w1591), .L(w812), .R(1'b0), .Q(w687), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w680), .CO(w698) );
	vdp_cnt_bit_load g701 (.D(w696), .nL(w793), .L(w794), .R(1'b0), .Q(w688), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w693), .CO(w686) );
	vdp_nand3 g702 (.Z(w701), .B(w699), .A(w700), .C(w687) );
	vdp_slatch g703 (.D(w716), .C(w614), .nC(w615), .nQ(w6688) );
	vdp_slatch g704 (.D(REG_BUS[4]), .C(w1546), .nC(w1547), .nQ(w6695) );
	vdp_slatch g705 (.D(w716), .C(w618), .nC(w619), .nQ(w6713) );
	vdp_slatch g706 (.D(REG_BUS[4]), .C(w1467), .nC(w621), .nQ(w6706) );
	vdp_slatch g707 (.D(w716), .C(w1466), .nC(w1548), .nQ(w6722) );
	vdp_slatch g708 (.D(w716), .C(w1465), .nC(w628), .nQ(w6747) );
	vdp_slatch g709 (.D(REG_BUS[4]), .C(w1464), .nC(w1463), .nQ(w6740) );
	vdp_slatch g710 (.D(VRAMA[12]), .C(w1462), .nC(w630), .nQ(w6756) );
	vdp_slatch g711 (.D(VRAMA[4]), .C(w631), .nC(w632), .nQ(w6763) );
	vdp_notif0 g712 (.nZ(VRAMA[4]), .nE(w847), .A(w6763) );
	vdp_notif0 g713 (.nZ(VRAMA[12]), .nE(w1461), .A(w6756) );
	vdp_notif0 g714 (.nZ(VRAMA[4]), .nE(w629), .A(w6740) );
	vdp_notif0 g715 (.nZ(VRAMA[12]), .nE(w1544), .A(w6747) );
	vdp_notif0 g716 (.nZ(VRAMA[4]), .nE(w624), .A(w6729) );
	vdp_notif0 g717 (.nZ(VRAMA[12]), .nE(w617), .A(w6713) );
	vdp_notif0 g718 (.nZ(VRAMA[4]), .nE(w1545), .A(w6706) );
	vdp_notif0 g719 (.nZ(VRAMA[12]), .nE(w622), .A(w6722) );
	vdp_notif0 g720 (.nZ(VRAMA[12]), .nE(w613), .A(w6688) );
	vdp_notif0 g721 (.nZ(VRAMA[4]), .nE(w846), .A(w6695) );
	vdp_bufif0 g722 (.A(w716), .Z(VRAMA[12]), .nE(w647) );
	vdp_bufif0 g723 (.A(REG_BUS[4]), .Z(VRAMA[4]), .nE(w1498) );
	vdp_bufif0 g724 (.A(w706), .Z(VRAMA[11]), .nE(w1497) );
	vdp_bufif0 g725 (.A(w706), .Z(CA[11]), .nE(w849) );
	vdp_bufif0 g726 (.A(w717), .Z(VRAMA[4]), .nE(w1495) );
	vdp_bufif0 g727 (.A(w717), .Z(CA[4]), .nE(w848) );
	vdp_slatch g728 (.Q(CA[19]), .D(REG_BUS[3]), .C(w1589), .nC(w1590) );
	vdp_not g729 (.A(REG_BUS[3]), .nZ(w718) );
	vdp_not g730 (.A(REG_BUS[4]), .nZ(w720) );
	vdp_and g731 (.Z(w584), .B(w695), .A(w728) );
	vdp_cnt_bit_load g732 (.D(REG_BUS[3]), .nL(w1592), .L(w1601), .R(1'b0), .Q(w706), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w707), .CO(w712) );
	vdp_cnt_bit_load g733 (.D(REG_BUS[4]), .nL(w1432), .L(w803), .R(1'b0), .Q(w717), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w722), .CO(w703) );
	vdp_cnt_bit_load g734 (.D(w718), .nL(w1591), .L(w812), .R(1'b0), .Q(w699), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w698), .CO(w723) );
	vdp_cnt_bit_load g735 (.D(w720), .nL(w793), .L(w794), .R(1'b0), .Q(w726), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w727), .CO(w693) );
	vdp_nor3 g736 (.Z(w695), .B(w701), .A(w725), .C(w690) );
	vdp_slatch g737 (.D(w734), .C(w614), .nC(w615), .nQ(w6687) );
	vdp_slatch g738 (.D(REG_BUS[3]), .C(w1546), .nC(w1547), .nQ(w6696) );
	vdp_slatch g739 (.D(w734), .C(w618), .nC(w619), .nQ(w6714) );
	vdp_slatch g740 (.D(REG_BUS[3]), .C(w1467), .nC(w621), .nQ(w6705) );
	vdp_slatch g741 (.D(w734), .C(w1466), .nC(w1548), .nQ(w6721) );
	vdp_slatch g742 (.D(REG_BUS[3]), .C(w625), .nC(w626), .nQ(w6731) );
	vdp_slatch g743 (.D(w734), .C(w1465), .nC(w628), .nQ(w6749) );
	vdp_slatch g744 (.D(REG_BUS[3]), .C(w1464), .nC(w1463), .nQ(w6739) );
	vdp_slatch g745 (.D(VRAMA[13]), .C(w1462), .nC(w630), .nQ(w6755) );
	vdp_slatch g746 (.D(VRAMA[3]), .C(w631), .nC(w632), .nQ(w6764) );
	vdp_notif0 g747 (.nZ(VRAMA[3]), .nE(w847), .A(w6764) );
	vdp_notif0 g748 (.nZ(VRAMA[13]), .nE(w1461), .A(w6755) );
	vdp_notif0 g749 (.nZ(VRAMA[3]), .nE(w629), .A(w6739) );
	vdp_notif0 g750 (.nZ(VRAMA[13]), .nE(w1544), .A(w6749) );
	vdp_notif0 g751 (.nZ(VRAMA[3]), .nE(w624), .A(w6731) );
	vdp_notif0 g752 (.nZ(VRAMA[13]), .nE(w617), .A(w6714) );
	vdp_notif0 g753 (.nZ(VRAMA[3]), .nE(w1545), .A(w6705) );
	vdp_notif0 g754 (.nZ(VRAMA[13]), .nE(w622), .A(w6721) );
	vdp_notif0 g755 (.nZ(VRAMA[13]), .nE(w613), .A(w6687) );
	vdp_notif0 g756 (.nZ(VRAMA[3]), .nE(w846), .A(w6696) );
	vdp_bufif0 g757 (.A(w734), .Z(VRAMA[13]), .nE(w647) );
	vdp_bufif0 g758 (.A(REG_BUS[3]), .Z(VRAMA[3]), .nE(w1498) );
	vdp_bufif0 g759 (.A(w711), .Z(VRAMA[12]), .nE(w1497) );
	vdp_bufif0 g760 (.A(w711), .Z(CA[12]), .nE(w849) );
	vdp_bufif0 g761 (.A(w742), .Z(VRAMA[3]), .nE(w1495) );
	vdp_bufif0 g762 (.A(w742), .Z(CA[3]), .nE(w848) );
	vdp_slatch g763 (.Q(w749), .D(REG_BUS[4]), .C(w1589), .nC(w1590) );
	vdp_not g764 (.A(REG_BUS[4]), .nZ(w736) );
	vdp_not g765 (.A(REG_BUS[3]), .nZ(w737) );
	vdp_cnt_bit_load g766 (.D(REG_BUS[4]), .nL(w1592), .L(w1601), .R(1'b0), .Q(w711), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w712), .CO(w733) );
	vdp_cnt_bit_load g767 (.D(REG_BUS[3]), .nL(w1432), .L(w803), .R(1'b0), .Q(w742), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w731), .CO(w722) );
	vdp_cnt_bit_load g768 (.D(w736), .nL(w1591), .L(w812), .R(1'b0), .Q(w700), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w723), .CO(w741) );
	vdp_cnt_bit_load g769 (.D(w737), .nL(w793), .L(w794), .R(1'b0), .Q(w746), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w738), .CO(w727) );
	vdp_nor3 g770 (.Z(w728), .B(w747), .A(w745), .C(w689) );
	vdp_bufif0 g771 (.A(w749), .Z(CA[20]), .nE(w791) );
	vdp_slatch g772 (.D(w753), .C(w614), .nC(w615), .nQ(w6686) );
	vdp_slatch g773 (.D(REG_BUS[2]), .C(w1546), .nC(w1547), .nQ(w6697) );
	vdp_slatch g774 (.D(w753), .C(w618), .nC(w619), .nQ(w6715) );
	vdp_slatch g775 (.D(REG_BUS[2]), .C(w1467), .nC(w621), .nQ(w6704) );
	vdp_slatch g776 (.D(w753), .C(w1466), .nC(w1548), .nQ(w6720) );
	vdp_slatch g777 (.D(REG_BUS[2]), .C(w625), .nC(w626), .nQ(w6730) );
	vdp_slatch g778 (.D(w753), .C(w1465), .nC(w628), .nQ(w6748) );
	vdp_slatch g779 (.D(REG_BUS[2]), .C(w1464), .nC(w1463), .nQ(w6738) );
	vdp_slatch g780 (.D(VRAMA[14]), .C(w1462), .nC(w630), .nQ(w6754) );
	vdp_slatch g781 (.D(VRAMA[2]), .nC(w632), .C(w631), .nQ(w6765) );
	vdp_notif0 g782 (.nZ(VRAMA[2]), .nE(w847), .A(w6765) );
	vdp_notif0 g783 (.nZ(VRAMA[14]), .nE(w1461), .A(w6754) );
	vdp_notif0 g784 (.nZ(VRAMA[2]), .nE(w629), .A(w6738) );
	vdp_notif0 g785 (.nZ(VRAMA[14]), .nE(w1544), .A(w6748) );
	vdp_notif0 g786 (.nZ(VRAMA[2]), .nE(w624), .A(w6730) );
	vdp_notif0 g787 (.nZ(VRAMA[14]), .nE(w617), .A(w6715) );
	vdp_notif0 g788 (.nZ(VRAMA[2]), .nE(w1545), .A(w6704) );
	vdp_notif0 g789 (.nZ(VRAMA[14]), .nE(w622), .A(w6720) );
	vdp_notif0 g790 (.nZ(VRAMA[14]), .nE(w613), .A(w6686) );
	vdp_notif0 g791 (.nZ(VRAMA[2]), .nE(w846), .A(w6697) );
	vdp_bufif0 g792 (.A(w753), .Z(VRAMA[14]), .nE(w1496) );
	vdp_bufif0 g793 (.A(REG_BUS[2]), .Z(VRAMA[2]), .nE(w1498) );
	vdp_bufif0 g794 (.A(w732), .Z(VRAMA[13]), .nE(w1497) );
	vdp_bufif0 g795 (.A(w732), .Z(CA[13]), .nE(w849) );
	vdp_bufif0 g796 (.A(w754), .Z(VRAMA[2]), .nE(w1495) );
	vdp_bufif0 g797 (.A(w754), .Z(CA[2]), .nE(w848) );
	vdp_slatch g798 (.Q(w761), .D(REG_BUS[5]), .C(w1589), .nC(w1590) );
	vdp_not g799 (.A(REG_BUS[5]), .nZ(w755) );
	vdp_not g800 (.A(REG_BUS[2]), .nZ(w756) );
	vdp_cnt_bit_load g801 (.D(REG_BUS[5]), .nL(w1592), .L(w1601), .R(1'b0), .Q(w732), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w733), .CO(w767) );
	vdp_cnt_bit_load g802 (.D(REG_BUS[2]), .nL(w1432), .L(w803), .R(1'b0), .Q(w754), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w766), .CO(w731) );
	vdp_cnt_bit_load g803 (.D(w755), .nL(w1591), .L(w812), .R(1'b0), .Q(w765), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w741), .CO(w757) );
	vdp_cnt_bit_load g804 (.D(w756), .nL(w793), .L(w794), .R(1'b0), .Q(w763), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w769), .CO(w738) );
	vdp_nand3 g805 (.Z(w747), .B(w746), .A(w763), .C(w726) );
	vdp_bufif0 g806 (.A(w761), .Z(CA[21]), .nE(w791) );
	vdp_slatch g807 (.D(w774), .C(w614), .nC(w615), .nQ(w6685) );
	vdp_slatch g808 (.D(REG_BUS[1]), .C(w1546), .nC(w1547), .nQ(w6698) );
	vdp_slatch g809 (.D(w774), .C(w618), .nC(w619), .nQ(w6717) );
	vdp_slatch g810 (.D(REG_BUS[1]), .C(w1467), .nC(w621), .nQ(w6703) );
	vdp_slatch g811 (.D(w774), .C(w1466), .nC(w1548), .nQ(w6719) );
	vdp_slatch g812 (.D(REG_BUS[1]), .C(w625), .nC(w626), .nQ(w6733) );
	vdp_slatch g813 (.D(w774), .C(w1465), .nC(w628), .nQ(w6750) );
	vdp_slatch g814 (.D(REG_BUS[1]), .C(w1464), .nC(w1463), .nQ(w6737) );
	vdp_slatch g815 (.D(VRAMA[15]), .C(w1462), .nC(w630), .nQ(w6753) );
	vdp_slatch g816 (.D(VRAMA[1]), .C(w631), .nC(w632), .nQ(w6766) );
	vdp_notif0 g817 (.nZ(VRAMA[1]), .nE(w847), .A(w6766) );
	vdp_notif0 g818 (.nZ(VRAMA[15]), .nE(w1461), .A(w6753) );
	vdp_notif0 g819 (.nZ(VRAMA[1]), .nE(w629), .A(w6737) );
	vdp_notif0 g820 (.nZ(VRAMA[15]), .nE(w1544), .A(w6750) );
	vdp_notif0 g821 (.nZ(VRAMA[1]), .nE(w624), .A(w6733) );
	vdp_notif0 g822 (.nZ(VRAMA[15]), .nE(w617), .A(w6717) );
	vdp_notif0 g823 (.nZ(VRAMA[1]), .nE(w1545), .A(w6703) );
	vdp_notif0 g824 (.nZ(VRAMA[15]), .nE(w622), .A(w6719) );
	vdp_notif0 g825 (.nZ(VRAMA[15]), .nE(w613), .A(w6685) );
	vdp_notif0 g826 (.nZ(VRAMA[1]), .nE(w846), .A(w6698) );
	vdp_bufif0 g827 (.A(w774), .Z(VRAMA[15]), .nE(w1496) );
	vdp_bufif0 g828 (.A(REG_BUS[1]), .Z(VRAMA[1]), .nE(w1498) );
	vdp_bufif0 g829 (.A(w750), .Z(VRAMA[14]), .nE(w1497) );
	vdp_bufif0 g830 (.A(w750), .Z(CA[14]), .nE(w849) );
	vdp_bufif0 g831 (.A(w776), .Z(VRAMA[1]), .nE(w1495) );
	vdp_bufif0 g832 (.A(w776), .Z(CA[1]), .nE(w848) );
	vdp_slatch g833 (.Q(w1499), .D(REG_BUS[1]), .C(w1589), .nC(w1590) );
	vdp_not g834 (.A(REG_BUS[6]), .nZ(w779) );
	vdp_not g835 (.A(REG_BUS[1]), .nZ(w782) );
	vdp_cnt_bit_load g836 (.D(REG_BUS[6]), .nL(w1592), .L(w1601), .R(1'b0), .Q(w750), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w767), .CO(w783) );
	vdp_cnt_bit_load g837 (.D(REG_BUS[1]), .nL(w1432), .L(w803), .R(1'b0), .Q(w776), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w784), .CO(w766) );
	vdp_cnt_bit_load g838 (.D(w779), .nL(w1591), .L(w812), .R(1'b0), .Q(w764), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w757), .CO(w777) );
	vdp_cnt_bit_load g839 (.D(w782), .nL(w793), .L(w794), .R(1'b0), .Q(w781), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w780), .CO(w769) );
	vdp_nand3 g840 (.Z(w725), .B(w764), .A(w765), .C(w778) );
	vdp_bufif0 g841 (.A(w1499), .Z(CA[17]), .nE(w791) );
	vdp_slatch g842 (.nQ(w775), .D(w788), .C(w614), .nC(w615) );
	vdp_slatch g843 (.D(REG_BUS[0]), .C(w1546), .nC(w1547), .nQ(w6699) );
	vdp_slatch g844 (.D(w788), .C(w618), .nC(w619), .nQ(w6716) );
	vdp_slatch g845 (.D(REG_BUS[0]), .C(w1467), .nC(w621), .nQ(w6702) );
	vdp_slatch g846 (.D(w788), .C(w1466), .nC(w1548), .nQ(w6718) );
	vdp_slatch g847 (.D(REG_BUS[0]), .C(w625), .nC(w626), .nQ(w6732) );
	vdp_slatch g848 (.D(w788), .C(w1465), .nC(w628), .nQ(w6751) );
	vdp_slatch g849 (.D(REG_BUS[0]), .C(w1464), .nC(w1463), .nQ(w6736) );
	vdp_slatch g850 (.D(VRAMA[16]), .C(w1462), .nC(w630), .nQ(w6752) );
	vdp_slatch g851 (.Q(w6767), .D(VRAMA[0]), .C(w631), .nC(w632) );
	vdp_notif0 g852 (.nZ(VRAMA[0]), .nE(w847), .A(w6767) );
	vdp_notif0 g853 (.nZ(VRAMA[16]), .nE(w1461), .A(w6752) );
	vdp_notif0 g854 (.nZ(VRAMA[0]), .nE(w629), .A(w6736) );
	vdp_notif0 g855 (.nZ(VRAMA[16]), .nE(w1544), .A(w6751) );
	vdp_notif0 g856 (.nZ(VRAMA[0]), .nE(w624), .A(w6732) );
	vdp_notif0 g857 (.nZ(VRAMA[16]), .nE(w617), .A(w6716) );
	vdp_notif0 g858 (.nZ(VRAMA[0]), .nE(w1545), .A(w6702) );
	vdp_notif0 g859 (.nZ(VRAMA[16]), .nE(w622), .A(w6718) );
	vdp_notif0 g860 (.A(w775), .nZ(VRAMA[16]), .nE(w613) );
	vdp_notif0 g861 (.nZ(VRAMA[0]), .nE(w846), .A(w6699) );
	vdp_bufif0 g862 (.A(w788), .Z(VRAMA[16]), .nE(w1496) );
	vdp_bufif0 g863 (.A(REG_BUS[0]), .Z(VRAMA[0]), .nE(w1498) );
	vdp_bufif0 g864 (.A(w770), .Z(VRAMA[15]), .nE(w1497) );
	vdp_bufif0 g865 (.A(w770), .Z(CA[15]), .nE(w849) );
	vdp_bufif0 g866 (.A(w798), .Z(VRAMA[0]), .nE(w1495) );
	vdp_bufif0 g867 (.A(w798), .Z(CA[0]), .nE(w848) );
	vdp_slatch g868 (.Q(w789), .D(REG_BUS[0]), .C(w1589), .nC(w1590) );
	vdp_not g869 (.A(REG_BUS[7]), .nZ(w1593) );
	vdp_not g870 (.A(REG_BUS[0]), .nZ(w1469) );
	vdp_cnt_bit_load g871 (.D(REG_BUS[7]), .nL(w1592), .L(w1601), .R(1'b0), .Q(w770), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w783) );
	vdp_cnt_bit_load g872 (.D(REG_BUS[0]), .nL(w1432), .L(w803), .R(1'b0), .Q(w798), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w796), .CO(w784) );
	vdp_cnt_bit_load g873 (.D(w1593), .nL(w1591), .L(w812), .R(1'b0), .Q(w778), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w777) );
	vdp_cnt_bit_load g874 (.D(w1469), .nL(w793), .L(w794), .R(1'b0), .Q(w1468), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w796), .CO(w780) );
	vdp_nand3 g875 (.Z(w745), .B(w781), .A(w592), .C(w1427) );
	vdp_bufif0 g876 (.A(w789), .Z(CA[16]), .nE(w791) );
	vdp_slatch g877 (.D(VRAMA[8]), .C(w631), .nC(w632), .nQ(w6768) );
	vdp_slatch g878 (.D(w591), .C(w1464), .nC(w1463), .nQ(w6735) );
	vdp_slatch g879 (.D(w591), .C(w625), .nC(w626), .nQ(w6734) );
	vdp_slatch g880 (.D(w591), .C(w1467), .nC(w621), .nQ(w6701) );
	vdp_slatch g881 (.D(w591), .C(w1546), .nC(w1547), .nQ(w6700) );
	vdp_notif0 g882 (.nZ(VRAMA[8]), .nE(w846), .A(w6700) );
	vdp_notif0 g883 (.nZ(VRAMA[8]), .nE(w1545), .A(w6701) );
	vdp_notif0 g884 (.nZ(VRAMA[8]), .nE(w624), .A(w6734) );
	vdp_notif0 g885 (.nZ(VRAMA[8]), .nE(w629), .A(w6735) );
	vdp_notif0 g886 (.nZ(VRAMA[8]), .nE(w847), .A(w6768) );
	vdp_bufif0 g887 (.A(w789), .Z(VRAMA[16]), .nE(w1497) );
	vdp_not g888 (.A(w1460), .nZ(w1496) );
	vdp_not g889 (.A(w580), .nZ(w1498) );
	vdp_not g890 (.A(w33), .nZ(w1497) );
	vdp_not g891 (.A(w588), .nZ(w849) );
	vdp_not g892 (.A(w33), .nZ(w1495) );
	vdp_not g893 (.A(w588), .nZ(w848) );
	vdp_not g894 (.A(w588), .nZ(w791) );
	vdp_not g895 (.A(w1468), .nZ(w1427) );
	vdp_not g896 (.A(w792), .nZ(w1431) );
	vdp_not g897 (.A(M5), .nZ(w808) );
	vdp_and4 g898 (.Z(w804), .B(w678), .A(w814), .D(w591), .C(w815) );
	vdp_and4 g899 (.Z(w805), .B(w678), .A(w814), .D(w817), .C(w658) );
	vdp_and4 g900 (.B(w818), .A(w799), .D(w817), .C(w815), .Z(w807) );
	vdp_and4 g901 (.B(w818), .A(w799), .D(w591), .C(w815), .Z(w806) );
	vdp_and4 g902 (.Z(w801), .B(w815), .A(w591), .D(w819), .C(w678) );
	vdp_and4 g903 (.Z(w809), .B(w658), .A(w817), .D(w799), .C(w818) );
	vdp_and4 g904 (.Z(w800), .B(w658), .A(w591), .D(w819), .C(w678) );
	vdp_and4 g905 (.B(w822), .A(M5), .D(w702), .C(w823), .Z(w814) );
	vdp_comp_str g906 (.A(w825), .Z(w1589), .nZ(w1590) );
	vdp_comp_we g907 (.A(w1473), .Z(w1601), .nZ(w1592) );
	vdp_comp_we g908 (.A(w802), .Z(w803), .nZ(w1432) );
	vdp_comp_we g909 (.A(w826), .Z(w812), .nZ(w1591) );
	vdp_comp_we g910 (.A(w827), .Z(w794), .nZ(w793) );
	vdp_and g911 (.Z(w601), .B(w592), .A(w792) );
	vdp_and g912 (.Z(w796), .B(w592), .A(w1431) );
	vdp_or g913 (.Z(w825), .B(w800), .A(SYSRES) );
	vdp_or g914 (.Z(w802), .B(w801), .A(SYSRES) );
	vdp_or g915 (.Z(w1460), .B(w808), .A(w580) );
	vdp_or g916 (.B(w806), .A(SYSRES), .Z(w171) );
	vdp_or g917 (.B(w807), .A(SYSRES), .Z(w170) );
	vdp_or g918 (.Z(w169), .B(w805), .A(SYSRES) );
	vdp_or g919 (.Z(w68), .B(w804), .A(SYSRES) );
	vdp_or g920 (.B(w1470), .A(SYSRES), .Z(w72) );
	vdp_and4 g921 (.B(w678), .A(w816), .D(w591), .C(w658), .Z(w833) );
	vdp_or g922 (.B(w833), .A(SYSRES), .Z(w73) );
	vdp_and4 g923 (.B(w818), .A(w819), .D(w817), .C(w658), .Z(w832) );
	vdp_or g924 (.B(w832), .A(SYSRES), .Z(w74) );
	vdp_and4 g925 (.B(w818), .A(w819), .D(w591), .C(w815), .Z(w831) );
	vdp_or g926 (.B(w831), .A(SYSRES), .Z(w168) );
	vdp_and4 g927 (.B(w818), .A(w819), .D(w817), .C(w815), .Z(w1471) );
	vdp_or g928 (.B(w1471), .A(SYSRES), .Z(w69) );
	vdp_and4 g929 (.B(w678), .A(w816), .D(w817), .C(w658), .Z(w830) );
	vdp_or g930 (.B(w830), .A(SYSRES), .Z(w138) );
	vdp_and4 g931 (.B(w678), .A(w816), .D(w591), .C(w815), .Z(w829) );
	vdp_or g932 (.B(w829), .A(SYSRES), .Z(w137) );
	vdp_or g933 (.B(w834), .A(SYSRES), .Z(w71) );
	vdp_and4 g934 (.B(w678), .A(w816), .D(w817), .C(w815), .Z(w1470) );
	vdp_or g935 (.B(w835), .A(SYSRES), .Z(w70) );
	vdp_and4 g936 (.B(w818), .A(w816), .D(w591), .C(w658), .Z(w834) );
	vdp_and4 g937 (.B(w818), .A(w816), .D(w817), .C(w658), .Z(w835) );
	vdp_and4 g938 (.B(w815), .A(w591), .D(w816), .C(w818), .Z(w837) );
	vdp_or g939 (.B(w837), .A(SYSRES), .Z(w1131) );
	vdp_and4 g940 (.B(w815), .A(w817), .D(w816), .C(w818), .Z(w1472) );
	vdp_or g941 (.B(w1472), .A(SYSRES), .Z(w1171) );
	vdp_and4 g942 (.B(w815), .A(w817), .D(w814), .C(w678), .Z(w836) );
	vdp_or g943 (.B(w836), .A(SYSRES), .Z(w1132) );
	vdp_and4 g944 (.B(w658), .A(w817), .D(w819), .C(w678), .Z(w838) );
	vdp_or g945 (.B(w838), .A(SYSRES), .Z(w1473) );
	vdp_and4 g946 (.B(w658), .A(w591), .D(w814), .C(w818), .Z(w1474) );
	vdp_or g947 (.B(w1474), .A(SYSRES), .Z(CA[14]) );
	vdp_and4 g948 (.B(w815), .A(w817), .D(w819), .C(w678), .Z(w839) );
	vdp_or g949 (.B(w839), .A(SYSRES), .Z(w826) );
	vdp_and4 g950 (.B(w658), .A(w591), .D(w819), .C(w818), .Z(w840) );
	vdp_or g951 (.B(w840), .A(SYSRES), .Z(w827) );
	vdp_and4 g952 (.B(w658), .A(w591), .D(w814), .C(w678), .Z(w841) );
	vdp_or g953 (.B(w841), .A(SYSRES), .Z(w842) );
	vdp_and4 g954 (.B(w824), .A(w822), .D(M5), .C(w716), .Z(w819) );
	vdp_and3 g955 (.B(w823), .A(w822), .C(w702), .Z(w799) );
	vdp_and3 g956 (.B(w824), .A(w822), .C(w823), .Z(w816) );
	vdp_or g957 (.Z(w843), .B(w844), .A(w6670) );
	vdp_and g958 (.B(w821), .A(HCLK1), .Z(w822) );
	vdp_dlatch_inv g959 (.D(w820), .C(DCLK2), .nQ(w844), .nC(nDCLK2) );
	vdp_dlatch_inv g960 (.D(w6669), .C(HCLK2), .nQ(w821), .nC(nHCLK2) );
	vdp_not g961 (.A(w716), .nZ(w823) );
	vdp_not g962 (.A(w702), .nZ(w824) );
	vdp_not g963 (.A(w658), .nZ(w815) );
	vdp_not g964 (.A(w678), .nZ(w818) );
	vdp_not g965 (.A(w591), .nZ(w817) );
	vdp_slatch g966 (.D(REG_BUS[5]), .C(w625), .nC(w626), .nQ(w6728) );
	vdp_slatch g967 (.D(REG_BUS[4]), .C(w625), .nC(w626), .nQ(w6729) );
	vdp_sr_bit g968 (.D(w844), .C2(DCLK2), .C1(DCLK1), .Q(w6670), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_dlatch_inv g969 (.D(w843), .C(DCLK1), .nQ(w6669), .nC(nDCLK1) );
	vdp_comp_str g970 (.A(w881), .Z(w851), .nZ(w859) );
	vdp_fa g971 (.SUM(w878), .A(REG_BUS[6]), .B(w1566), .CO(w880), .CI(w876) );
	vdp_fa g972 (.SUM(w874), .A(REG_BUS[5]), .B(w875), .CO(w876), .CI(w873) );
	vdp_fa g973 (.SUM(w871), .A(REG_BUS[4]), .B(w872), .CO(w873), .CI(w868) );
	vdp_fa g974 (.SUM(w867), .A(REG_BUS[3]), .B(w870), .CO(w868), .CI(w865) );
	vdp_fa g975 (.SUM(w863), .A(REG_BUS[2]), .B(w864), .CO(w865), .CI(w862) );
	vdp_fa g976 (.SUM(w6673), .A(REG_BUS[1]), .B(w861), .CO(w862), .CI(w858) );
	vdp_fa g977 (.SUM(w6674), .A(REG_BUS[0]), .B(w855), .CO(w858), .CI(w853) );
	vdp_fa g978 (.SUM(w1475), .A(REG_BUS[7]), .B(w1565), .CO(w882), .CI(w880) );
	vdp_slatch g979 (.Q(w879), .D(DB[7]), .C(w851), .nC(w859) );
	vdp_aon22 g980 (.Z(w1576), .A1(w879), .A2(w850), .B1(w856), .B2(w1475) );
	vdp_slatch g981 (.Q(w877), .D(DB[6]), .C(w851), .nC(w859) );
	vdp_aon22 g982 (.Z(w1577), .A1(w877), .A2(w850), .B1(w856), .B2(w878) );
	vdp_slatch g983 (.Q(w1518), .D(DB[5]), .C(w851), .nC(w859) );
	vdp_aon22 g984 (.Z(w1578), .A1(w1518), .A2(w850), .B1(w856), .B2(w874) );
	vdp_slatch g985 (.Q(w869), .D(DB[4]), .C(w851), .nC(w859) );
	vdp_aon22 g986 (.Z(w1579), .A1(w869), .A2(w850), .B1(w856), .B2(w871) );
	vdp_slatch g987 (.Q(w866), .D(DB[3]), .C(w851), .nC(w859) );
	vdp_aon22 g988 (.Z(w1580), .A1(w866), .A2(w850), .B1(w856), .B2(w867) );
	vdp_slatch g989 (.Q(w860), .D(DB[2]), .C(w851), .nC(w859) );
	vdp_aon22 g990 (.Z(w1581), .A1(w860), .A2(w850), .B1(w856), .B2(w863) );
	vdp_slatch g991 (.Q(w857), .D(DB[1]), .C(w851), .nC(w859) );
	vdp_aon22 g992 (.Z(w1582), .A1(w857), .A2(w850), .B1(w856), .B2(w6673) );
	vdp_slatch g993 (.Q(w852), .D(DB[0]), .C(w851), .nC(w859) );
	vdp_aon22 g994 (.Z(w1583), .A1(w852), .A2(w850), .B1(w856), .B2(w6674) );
	vdp_dff g995 (.Q(REG_BUS[0]), .R(SYSRES), .C(w884), .D(w1583) );
	vdp_slatch g996 (.Q(w855), .D(REG_BUS[0]), .C(w883), .nC(w854) );
	vdp_dff g997 (.Q(REG_BUS[1]), .R(SYSRES), .D(w1582), .C(w884) );
	vdp_slatch g998 (.Q(w861), .D(REG_BUS[1]), .C(w883), .nC(w854) );
	vdp_dff g999 (.Q(REG_BUS[2]), .R(SYSRES), .C(w884), .D(w1581) );
	vdp_slatch g1000 (.Q(w864), .D(REG_BUS[2]), .C(w883), .nC(w854) );
	vdp_dff g1001 (.Q(REG_BUS[3]), .R(SYSRES), .D(w1580), .C(w884) );
	vdp_slatch g1002 (.Q(w870), .D(REG_BUS[3]), .C(w883), .nC(w854) );
	vdp_dff g1003 (.Q(REG_BUS[4]), .R(SYSRES), .C(w884), .D(w1579) );
	vdp_slatch g1004 (.Q(w872), .D(REG_BUS[4]), .C(w883), .nC(w854) );
	vdp_dff g1005 (.Q(REG_BUS[5]), .R(SYSRES), .C(w884), .D(w1578) );
	vdp_slatch g1006 (.Q(w875), .D(REG_BUS[5]), .C(w883), .nC(w854) );
	vdp_dff g1007 (.Q(REG_BUS[6]), .R(SYSRES), .C(w884), .D(w1577) );
	vdp_slatch g1008 (.Q(w1566), .D(REG_BUS[6]), .C(w883), .nC(w854) );
	vdp_dff g1009 (.Q(REG_BUS[7]), .R(SYSRES), .D(w1576), .C(w884) );
	vdp_slatch g1010 (.Q(w1565), .D(REG_BUS[7]), .C(w883), .nC(w854) );
	vdp_comp_str g1011 (.A(w842), .Z(w883), .nZ(w854) );
	vdp_comp_we g1012 (.A(w887), .Z(w850), .nZ(w856) );
	vdp_dff g1013 (.Q(w788), .R(w891), .C(w884), .D(w1567) );
	vdp_dff g1014 (.Q(w774), .R(w891), .C(w884), .D(w1568) );
	vdp_dff g1015 (.Q(w753), .R(w891), .C(w884), .D(w1569) );
	vdp_dff g1016 (.Q(w734), .R(SYSRES), .C(w884), .D(w1570) );
	vdp_dff g1017 (.Q(w716), .R(SYSRES), .C(w884), .D(w1571) );
	vdp_dff g1018 (.Q(w702), .R(SYSRES), .C(w884), .D(w1572) );
	vdp_dff g1019 (.Q(w678), .R(SYSRES), .C(w884), .D(w1573) );
	vdp_dff g1020 (.Q(w658), .R(SYSRES), .C(w884), .D(w1574) );
	vdp_dff g1021 (.Q(w591), .R(SYSRES), .C(w884), .D(w1575) );
	vdp_not g1022 (.A(w913), .nZ(w884) );
	vdp_or g1023 (.Z(w891), .B(SYSRES), .A(w853) );
	vdp_not g1024 (.A(M5), .nZ(w853) );
	vdp_slatch g1025 (.Q(w910), .D(w278), .C(w924), .nC(w901) );
	vdp_aon22 g1026 (.Z(w1575), .A1(w914), .A2(w922), .B1(w888), .B2(w912) );
	vdp_slatch g1027 (.Q(w914), .D(w243), .C(w924), .nC(w901) );
	vdp_comp_str g1028 (.A(w928), .Z(w924), .nZ(w901) );
	vdp_comp_we g1029 (.A(w887), .Z(w922), .nZ(w888) );
	vdp_ha g1030 (.SUM(w912), .A(w591), .B(w882), .CO(w909) );
	vdp_slatch g1031 (.Q(w908), .D(w251), .C(w924), .nC(w901) );
	vdp_aon22 g1032 (.Z(w1574), .A1(w910), .A2(w922), .B1(w888), .B2(w911) );
	vdp_ha g1033 (.SUM(w911), .A(w658), .B(w909), .CO(w1586) );
	vdp_slatch g1034 (.Q(w906), .D(w287), .C(w924), .nC(w901) );
	vdp_aon22 g1035 (.Z(w1573), .A1(w908), .A2(w922), .B1(w888), .B2(w907) );
	vdp_ha g1036 (.SUM(w907), .A(w678), .B(w1586), .CO(w905) );
	vdp_slatch g1037 (.Q(w903), .D(w260), .C(w924), .nC(w901) );
	vdp_aon22 g1038 (.Z(w1572), .A1(w906), .A2(w922), .B1(w888), .B2(w904) );
	vdp_ha g1039 (.SUM(w904), .A(w702), .B(w905), .CO(w1585) );
	vdp_slatch g1040 (.Q(w900), .D(w296), .C(w924), .nC(w901) );
	vdp_aon22 g1041 (.Z(w1571), .A1(w903), .A2(w922), .B1(w888), .B2(w902) );
	vdp_ha g1042 (.SUM(w902), .A(w716), .B(w1585), .CO(w899) );
	vdp_aon22 g1043 (.Z(w1570), .A1(w900), .A2(w922), .B1(w888), .B2(w897) );
	vdp_ha g1044 (.SUM(w897), .A(w734), .B(w899), .CO(w898) );
	vdp_comp_str g1045 (.A(w923), .Z(w921), .nZ(w890) );
	vdp_aon22 g1046 (.Z(w1569), .A1(w896), .A2(w922), .B1(w888), .B2(w1584) );
	vdp_ha g1047 (.SUM(w1584), .A(w753), .B(w898), .CO(w893) );
	vdp_slatch_r g1048 (.Q(w896), .D(DB[0]), .R(w891), .C(w921), .nC(w890) );
	vdp_slatch_r g1049 (.Q(w895), .D(DB[1]), .R(w891), .C(w921), .nC(w890) );
	vdp_aon22 g1050 (.Z(w1568), .A1(w895), .A2(w922), .B1(w888), .B2(w894) );
	vdp_ha g1051 (.SUM(w894), .A(w774), .B(w893), .CO(w892) );
	vdp_slatch_r g1052 (.Q(w889), .D(DB[2]), .R(w891), .C(w921), .nC(w890) );
	vdp_aon22 g1053 (.Z(w1567), .A1(w889), .A2(w922), .B1(w888), .B2(w1517) );
	vdp_ha g1054 (.SUM(w1517), .A(w788), .B(w892) );
	vdp_and3 g1055 (.C(w918), .A(w916), .B(w917), .Z(w920) );
	vdp_sr_bit g1056 (.D(w1481), .C2(HCLK2), .C1(HCLK1), .nQ(w105), .nC1(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1057 (.D(w937), .Q(w1481), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK2), .nC1(nHCLK1) );
	vdp_not g1058 (.A(w963), .nZ(w939) );
	vdp_not g1059 (.A(w466), .nZ(w1482) );
	vdp_not g1060 (.A(w467), .nZ(w950) );
	vdp_not g1061 (.A(w916), .nZ(w951) );
	vdp_not g1062 (.A(w948), .nZ(w956) );
	vdp_not g1063 (.A(w509), .nZ(w933) );
	vdp_not g1064 (.A(w585), .nZ(w945) );
	vdp_not g1065 (.A(w970), .nZ(w959) );
	vdp_not g1066 (.A(w1483), .nZ(w962) );
	vdp_not g1067 (.A(w960), .nZ(w929) );
	vdp_slatch g1068 (.Q(w493), .D(w926), .C(w927), .nC(w940) );
	vdp_slatch g1069 (.Q(w509), .D(w269), .C(w927), .nC(w940) );
	vdp_comp_str g1070 (.A(w928), .Z(w927), .nZ(w940) );
	vdp_dlatch_inv g1071 (.D(w593), .C(DCLK1), .nQ(w960), .nC(nDCLK1) );
	vdp_dlatch_inv g1072 (.D(w959), .C(DCLK1), .nQ(w958), .nC(nDCLK1) );
	vdp_dlatch_inv g1073 (.D(w972), .C(DCLK2), .nQ(w970), .nC(nDCLK2) );
	vdp_dlatch_inv g1074 (.D(w977), .C(DCLK1), .nQ(w972), .nC(nDCLK1) );
	vdp_slatch g1075 (.Q(w977), .D(w935), .C(DCLK2), .nC(nDCLK2) );
	vdp_slatch g1076 (.Q(w935), .D(w971), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g1077 (.D(w580), .C(HCLK1), .nQ(w934), .nC(nHCLK1) );
	vdp_rs_ff g1078 (.nQ(w931), .R(w979), .S(w978), .Q(w943) );
	vdp_rs_ff g1079 (.Q(w955), .R(w953), .S(w932) );
	vdp_and3 g1080 (.C(w420), .A(w467), .B(w1482), .Z(w938) );
	vdp_and3 g1081 (.C(w950), .A(w466), .B(w420), .Z(w104) );
	vdp_comp_dff g1082 (.D(w954), .C2(HCLK2), .C1(HCLK1), .Q(w947), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_comp_dff g1083 (.D(w944), .C2(HCLK2), .C1(HCLK1), .Q(w946), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g1084 (.C(w32), .A(w943), .B(w587), .Z(w944) );
	vdp_and g1085 (.A(DB[7]), .B(w923), .Z(w925) );
	vdp_and g1086 (.A(w934), .B(w977), .Z(w887) );
	vdp_and g1087 (.A(w946), .B(w945), .Z(w568) );
	vdp_and g1088 (.A(w585), .B(w946), .Z(w589) );
	vdp_and g1089 (.A(w947), .B(w945), .Z(w957) );
	vdp_and g1090 (.A(w585), .B(w947), .Z(w33) );
	vdp_or g1091 (.A(w947), .B(w968), .Z(w953) );
	vdp_or g1092 (.A(w947), .B(w568), .Z(w420) );
	vdp_or g1093 (.A(w585), .B(w448), .Z(w976) );
	vdp_aoi21 g1094 (.A1(w958), .B(SYSRES), .Z(w1483), .A2(w959) );
	vdp_or3 g1095 (.C(w930), .A(w952), .B(w920), .Z(w932) );
	vdp_or3 g1096 (.C(w589), .A(w957), .B(w583), .Z(w580) );
	vdp_or5 g1097 (.C(w941), .A(w929), .B(w580), .Z(w913), .D(w928), .E(w923) );
	vdp_nand3 g1098 (.C(w919), .A(w956), .B(w966), .Z(w820) );
	vdp_2a3oi g1099 (.A1(w918), .B(w973), .Z(w967), .A2(w966), .C(w917) );
	vdp_nand g1100 (.A(w493), .B(w933), .Z(w948) );
	vdp_nor g1101 (.A(w935), .B(w972), .Z(w919) );
	vdp_and4 g1102 (.C(w931), .A(w587), .B(w32), .Z(w954), .D(w955) );
	vdp_nor5 g1103 (.C(w509), .A(w981), .B(w967), .Z(w930), .D(w493), .E(w951) );
	vdp_and g1104 (.A(w585), .B(w981), .Z(w952) );
	vdp_not g1105 (.A(w573), .nZ(w1535) );
	vdp_not g1106 (.A(w1535), .nZ(w1015) );
	vdp_not g1107 (.A(w996), .nZ(w1032) );
	vdp_not g1108 (.A(w972), .nZ(w1488) );
	vdp_not g1109 (.A(w977), .nZ(w1017) );
	vdp_not g1110 (.A(w1020), .nZ(w928) );
	vdp_not g1111 (.A(w403), .nZ(w949) );
	vdp_not g1112 (.A(w1005), .nZ(w1013) );
	vdp_not g1113 (.A(M5), .nZ(w918) );
	vdp_rs_ff g1114 (.Q(w966), .R(w964), .S(w928) );
	vdp_rs_ff g1115 (.Q(w917), .R(w964), .S(w1040) );
	vdp_rs_ff g1116 (.Q(w973), .R(w964), .S(w923) );
	vdp_rs_ff g1117 (.nQ(w975), .R(w974), .S(w942) );
	vdp_rs_ff g1118 (.Q(w1037), .R(w962), .S(w969) );
	vdp_rs_ff g1119 (.Q(w563), .R(w962), .S(w1030) );
	vdp_rs_ff g1120 (.Q(w562), .R(w962), .S(w987) );
	vdp_or g1121 (.A(w987), .B(w1030), .Z(w1039) );
	vdp_and g1122 (.A(w1037), .B(w916), .Z(w570) );
	vdp_and g1123 (.A(w1036), .B(w1037), .Z(w573) );
	vdp_and g1124 (.A(w1017), .B(w1488), .Z(w916) );
	vdp_and g1125 (.A(w1017), .B(w970), .Z(w1036) );
	vdp_and g1126 (.A(w972), .B(w970), .Z(w1003) );
	vdp_and g1127 (.A(w947), .B(w976), .Z(w978) );
	vdp_and g1128 (.A(w999), .B(w988), .Z(w411) );
	vdp_and g1129 (.A(w949), .B(w881), .Z(w1046) );
	vdp_and g1130 (.A(w1023), .B(w1022), .Z(w969) );
	vdp_or g1131 (.A(w946), .B(w968), .Z(w979) );
	vdp_or g1132 (.A(w1016), .B(w1019), .Z(w961) );
	vdp_or g1133 (.A(SYSRES), .B(w916), .Z(w974) );
	vdp_or g1134 (.A(SYSRES), .B(w977), .Z(w1043) );
	vdp_or g1135 (.A(w972), .B(w971), .Z(w1038) );
	vdp_or g1136 (.A(w999), .B(w1023), .Z(w1044) );
	vdp_or g1137 (.A(w965), .B(SYSRES), .Z(w1009) );
	vdp_or g1138 (.A(SYSRES), .B(w1004), .Z(w1048) );
	vdp_or g1139 (.A(SYSRES), .B(w1003), .Z(w964) );
	vdp_and g1140 (.A(w963), .B(w938), .Z(w126) );
	vdp_and g1141 (.A(w938), .B(w939), .Z(w103) );
	vdp_and g1142 (.A(w916), .B(w1011), .Z(w1047) );
	vdp_nand g1143 (.A(w411), .B(w975), .Z(w1028) );
	vdp_nor g1144 (.A(w1033), .B(w1015), .Z(w1029) );
	vdp_or5 g1145 (.C(w928), .A(w1014), .B(w1027), .Z(w1026), .D(w881), .E(w1031) );
	vdp_or3 g1146 (.C(w1018), .A(w999), .B(w406), .Z(w1019) );
	vdp_nor g1147 (.A(w104), .B(w938), .Z(w937) );
	vdp_and3 g1148 (.C(w1049), .A(w1045), .B(w1001), .Z(w1021) );
	vdp_or4 g1149 (.C(w969), .A(w923), .B(w998), .Z(w965), .D(w411) );
	vdp_and4 g1150 (.C(w1045), .A(w1023), .B(w1006), .Z(w881), .D(w1024) );
	vdp_aoi21 g1151 (.A1(w916), .B(SYSRES), .Z(w1005), .A2(w1012) );
	vdp_aoi21 g1152 (.A1(w881), .B(w1021), .Z(w1020), .A2(w403) );
	vdp_or5 g1153 (.C(w411), .A(w998), .B(w923), .Z(w1004), .D(w969), .E(w928) );
	vdp_and5 g1154 (.C(w1010), .A(M5), .B(w1045), .Z(w923), .D(w1024), .E(w1023) );
	vdp_not g1155 (.A(CA[7]), .nZ(w992) );
	vdp_not g1156 (.A(w1023), .nZ(w1000) );
	vdp_not g1157 (.A(w1000), .nZ(w985) );
	vdp_not g1158 (.A(w999), .nZ(w984) );
	vdp_not g1159 (.A(w984), .nZ(w983) );
	vdp_slatch g1160 (.Q(w1025), .D(w986), .nC(w983), .C(w984) );
	vdp_slatch g1161 (.Q(w1045), .D(w986), .nC(w985), .C(w1000), .nQ(w1022) );
	vdp_rs_ff g1162 (.Q(w1007), .R(w1003), .S(w1009) );
	vdp_rs_ff g1163 (.Q(w1011), .R(w1048), .S(w1046), .nQ(w1012) );
	vdp_rs_ff g1164 (.Q(w1049), .R(w1013), .S(w1047), .nQ(w1024) );
	vdp_rs_ff g1165 (.Q(w1010), .R(w1008), .S(w1479), .nQ(w1006) );
	vdp_slatch_r g1166 (.Q(w981), .D(DB[6]), .C(w1002), .nC(w982), .R(w891) );
	vdp_slatch_r g1167 (.Q(w467), .D(DB[5]), .R(w891), .C(w1002), .nC(w982) );
	vdp_slatch_r g1168 (.Q(w466), .D(DB[4]), .R(w891), .C(w1002), .nC(w982) );
	vdp_comp_str g1169 (.A(w923), .Z(w1002), .nZ(w982) );
	vdp_not g1170 (.A(w1480), .nZ(w1008) );
	vdp_aoi21 g1171 (.A1(w916), .B(SYSRES), .Z(w1480), .A2(w1007) );
	vdp_and4 g1172 (.C(w948), .A(M5), .B(w966), .Z(w1479), .D(w916) );
	vdp_and g1173 (.A(w999), .B(w1025), .Z(w1040) );
	vdp_rs_ff g1174 (.nQ(w1042), .R(w1041), .S(w1040) );
	vdp_rs_ff g1175 (.Q(w971), .R(w1043), .S(w1044) );
	vdp_not g1176 (.A(w986), .nZ(w1587) );
	vdp_not g1177 (.A(CA[2]), .nZ(w1073) );
	vdp_not g1178 (.A(CA[3]), .nZ(w1074) );
	vdp_aon22 g1179 (.Z(w986), .A1(CA[0]), .A2(w1100), .B1(w403), .B2(CA[1]) );
	vdp_and4 g1180 (.C(w991), .A(w992), .B(CA[6]), .Z(w1035), .D(w990) );
	vdp_and4 g1181 (.C(w995), .A(w994), .B(CA[7]), .Z(w1001), .D(w990) );
	vdp_and4 g1182 (.C(CA[3]), .A(w1032), .B(w1034), .Z(w1018), .D(CA[9]) );
	vdp_and4 g1183 (.C(CA[2]), .A(w1032), .B(w1034), .Z(w402), .D(w1074) );
	vdp_and4 g1184 (.C(w996), .A(w1073), .B(CA[3]), .Z(w993), .D(w1034) );
	vdp_or g1185 (.A(w1035), .B(w402), .Z(w406) );
	vdp_and g1186 (.A(w969), .B(w1029), .Z(w1027) );
	vdp_and g1187 (.A(w1019), .B(w1028), .Z(w1031) );
	vdp_and g1188 (.A(w403), .B(w1026), .Z(w1064) );
	vdp_or g1189 (.A(SYSRES), .B(w942), .Z(w1041) );
	vdp_or g1190 (.A(w1001), .B(w989), .Z(w1023) );
	vdp_or g1191 (.A(SYSRES), .B(w590), .Z(w968) );
	vdp_and3 g1192 (.C(w1072), .A(w923), .B(w1042), .Z(w1014) );
	vdp_and3 g1193 (.C(w1075), .A(w1038), .B(w1205), .Z(w1034) );
	vdp_and5 g1194 (.C(CA[2]), .A(w996), .B(CA[3]), .Z(w1069), .D(w1587), .E(w1034) );
	vdp_and5 g1195 (.C(CA[2]), .A(w996), .B(w986), .Z(w1068), .D(CA[3]), .E(w1034) );
	vdp_and5 g1196 (.C(w1073), .A(w1039), .B(w1032), .Z(w997), .D(w1074), .E(w1034) );
	vdp_and5 g1197 (.C(w1074), .A(w1073), .B(w1039), .Z(w989), .D(w996), .E(w1034) );
	vdp_nor5 g1198 (.C(w1065), .A(w1068), .B(w1069), .Z(w1051), .D(w993), .E(w1064) );
	vdp_aon22 g1199 (.Z(w1062), .A1(w4), .A2(w1071), .B1(w27), .B2(w403) );
	vdp_aon22 g1200 (.Z(w174), .A1(LS0), .A2(VPOS[8]), .B1(w1059), .B2(VPOS[0]) );
	vdp_not g1201 (.A(LS0), .nZ(w1059) );
	vdp_not g1202 (.A(w403), .nZ(w1055) );
	vdp_not g1203 (.A(w403), .nZ(w1071) );
	vdp_not g1204 (.A(w1532), .nZ(w109) );
	vdp_not g1205 (.A(CA[6]), .nZ(w994) );
	vdp_not g1206 (.A(w1477), .nZ(w1060) );
	vdp_not g1207 (.A(w986), .nZ(w988) );
	vdp_aoi21 g1208 (.A1(w987), .B(w1478), .Z(w1477), .A2(w993) );
	vdp_and4 g1209 (.C(w991), .A(w994), .B(CA[7]), .Z(w1476), .D(w990) );
	vdp_and4 g1210 (.C(w995), .A(w992), .B(CA[6]), .Z(w1478), .D(w990) );
	vdp_slatch g1211 (.Q(w111), .D(w991), .C(w1588), .nC(w1533) );
	vdp_comp_we g1212 (.A(PSG_Z80_CLK), .Z(w1588), .nZ(w1533) );
	vdp_and g1213 (.A(w47), .B(w1066), .Z(w1534) );
	vdp_and g1214 (.A(w986), .B(w999), .Z(w998) );
	vdp_or g1215 (.A(w997), .B(w1476), .Z(w999) );
	vdp_or g1216 (.A(w1065), .B(w1534), .Z(w1067) );
	vdp_or g1217 (.Z(w1061), .A(w7), .B(SYSRES) );
	vdp_and g1218 (.Z(w107), .A(w58), .B(w1062) );
	vdp_rs_ff g1219 (.Q(w1057), .R(w1061), .S(w107) );
	vdp_aoi221 g1220 (.Z(w1532), .A1(w108), .A2(1'b0), .B1(w1063), .B2(w1067), .C(w110) );
	vdp_aoi22 g1221 (.Z(w1052), .A1(w1058), .A2(w1055), .B1(w403), .B2(w1057) );
	vdp_comp_str g1222 (.Z(w1088), .A(w58), .nZ(w1089) );
	vdp_comp_str g1223 (.Z(w1114), .A(CA[14]), .nZ(w1115) );
	vdp_comp_str g1224 (.Z(w1124), .A(w1132), .nZ(w1125) );
	vdp_comp_str g1225 (.Z(w1121), .A(w1131), .nZ(w1120) );
	vdp_not g1226 (.A(w1130), .nZ(w1133) );
	vdp_not g1227 (.A(w1122), .nZ(w1135) );
	vdp_not g1228 (.A(w1119), .nZ(w1134) );
	vdp_not g1229 (.A(w1134), .nZ(w1099) );
	vdp_not g1230 (.A(w403), .nZ(w1100) );
	vdp_not g1231 (.A(w1135), .nZ(w1118) );
	vdp_not g1232 (.A(w1137), .nZ(w1117) );
	vdp_not g1233 (.A(w1136), .nZ(w1116) );
	vdp_aon222 g1234 (.C2(w1116), .B2(w1117), .A2(w1118), .C1(w1097), .B1(CA[15]), .A1(CA[7]), .Z(w1109) );
	vdp_aon222 g1235 (.C2(w1116), .B2(w1117), .A2(w1118), .C1(w1096), .B1(CA[13]), .A1(CA[6]), .Z(w1108) );
	vdp_aon222 g1236 (.C2(w1116), .B2(w1117), .A2(w1118), .C1(w1095), .B1(CA[12]), .A1(CA[5]), .Z(w1107) );
	vdp_aon222 g1237 (.C2(w1116), .B2(w1117), .A2(w1118), .C1(w1094), .B1(CA[11]), .A1(CA[4]), .Z(w1106) );
	vdp_aon222 g1238 (.C2(w1116), .B2(w1117), .A2(w1118), .C1(w1098), .B1(CA[10]), .A1(CA[3]), .Z(w1105) );
	vdp_aon222 g1239 (.C2(w1116), .B2(w1117), .A2(w1118), .C1(w1516), .B1(CA[9]), .A1(CA[2]), .Z(w1104) );
	vdp_aon222 g1240 (.C2(w1116), .B2(w1117), .A2(w1118), .C1(w1101), .B1(CA[8]), .A1(CA[1]), .Z(w1103) );
	vdp_aon222 g1241 (.C2(w1116), .B2(w1117), .A2(w1118), .C1(w1091), .B1(CA[14]), .A1(CA[0]), .Z(w1102) );
	vdp_aon222 g1242 (.C2(w1116), .B2(w1117), .A2(w1118), .C1(nHCLK1), .B1(1'b1), .A1(1'b0), .Z(w1119) );
	vdp_slatch g1243 (.Q(LS0), .D(w1111), .C(w1088), .nC(w1089) );
	vdp_slatch g1244 (.Q(w1087), .D(w1123), .C(w1088), .nC(w1089) );
	vdp_aon22 g1245 (.Z(w1090), .A1(COL[6]), .A2(w1126), .B1(w124), .B2(w1486) );
	vdp_not g1246 (.A(w1113), .nZ(w1085) );
	vdp_not g1247 (.A(w1126), .nZ(w1486) );
	vdp_and g1248 (.Z(w1), .A(w1087), .B(LS0) );
	vdp_and g1249 (.Z(w1086), .A(M5), .B(w1085) );
	vdp_and g1250 (.Z(w1487), .A(M5), .B(w1113) );
	vdp_and g1251 (.Z(128k), .A(M5), .B(w1112) );
	vdp_or3 g1252 (.Z(w1130), .A(w1127), .B(w1128), .C(w1393) );
	vdp_and g1253 (.Z(w1129), .A(w1127), .B(w1099) );
	vdp_nand g1254 (.Z(w1137), .A(w1135), .B(w1130) );
	vdp_nand g1255 (.Z(w1136), .A(w1135), .B(w1133) );
	vdp_slatch g1256 (.Q(w86), .D(REG_BUS[0]), .C(w1114), .nC(w1115) );
	vdp_slatch g1257 (.Q(w88), .D(REG_BUS[1]), .C(w1114), .nC(w1115) );
	vdp_slatch g1258 (.Q(w44), .D(REG_BUS[2]), .C(w1114), .nC(w1115) );
	vdp_slatch g1259 (.Q(w1138), .D(REG_BUS[3]), .C(w1114), .nC(w1115) );
	vdp_slatch g1260 (.Q(w106), .D(REG_BUS[4]), .C(w1114), .nC(w1115) );
	vdp_slatch g1261 (.Q(w89), .D(REG_BUS[5]), .C(w1114), .nC(w1115) );
	vdp_slatch g1262 (.Q(w1066), .D(REG_BUS[6]), .C(w1114), .nC(w1115) );
	vdp_slatch g1263 (.Q(w1122), .D(REG_BUS[7]), .C(w1114), .nC(w1115) );
	vdp_slatch g1264 (.Q(w1113), .D(REG_BUS[3]), .C(w1121), .nC(w1120) );
	vdp_slatch g1265 (.Q(w1112), .D(REG_BUS[7]), .C(w1121), .nC(w1120) );
	vdp_slatch g1266 (.Q(w19), .D(REG_BUS[4]), .C(w1124), .nC(w1125) );
	vdp_slatch g1267 (.Q(w84), .D(REG_BUS[3]), .C(w1124), .nC(w1125) );
	vdp_slatch g1268 (.Q(w1123), .D(REG_BUS[2]), .C(w1124), .nC(w1125) );
	vdp_slatch g1269 (.Q(w1111), .D(REG_BUS[1]), .C(w1124), .nC(w1125) );
	vdp_slatch g1270 (.Q(H40), .D(REG_BUS[0]), .C(w1124), .nC(w1125) );
	vdp_slatch g1271 (.Q(w45), .D(REG_BUS[0]), .C(w1121), .nC(w1120) );
	vdp_slatch g1272 (.Q(w127), .D(REG_BUS[1]), .C(w1121), .nC(w1120) );
	vdp_slatch g1273 (.Q(M5), .D(REG_BUS[2]), .C(w1121), .nC(w1120) );
	vdp_slatch g1274 (.Q(w1140), .D(REG_BUS[4]), .C(w1121), .nC(w1120) );
	vdp_slatch g1275 (.Q(w1139), .D(REG_BUS[5]), .C(w1121), .nC(w1120) );
	vdp_slatch g1276 (.Q(w1110), .D(REG_BUS[6]), .C(w1121), .nC(w1120) );
	vdp_and g1277 (.Z(w114), .A(w1068), .B(w1149) );
	vdp_and g1278 (.Z(w118), .A(w1018), .B(w1149) );
	vdp_and g1279 (.Z(w113), .A(w1068), .B(w1150) );
	vdp_and g1280 (.Z(w117), .A(w1018), .B(w1150) );
	vdp_and g1281 (.Z(w115), .A(w1068), .B(w1144) );
	vdp_and g1282 (.Z(w116), .A(w1018), .B(w1144) );
	vdp_and g1283 (.Z(w57), .A(w1068), .B(w1145) );
	vdp_and g1284 (.Z(w48), .A(w1018), .B(w1145) );
	vdp_and g1285 (.Z(w85), .A(w1068), .B(w1147) );
	vdp_and g1286 (.Z(w83), .A(w1018), .B(w1147) );
	vdp_and g1287 (.Z(w87), .A(w1068), .B(w1148) );
	vdp_and g1288 (.Z(PSG_TEST_OE), .A(w1018), .B(w1148) );
	vdp_and g1289 (.Z(w1167), .A(w1068), .B(w1152) );
	vdp_and g1290 (.Z(w1141), .A(w1068), .B(w1153) );
	vdp_and g1291 (.Z(w56), .A(w1068), .B(w1146) );
	vdp_and g1292 (.Z(w54), .A(w1018), .B(w1146) );
	vdp_dlatch g1293 (.D(COL[0]), .C(HCLK1), .Q(w1091), .nC(nHCLK1) );
	vdp_dlatch g1294 (.D(COL[1]), .Q(w1101), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch g1295 (.D(COL[2]), .Q(w1516), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch g1296 (.D(COL[3]), .Q(w1098), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch g1297 (.D(COL[4]), .Q(w1094), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch g1298 (.D(COL[5]), .Q(w1095), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch g1299 (.D(w1090), .Q(w1096), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch g1300 (.D(w125), .Q(w1097), .C(HCLK1), .nC(nHCLK1) );
	vdp_slatch g1301 (.Q(w52), .D(REG_BUS[5]), .C(w1125), .nC(w1124) );
	vdp_slatch g1302 (.Q(w39), .D(REG_BUS[6]), .C(w1125), .nC(w1124) );
	vdp_slatch g1303 (.Q(w1142), .D(REG_BUS[7]), .C(w1125), .nC(w1124) );
	vdp_slatch g1304 (.Q(w23), .D(REG_BUS[3]), .nC(w1175), .C(w1173) );
	vdp_slatch g1305 (.Q(w92), .D(REG_BUS[2]), .nC(w1175), .C(w1173) );
	vdp_slatch g1306 (.Q(w472), .D(REG_BUS[1]), .nC(w1175), .C(w1173) );
	vdp_slatch g1307 (.Q(w53), .D(REG_BUS[0]), .nC(w1175), .C(w1173) );
	vdp_slatch g1308 (.Q(w90), .D(REG_BUS[7]), .nC(w1175), .C(w1173) );
	vdp_slatch g1309 (.Q(w91), .D(REG_BUS[6]), .nC(w1175), .C(w1173) );
	vdp_slatch g1310 (.Q(w59), .D(REG_BUS[5]), .nC(w1175), .C(w1173) );
	vdp_slatch g1311 (.Q(w1172), .D(REG_BUS[4]), .nC(w1175), .C(w1173) );
	vdp_slatch_r g1312 (.Q(w119), .D(DB[14]), .nC(w1166), .R(w1161), .C(w1170) );
	vdp_slatch_r g1313 (.Q(w123), .D(DB[13]), .R(w1161), .nC(w1166), .C(w1170) );
	vdp_slatch_r g1314 (.Q(w120), .D(DB[12]), .R(w1161), .nC(w1166), .C(w1170) );
	vdp_comp_str g1315 (.Z(w1173), .A(w1171), .nZ(w1175) );
	vdp_comp_str g1316 (.Z(w1169), .A(w1141), .nZ(w1168) );
	vdp_not g1317 (.A(REG_BUS[6]), .nZ(w1484) );
	vdp_not g1318 (.A(REG_BUS[7]), .nZ(w1189) );
	vdp_not g1319 (.A(REG_BUS[4]), .nZ(w1176) );
	vdp_not g1320 (.A(REG_BUS[5]), .nZ(w1174) );
	vdp_not g1321 (.A(REG_BUS[2]), .nZ(w1190) );
	vdp_not g1322 (.A(REG_BUS[3]), .nZ(w1177) );
	vdp_not g1323 (.A(REG_BUS[0]), .nZ(w1184) );
	vdp_not g1324 (.A(REG_BUS[1]), .nZ(w1185) );
	vdp_not g1325 (.A(w1159), .nZ(w1179) );
	vdp_not g1326 (.A(w1160), .nZ(w1164) );
	vdp_not g1327 (.A(w1151), .nZ(w1178) );
	vdp_not g1328 (.A(w1165), .nZ(w1180) );
	vdp_comp_str g1329 (.Z(w1163), .nZ(w1162), .A(w1069) );
	vdp_slatch_r g1330 (.Q(w1165), .R(w1161), .D(DB[11]), .nC(w1162), .C(w1163) );
	vdp_slatch_r g1331 (.Q(w1151), .D(DB[10]), .nC(w1162), .R(w1161), .C(w1163) );
	vdp_and4 g1332 (.Z(w1493), .A(w1159), .B(w1160), .C(w1165), .D(w1151) );
	vdp_and4 g1333 (.Z(w1144), .A(w1165), .B(w1178), .C(w1164), .D(w1179) );
	vdp_and4 g1334 (.Z(w1150), .A(w1180), .B(w1151), .C(w1160), .D(w1159) );
	vdp_and4 g1335 (.Z(w1149), .A(w1180), .B(w1151), .C(w1160), .D(w1179) );
	vdp_and4 g1336 (.Z(w1148), .A(w1180), .B(w1151), .C(w1164), .D(w1159) );
	vdp_and4 g1337 (.Z(w1147), .A(w1180), .B(w1151), .C(w1164), .D(w1179) );
	vdp_and4 g1338 (.Z(w1145), .A(w1180), .B(w1178), .C(w1160), .D(w1159) );
	vdp_and4 g1339 (.Z(w1146), .A(w1180), .B(w1178), .C(w1160), .D(w1179) );
	vdp_and4 g1340 (.Z(w1153), .A(w1180), .B(w1178), .C(w1164), .D(w1159) );
	vdp_and4 g1341 (.Z(w1152), .A(w1180), .B(w1178), .C(w1164), .D(w1179) );
	vdp_nand g1342 (.Z(w1430), .A(w1493), .B(w1068) );
	vdp_slatch_r g1343 (.Q(w1159), .D(DB[8]), .R(w1161), .C(w1163), .nC(w1162) );
	vdp_slatch_r g1344 (.Q(w1158), .D(DB[11]), .R(w1161), .C(w1170), .nC(w1166) );
	vdp_slatch_r g1345 (.nC(w1162), .Q(w1160), .D(DB[9]), .R(w1161), .C(w1163) );
	vdp_slatch_r g1346 (.Q(w1157), .D(DB[10]), .R(w1161), .C(w1170), .nC(w1166) );
	vdp_slatch_r g1347 (.Q(w94), .D(DB[8]), .R(w1161), .C(w1170), .nC(w1166) );
	vdp_slatch_r g1348 (.Q(w1156), .D(DB[9]), .R(w1161), .C(w1170), .nC(w1166) );
	vdp_slatch_r g1349 (.Q(w93), .D(DB[7]), .R(w1161), .C(w1170), .nC(w1166) );
	vdp_slatch_r g1350 (.Q(w95), .D(DB[5]), .R(w1161), .C(w1170), .nC(w1166) );
	vdp_slatch_r g1351 (.Q(w96), .D(DB[6]), .R(w1161), .C(w1170), .nC(w1166) );
	vdp_slatch_r g1352 (.Q(w963), .D(DB[4]), .R(w1161), .C(w1170), .nC(w1166) );
	vdp_slatch_r g1353 (.Q(w1187), .D(DB[2]), .R(w1161), .C(w1170), .nC(w1166) );
	vdp_slatch_r g1354 (.Q(w1188), .D(DB[3]), .R(w1161), .C(w1170), .nC(w1166) );
	vdp_slatch_r g1355 (.Q(w1126), .D(DB[0]), .R(w1161), .C(w1170), .nC(w1166) );
	vdp_slatch_r g1356 (.Q(w792), .D(DB[1]), .R(w1161), .C(w1170), .nC(w1166) );
	vdp_slatch_r g1357 (.Q(w100), .D(DB[9]), .R(w1161), .C(w1169), .nC(w1168) );
	vdp_slatch_r g1358 (.Q(w101), .D(DB[10]), .R(w1161), .C(w1169), .nC(w1168) );
	vdp_slatch_r g1359 (.Q(w98), .D(DB[7]), .R(w1161), .C(w1169), .nC(w1168) );
	vdp_slatch_r g1360 (.Q(w99), .D(DB[8]), .R(w1161), .C(w1169), .nC(w1168) );
	vdp_slatch_r g1361 (.Q(w51), .D(DB[5]), .R(w1161), .C(w1169), .nC(w1168) );
	vdp_slatch_r g1362 (.Q(w41), .D(DB[6]), .R(w1161), .C(w1169), .nC(w1168) );
	vdp_slatch_r g1363 (.Q(w40), .D(DB[3]), .R(w1161), .C(w1169), .nC(w1168) );
	vdp_slatch_r g1364 (.Q(w42), .D(DB[4]), .R(w1161), .C(w1169), .nC(w1168) );
	vdp_slatch_r g1365 (.Q(w1485), .D(DB[1]), .R(w1161), .C(w1169), .nC(w1168) );
	vdp_slatch_r g1366 (.Q(w55), .D(DB[2]), .R(w1161), .C(w1169), .nC(w1168) );
	vdp_slatch_r g1367 (.Q(w43), .D(DB[0]), .R(w1161), .C(w1169), .nC(w1168) );
	vdp_comp_str g1368 (.Z(w1170), .nZ(w1166), .A(w1167) );
	vdp_notif0 g1369 (.A(VPOS[9]), .nZ(DB[10]), .nE(w1182) );
	vdp_notif0 g1370 (.A(VPOS[8]), .nZ(DB[9]), .nE(w1182) );
	vdp_bufif0 g1371 (.A(w587), .Z(DB[9]), .nE(w1213) );
	vdp_bufif0 g1372 (.A(w1033), .Z(DB[8]), .nE(w1213) );
	vdp_bufif0 g1373 (.A(w1212), .Z(DB[1]), .nE(w1213) );
	vdp_bufif0 g1374 (.A(w1214), .Z(DB[0]), .nE(w1213) );
	vdp_bufif0 g1375 (.A(w1195), .Z(DB[7]), .nE(w1213) );
	vdp_bufif0 g1376 (.A(w1194), .Z(DB[6]), .nE(w1213) );
	vdp_bufif0 g1377 (.A(w1193), .Z(DB[5]), .nE(w1213) );
	vdp_bufif0 g1378 (.A(ODD_EVEN), .Z(DB[4]), .nE(w1213) );
	vdp_bufif0 g1379 (.A(w46), .Z(DB[3]), .nE(w1213) );
	vdp_bufif0 g1380 (.A(w21), .Z(DB[2]), .nE(w1213) );
	vdp_slatch_r g1381 (.Q(w79), .D(DB[4]), .R(w1161), .C(w1163), .nC(w1162) );
	vdp_slatch_r g1382 (.Q(w80), .D(DB[5]), .R(w1161), .C(w1163), .nC(w1162) );
	vdp_slatch_r g1383 (.Q(w82), .D(DB[7]), .R(w1161), .C(w1163), .nC(w1162) );
	vdp_slatch_r g1384 (.Q(w81), .D(DB[6]), .R(w1161), .C(w1163), .nC(w1162) );
	vdp_slatch_r g1385 (.Q(w75), .D(DB[0]), .R(w1161), .C(w1163), .nC(w1162) );
	vdp_slatch_r g1386 (.Q(w76), .D(DB[1]), .R(w1161), .C(w1163), .nC(w1162) );
	vdp_slatch_r g1387 (.Q(w78), .D(DB[3]), .R(w1161), .C(w1163), .nC(w1162) );
	vdp_slatch_r g1388 (.Q(w77), .D(DB[2]), .R(w1161), .C(w1163), .nC(w1162) );
	vdp_notif0 g1389 (.A(HPOS[0]), .nZ(DB[8]), .nE(w1182) );
	vdp_not g1390 (.A(w403), .nZ(w1494) );
	vdp_comp_str g1391 (.Z(w1183), .A(w809), .nZ(w1186) );
	vdp_slatch_r g1392 (.Q(w1199), .D(w1184), .R(SYSRES), .C(w1183), .nC(w1186) );
	vdp_slatch_r g1393 (.Q(w1209), .D(w1190), .R(SYSRES), .C(w1183), .nC(w1186) );
	vdp_slatch_r g1394 (.Q(w1215), .D(w1185), .R(SYSRES), .C(w1183), .nC(w1186) );
	vdp_slatch_r g1395 (.Q(w1203), .D(w1484), .R(SYSRES), .C(w1183), .nC(w1186) );
	vdp_slatch_r g1396 (.Q(w1210), .D(w1177), .R(SYSRES), .C(w1183), .nC(w1186) );
	vdp_slatch_r g1397 (.Q(w1202), .D(w1174), .R(SYSRES), .C(w1183), .nC(w1186) );
	vdp_slatch_r g1398 (.Q(w1211), .D(w1176), .R(SYSRES), .C(w1183), .nC(w1186) );
	vdp_slatch_r g1399 (.Q(w1204), .D(w1189), .R(SYSRES), .C(w1183), .nC(w1186) );
	vdp_aon22 g1400 (.Z(w1212), .A1(w587), .A2(w1197), .B1(w1198), .B2(DMA_BUSY) );
	vdp_aon22 g1401 (.Z(w1214), .A1(w1033), .A2(w1197), .B1(w1198), .B2(PAL) );
	vdp_and3 g1402 (.C(w1187), .A(w406), .B(w1494), .Z(w1192) );
	vdp_not g1403 (.A(w1192), .nZ(w1182) );
	vdp_not g1404 (.A(w998), .nZ(w1213) );
	vdp_cnt_bit_load g1405 (.V(w1204), .nL(w1220), .L(w1200), .R(1'b0), .Q(w1221), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1249) );
	vdp_cnt_bit_load g1406 (.V(w1203), .nL(w1220), .L(w1200), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1526), .CO(w1249) );
	vdp_cnt_bit_load g1407 (.V(w1202), .nL(w1220), .L(w1200), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1248), .CO(w1526) );
	vdp_cnt_bit_load g1408 (.V(w1211), .nL(w1220), .L(w1200), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1247), .CO(w1248) );
	vdp_cnt_bit_load g1409 (.V(w1210), .nL(w1220), .L(w1200), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1246), .CO(w1247) );
	vdp_cnt_bit_load g1410 (.V(w1209), .nL(w1220), .L(w1200), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1536), .CO(w1246) );
	vdp_cnt_bit_load g1411 (.V(w1215), .nL(w1220), .L(w1200), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1245), .CO(w1536) );
	vdp_cnt_bit_load g1412 (.V(w1199), .nL(w1220), .L(w1200), .R(1'b0), .CI(w1217), .CO(w1245), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g1413 (.D(w1490), .C2(HCLK2), .C1(HCLK1), .Q(w1222), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_rs_ff g1414 (.Q(w1194), .R(w1238), .S(w1239) );
	vdp_rs_ff g1415 (.Q(w1195), .R(w1237), .S(w107) );
	vdp_rs_ff g1416 (.Q(w1193), .R(w1238), .S(w121) );
	vdp_not g1417 (.A(M5), .nZ(w1236) );
	vdp_not g1418 (.A(w1195), .nZ(w1216) );
	vdp_not g1419 (.A(w1201), .nZ(w1206) );
	vdp_not g1420 (.A(CA[21]), .nZ(w1491) );
	vdp_not g1421 (.A(w403), .nZ(w1207) );
	vdp_not g1422 (.A(w1241), .nZ(w1208) );
	vdp_comp_we g1423 (.Z(w1220), .A(w1489), .nZ(w1200) );
	vdp_or g1424 (.A(w1241), .B(w1222), .Z(w1489) );
	vdp_and g1425 (.A(w1208), .B(w1221), .Z(w1490) );
	vdp_and g1426 (.A(w1216), .B(w122), .Z(w1239) );
	vdp_or g1427 (.A(w1188), .B(w4), .Z(w1217) );
	vdp_not g1428 (.A(w1197), .nZ(w1198) );
	vdp_nor3 g1429 (.A(w403), .B(w1236), .Z(w1197), .C(CA[1]) );
	vdp_nor3 g1430 (.A(w1188), .B(w5), .Z(w1241), .C(w31) );
	vdp_nor g1431 (.A(w1244), .B(w1223), .Z(w1205) );
	vdp_or5 g1432 (.A(w1207), .B(CA[4]), .C(CA[5]), .D(CA[15]), .Z(w1244), .E(CA[6]) );
	vdp_or5 g1433 (.A(CA[16]), .B(CA[17]), .C(CA[20]), .D(w1206), .Z(w1223), .E(w1491) );
	vdp_rs_ff g1434 (.Q(w1229), .R(w1281), .S(w1490) );
	vdp_rs_ff g1435 (.Q(w1282), .R(w1265), .S(w1492) );
	vdp_dff g1436 (.Q(w1285), .R(w1242), .C(w1232), .D(w1225) );
	vdp_dff g1437 (.Q(w1284), .R(w1242), .C(w1232), .D(w1224) );
	vdp_dff g1438 (.Q(w1286), .R(w1242), .C(w1232), .D(w1226) );
	vdp_rs_ff g1439 (.Q(w1542), .R(w1280), .S(w1541) );
	vdp_rs_ff g1440 (.Q(w1253), .R(w1254), .S(w1539) );
	vdp_dlatch_inv g1441 (.D(w1260), .Q(w1261), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g1442 (.D(w1254), .C(DCLK1), .Q(w1260), .nC(nDCLK1) );
	vdp_dlatch_inv g1443 (.D(w1263), .Q(w1238), .C(HCLK1), .nC(nHCLK1) );
	vdp_not g1444 (.A(w1276), .nZ(w1250) );
	vdp_not g1445 (.A(w668), .nZ(w1228) );
	vdp_not g1446 (.A(w1231), .nZ(w1226) );
	vdp_not g1447 (.A(w1230), .nZ(w1225) );
	vdp_not g1448 (.A(w1240), .nZ(w1242) );
	vdp_not g1449 (.A(w1257), .nZ(w1232) );
	vdp_not g1450 (.A(w1233), .nZ(w50) );
	vdp_not g1451 (.A(w1235), .nZ(w1234) );
	vdp_sr_bit g1452 (.D(w1262), .C2(HCLK2), .C1(HCLK1), .Q(w1280), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and g1453 (.A(M5), .B(w1253), .Z(w1257) );
	vdp_and g1454 (.A(w403), .B(w1252), .Z(w1075) );
	vdp_and g1455 (.A(w1233), .B(w1075), .Z(w1540) );
	vdp_or g1456 (.A(w1016), .B(w1540), .Z(w1539) );
	vdp_or g1457 (.A(w998), .B(SYSRES), .Z(w1541) );
	vdp_and g1458 (.A(w1236), .B(w1238), .Z(w1264) );
	vdp_or g1459 (.A(w1284), .B(w1264), .Z(w1265) );
	vdp_and g1460 (.A(M5), .B(w469), .Z(w1492) );
	vdp_and g1461 (.A(w1140), .B(M5), .Z(w1227) );
	vdp_or g1462 (.A(w1286), .B(w1264), .Z(w1237) );
	vdp_or g1463 (.A(w1285), .B(w1264), .Z(w1281) );
	vdp_comp_dff g1464 (.D(w1542), .C2(HCLK2), .C1(HCLK1), .Q(w1262), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_comp_dff g1465 (.D(w1257), .C2(DCLK2), .C1(DCLK1), .Q(w1254), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_nor g1466 (.A(w1262), .B(SYSRES), .Z(w1564) );
	vdp_nand g1467 (.A(w1280), .B(w1564), .Z(w1263) );
	vdp_nand g1468 (.A(w1195), .B(w1139), .Z(w1231) );
	vdp_and3 g1469 (.A(w1227), .B(w925), .Z(w1275), .C(w1228) );
	vdp_and3 g1470 (.A(w1227), .B(w925), .Z(w1274), .C(w668) );
	vdp_and4 g1471 (.A(w1230), .B(w1138), .C(w1231), .D(w1282), .Z(w1224) );
	vdp_nand3 g1472 (.C(w1229), .A(w1231), .B(w1172), .Z(w1230) );
	vdp_aoi21 g1473 (.A1(w1261), .B(SYSRES), .Z(w1240), .A2(w1260) );
	vdp_dff g1474 (.Q(w1305), .R(w1291), .C(w1288), .D(w1273) );
	vdp_dff g1475 (.Q(w1301), .R(w1291), .C(w1288), .D(w1300) );
	vdp_dff g1476 (.Q(w1270), .R(w1291), .C(w1288), .D(w1268) );
	vdp_dff g1477 (.Q(w1278), .R(w1291), .C(w1288), .D(w1277) );
	vdp_dff g1478 (.Q(w1279), .R(w1291), .C(w1288), .D(w1267) );
	vdp_dff g1479 (.Q(w1258), .R(w1291), .C(w1288), .D(w1296) );
	vdp_dff g1480 (.Q(w1255), .R(w1291), .C(w1288), .D(w1294) );
	vdp_dff g1481 (.Q(w1287), .R(1'b0), .C(w1288), .D(w1251) );
	vdp_ha g1482 (.SUM(w1294), .A(w1255), .B(w1250), .CO(w1256) );
	vdp_ha g1483 (.SUM(w1296), .A(w1258), .B(w1256), .CO(w1259) );
	vdp_ha g1484 (.SUM(w1267), .A(w1279), .B(w1259), .CO(w1266) );
	vdp_ha g1485 (.SUM(w1277), .A(w1278), .B(w1266), .CO(w1271) );
	vdp_ha g1486 (.SUM(w1268), .A(w1270), .B(w1271), .CO(w1269) );
	vdp_ha g1487 (.SUM(w1273), .A(w1305), .B(w1269), .CO(w1272) );
	vdp_ha g1488 (.SUM(w1300), .A(w1301), .B(w1272) );
	vdp_and3 g1489 (.A(w1301), .B(w1270), .Z(w1298), .C(w1305) );
	vdp_and4 g1490 (.C(w1258), .A(w1278), .B(w1298), .Z(w1304), .D(w1279) );
	vdp_nand g1491 (.A(w1287), .B(w403), .Z(w1428) );
	vdp_dff g1492 (.Q(w1313), .R(1'b0), .C(w1288), .D(w1293) );
	vdp_dff g1493 (.Q(w1293), .R(w1295), .C(w1288), .D(w1318) );
	vdp_dff g1494 (.Q(w1318), .R(w1295), .C(w1316), .D(w1297) );
	vdp_dff g1495 (.Q(w1297), .R(w1295), .C(w1288), .D(w1322) );
	vdp_dff g1496 (.Q(w1322), .R(w1295), .C(w1288), .D(w1323) );
	vdp_dff g1497 (.Q(w1323), .R(w1295), .C(w1288), .D(1'b1) );
	vdp_dff g1498 (.Q(w1529), .R(w1332), .C(w1306), .D(w1298) );
	vdp_dff g1499 (.Q(w1306), .R(1'b0), .C(w1288), .D(w1304) );
	vdp_dff g1500 (.Q(w1325), .R(w1303), .C(w1326), .D(w1298) );
	vdp_dff g1501 (.Q(w1302), .R(w1317), .C(w1330), .D(1'b1) );
	vdp_or g1502 (.A(SYSRES), .B(w1302), .Z(w1303) );
	vdp_or g1503 (.A(w1295), .B(w1313), .Z(w1328) );
	vdp_not g1504 (.A(w1313), .nZ(w1290) );
	vdp_not g1505 (.A(w1529), .nZ(w1295) );
	vdp_nand3 g1506 (.A(w403), .B(w1311), .Z(w1291), .C(w1290) );
	vdp_not g1507 (.nZ(w1316), .A(w1312) );
	vdp_not g1508 (.nZ(w1288), .A(w1289) );
	vdp_dff g1509 (.Q(w1315), .R(1'b0), .C(w1316), .D(w1338) );
	vdp_dff g1510 (.Q(w1341), .R(w1317), .C(w1316), .D(w1321) );
	vdp_dff g1511 (.Q(w1321), .R(w1317), .C(w1288), .D(w1343) );
	vdp_dff g1512 (.Q(w1343), .R(w1317), .C(w1316), .D(w1320) );
	vdp_dff g1513 (.Q(w1320), .R(w1317), .C(w1316), .D(w1331) );
	vdp_dff g1514 (.Q(w1331), .R(w1317), .C(w1288), .D(w47) );
	vdp_dff g1515 (.Q(w1348), .R(w1347), .C(w1316), .D(w1128) );
	vdp_dff g1516 (.Q(w1128), .R(w1347), .C(w1288), .D(w1327) );
	vdp_not g1517 (.A(w1335), .nZ(w108) );
	vdp_not g1518 (.A(w996), .nZ(w1310) );
	vdp_not g1519 (.A(w1321), .nZ(w1319) );
	vdp_not g1520 (.A(w1318), .nZ(w1537) );
	vdp_not g1521 (.A(w1327), .nZ(w1347) );
	vdp_not g1522 (.A(w1075), .nZ(w1330) );
	vdp_not g1523 (.A(w1233), .nZ(w1530) );
	vdp_and g1524 (.A(w1328), .B(w1075), .Z(w1327) );
	vdp_and g1525 (.A(w1329), .B(w1327), .Z(w1326) );
	vdp_and g1526 (.A(w1348), .B(w1326), .Z(w47) );
	vdp_and g1527 (.A(w1322), .B(w1537), .Z(w1339) );
	vdp_and g1528 (.A(w1323), .B(w1537), .Z(w1340) );
	vdp_and g1529 (.A(w1314), .B(w987), .Z(w1337) );
	vdp_and g1530 (.A(w1314), .B(w1030), .Z(w1309) );
	vdp_and g1531 (.A(w996), .B(w1315), .Z(w1314) );
	vdp_and g1532 (.A(w108), .B(w1128), .Z(w1063) );
	vdp_nand g1533 (.A(w1320), .B(w1319), .Z(w1311) );
	vdp_nor g1534 (.A(w1317), .B(w1331), .Z(w1342) );
	vdp_or3 g1535 (.C(w1325), .A(SYSRES), .B(w1313), .Z(w1332) );
	vdp_oai21 g1536 (.A1(w1030), .B(w1310), .Z(w1335), .A2(w987) );
	vdp_dff g1537 (.Q(w1356), .R(1'b0), .C(w1288), .D(w1235) );
	vdp_rs_ff g1538 (.nQ(w1072), .R(w1357), .S(w1354) );
	vdp_not g1539 (.A(w1362), .nZ(PSG_Z80_CLK) );
	vdp_not g1540 (.A(REG_BUS[7]), .nZ(w1353) );
	vdp_and3 g1541 (.C(w1353), .A(w825), .B(M5), .Z(w1354) );
	vdp_or g1542 (.A(w1235), .B(SYSRES), .Z(w1357) );
	vdp_and g1543 (.A(w1374), .B(w588), .Z(w1375) );
	vdp_not g1544 (.A(w1329), .nZ(w1377) );
	vdp_and4 g1545 (.C(CA[21]), .A(w1201), .B(CA[20]), .Z(w1329), .D(w1530) );
	vdp_dff g1546 (.Q(w1417), .R(1'b0), .C(w1362), .D(w1402) );
	vdp_dff g1547 (.Q(w1397), .R(1'b0), .C(w1362), .D(w1396) );
	vdp_dff g1548 (.Q(w1336), .R(1'b0), .C(w1383), .D(w1384) );
	vdp_dff g1549 (.Q(w1396), .R(1'b0), .C(w1383), .D(w1336) );
	vdp_dff g1550 (.Q(w1409), .R(w1410), .C(HCLK2), .D(w1412) );
	vdp_dff g1551 (.Q(DMA_BUSY), .R(w1410), .C(HCLK2), .D(w1409) );
	vdp_rs_ff g1552 (.Q(w1276), .R(w1410), .S(w1345) );
	vdp_rs_ff g1553 (.Q(w1531), .R(w1410), .S(w1274) );
	vdp_rs_ff g1554 (.Q(w1251), .R(w1346), .S(w1275) );
	vdp_sr_bit g1555 (.D(w588), .Q(w1374), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1556 (.D(w1538), .Q(w1408), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_dlatch_inv g1557 (.D(w1373), .nQ(w1351), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g1558 (.D(w1372), .nQ(w1373), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g1559 (.D(w1359), .C(HCLK1), .nQ(w1372), .nC(nHCLK1) );
	vdp_aon22 g1560 (.Z(w1404), .A2(w1350), .B1(w1372), .B2(w1413), .A1(w1351) );
	vdp_sr_bit g1561 (.D(w1414), .Q(w1419), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1562 (.D(w1376), .Q(w1414), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1563 (.D(VRAM_REFRESH), .C2(HCLK2), .C1(HCLK1), .Q(w1376), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_aon22 g1564 (.Z(w1392), .A2(w1342), .B1(w1420), .B2(w1423), .A1(w1390) );
	vdp_not g1565 (.A(w1528), .nZ(w1065) );
	vdp_not g1566 (.A(w1342), .nZ(w1423) );
	vdp_not g1567 (.A(w1408), .nZ(w1413) );
	vdp_not g1568 (.A(w1349), .nZ(w1391) );
	vdp_not g1569 (.A(w1325), .nZ(w1317) );
	vdp_or g1570 (.A(w1276), .B(w1531), .Z(w1412) );
	vdp_or g1571 (.A(SYSRES), .B(w590), .Z(w1410) );
	vdp_or g1572 (.A(w1345), .B(w1410), .Z(w1346) );
	vdp_or g1573 (.A(w1226), .B(w1224), .Z(w277) );
	vdp_or g1574 (.A(w1226), .B(w1225), .Z(w252) );
	vdp_and g1575 (.A(w1408), .B(w642), .Z(w1350) );
	vdp_or g1576 (.A(w1351), .B(w1414) );
	vdp_and g1577 (.A(w1311), .B(w1326), .Z(w1390) );
	vdp_and g1578 (.A(w1343), .B(w1326), .Z(w1420) );
	vdp_and g1579 (.A(w1326), .B(w1317), .Z(w110) );
	vdp_and g1580 (.A(w991), .B(w111), .Z(w1403) );
	vdp_or g1581 (.A(w1337), .B(w995), .Z(w1399) );
	vdp_aon22 g1582 (.Z(w1407), .A2(w1066), .B1(w1344), .B2(w1395), .A1(w1394) );
	vdp_and g1583 (.A(w1402), .B(w1417), .Z(w1127) );
	vdp_and g1584 (.A(w1415), .B(w1424), .Z(w1405) );
	vdp_and g1585 (.A(w1424), .B(w1418), .Z(w1402) );
	vdp_not g1586 (.A(w1418), .nZ(w1415) );
	vdp_not g1587 (.A(w1416), .nZ(w1424) );
	vdp_not g1588 (.A(w1373), .nZ(w1411) );
	vdp_not g1589 (.A(w1388), .nZ(w1406) );
	vdp_and g1590 (.A(w1400), .B(w1364), .Z(w1363) );
	vdp_and g1591 (.A(w1400), .B(w1366), .Z(w990) );
	vdp_and g1592 (.A(w1400), .B(w1368), .Z(w995) );
	vdp_and g1593 (.A(w1400), .B(w1365), .Z(w991) );
	vdp_and g1594 (.A(w1400), .B(w1367), .Z(w1384) );
	vdp_and g1595 (.A(w990), .B(w1384), .Z(w1016) );
	vdp_and g1596 (.A(w403), .B(w1378), .Z(w987) );
	vdp_and g1597 (.A(w403), .B(w1369), .Z(w1030) );
	vdp_not g1598 (.A(w403), .nZ(w1400) );
	vdp_nand g1599 (.A(w1396), .B(w1397), .Z(w1418) );
	vdp_nand g1600 (.A(w1033), .B(w1361), .Z(w1360) );
	vdp_nand g1601 (.A(w403), .B(w252), .Z(w1371) );
	vdp_nand g1602 (.A(w277), .B(w403), .Z(w1370) );
	vdp_or3 g1603 (.C(w1226), .A(w1225), .B(w1224), .Z(w1058) );
	vdp_and3 g1604 (.C(w1351), .A(w588), .B(w1408), .Z(w593) );
	vdp_aoi21 g1605 (.A2(w1350), .B(w1411), .Z(w1349), .A1(w1372) );
	vdp_nor g1606 (.A(w1376), .B(w1419), .Z(w1361) );
	vdp_nand g1607 (.A(w108), .B(w1377), .Z(w1388) );
	vdp_nand3 g1608 (.C(w1360), .A(w3), .B(w1375), .Z(w1359) );
	vdp_2a3oi g1609 (.A1(w1411), .B(w669), .Z(w1358), .A2(w1372), .C(w1408) );
	vdp_nor4 g1610 (.C(VRAM_REFRESH), .A(w1414), .B(w1376), .Z(w1538), .D(w1419) );
	vdp_comb1 g1611 (.A1(CA[15]), .B(w1415), .Z(w1416), .A2(CA[14]), .C(w1363) );
	vdp_aon22 g1612 (.Z(w1334), .A2(w1066), .B1(w1344), .B2(w1389), .A1(w1527) );
	vdp_not g1613 (.A(w1066), .nZ(w1344) );
	vdp_or4 g1614 (.C(w1391), .A(w1424), .B(w1390), .Z(w1527), .D(w1339) );
	vdp_or4 g1615 (.C(w1351), .A(w1406), .B(w1403), .Z(w1395), .D(w1351) );
	vdp_or3 g1616 (.C(w1392), .A(w1402), .B(w1393), .Z(w1389) );
	vdp_comb1 g1617 (.A1(w1128), .B(w1321), .Z(w1528), .A2(w1342), .C(w1326) );
	vdp_and6 g1618 (.C(w1386), .A(w1287), .B(w1385), .Z(w1345), .D(w1356), .E(w403), .F(w1330) );
	vdp_or5 g1619 (.C(w1404), .A(w1396), .B(w47), .Z(w1394), .D(w1340), .E(w1129) );
	vdp_or5 g1620 (.C(w1351), .A(w1405), .B(w109), .Z(w1398), .D(w1339), .E(w1403) );
	vdp_aoi22 g1621 (.Z(w1338), .A2(w47), .B1(w1341), .B2(w1326), .A1(w1342) );
	vdp_n_fet g1622 (.Z(w305), .A(w423) );
	vdp_n_fet g1623 (.Z(w262), .A(w423) );
	vdp_n_fet g1624 (.A(w423), .Z(w297) );
	vdp_n_fet g1625 (.A(w423), .Z(w254) );
	vdp_n_fet g1626 (.Z(w288), .A(w423) );
	vdp_n_fet g1627 (.Z(w245), .A(w423) );
	vdp_n_fet g1628 (.Z(w279), .A(w423) );
	vdp_n_fet g1629 (.Z(w237), .A(w423) );
	vdp_aon22 g1630 (.Z(w1393), .A2(w1350), .B1(w1350), .B2(w1411), .A1(w1351) );
	vdp_comp_we g1631 (.nZ(w1362), .Z(w1383), .A(w1401) );
	vdp_comp_we g1632 (.nZ(w1289), .Z(w1312), .A(w1429) );
	vdp_not g1633 (.nZ(w1619), .A(w1973) );
	vdp_not g1634 (.nZ(w1621), .A(w1622) );
	vdp_sr_bit g1635 (.Q(w5), .D(w1968), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1636 (.Q(w1627), .D(w1823), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1637 (.Q(w1603), .D(w1824), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1638 (.Q(w1659), .D(w1624), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1639 (.Q(w1604), .D(w1825), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1640 (.Q(w1608), .D(w1826), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1641 (.Q(w1801), .D(w1813), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1642 (.Q(w1635), .D(w1633), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1643 (.Q(w1632), .D(w1814), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1644 (.Q(w1609), .D(w1815), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1645 (.Q(w1642), .D(w1840), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1646 (.Q(w1640), .D(w1637), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1647 (.Q(w1637), .D(w1984), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1648 (.Q(w1641), .D(w1644), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1649 (.Q(w1614), .D(w1934), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_not g1650 (.nZ(w1633), .A(w1643) );
	vdp_not g1651 (.nZ(w58), .A(w1632) );
	vdp_not g1652 (.nZ(w1618), .A(w1632) );
	vdp_not g1653 (.nZ(w1611), .A(ODD_EVEN) );
	vdp_not g1654 (.nZ(w1620), .A(LS0) );
	vdp_not g1655 (.nZ(w1984), .A(w1969) );
	vdp_not g1656 (.nZ(w1646), .A(w1647) );
	vdp_not g1657 (.nZ(w1634), .A(w1970) );
	vdp_not g1658 (.nZ(w1639), .A(w1640) );
	vdp_not g1659 (.nZ(w1616), .A(w53) );
	vdp_and g1660 (.Z(w1638), .A(w1836), .B(w1642) );
	vdp_nor g1661 (.Z(w1636), .A(SYSRES), .B(w1608) );
	vdp_oai21 g1662 (.Z(w1969), .B(w1636), .A2(w1646), .A1(w1637) );
	vdp_oai21 g1663 (.Z(w1647), .B(w1645), .A2(w1644), .A1(w1840) );
	vdp_aoi21 g1664 (.Z(w1970), .B(SYSRES), .A2(w1641), .A1(w1836) );
	vdp_and g1665 (.Z(w1615), .A(w1618), .B(w27) );
	vdp_and3 g1666 (.Z(w1836), .A(w1639), .B(w53), .C(w1637) );
	vdp_or g1667 (.Z(w1617), .A(SYSRES), .B(w1618) );
	vdp_and g1668 (.Z(w1934), .A(w1612), .B(w1622) );
	vdp_and g1669 (.Z(w1623), .A(w1615), .B(w1616) );
	vdp_and g1670 (.Z(w1612), .A(w1615), .B(w53) );
	vdp_and g1671 (.Z(w1607), .A(w1602), .B(w1609) );
	vdp_or g1672 (.Z(w1606), .A(SYSRES), .B(w1607) );
	vdp_2A3OI g1673 (.Z(w1973), .A1(w1621), .A2(w1612), .C(SYSRES), .B(w1620) );
	vdp_or g1674 (.Z(w1602), .A(w1610), .B(w1611) );
	vdp_or g1675 (.Z(w1605), .A(SYSRES), .B(w1657) );
	vdp_and g1676 (.Z(w1657), .A(w1602), .B(w1604) );
	vdp_and g1677 (.Z(w1628), .A(w1602), .B(w1627) );
	vdp_and g1678 (.Z(w1626), .A(w1602), .B(w1603) );
	vdp_or g1679 (.Z(w1924), .A(w1657), .B(SYSRES) );
	vdp_and g1680 (.Z(w1842), .A(w1624), .B(M5) );
	vdp_not g1681 (.nZ(w46), .A(w1630) );
	vdp_not g1682 (.nZ(w1630), .A(w1629) );
	vdp_not g1683 (.nZ(w1663), .A(w1629) );
	vdp_not g1684 (.nZ(w1968), .A(w1812) );
	vdp_and g1685 (.Z(w1729), .A(M5), .B(w1625) );
	vdp_or g1686 (.Z(w1631), .A(SYSRES), .B(w1628) );
	vdp_oai21 g1687 (.Z(w1629), .B(w1110), .A2(w31), .A1(w5) );
	vdp_rs_ff g1688 (.Q(w1625), .S(w1626), .R(w1631) );
	vdp_rs_ff g1689 (.Q(w1613), .R(w1605), .S(w1607) );
	vdp_rs_ff g1690 (.Q(w31), .S(w1635), .R(w1617) );
	vdp_rs_ff g1691 (.Q(w20), .R(w1608), .S(w1606) );
	vdp_tff g1692 (.C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .CI(w1623), .R(w1619), .A(w1614), .Q(ODD_EVEN) );
	vdp_cnt_bit_load g1693 (.D(w1832), .Q(w1695), .nL(w1951), .L(w1817), .CI(w1834), .nC1(nHCLK1), .CO(w1922), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g1694 (.Q(w1610), .D(w1913), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1695 (.Q(w1982), .D(w1931), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1696 (.Q(w32), .D(w1997), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1697 (.Q(w27), .D(w1909), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1698 (.Q(VRAM_REFRESH), .D(w1682), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1699 (.Q(w1697), .D(w1681), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1700 (.Q(w1691), .D(w1680), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1701 (.Q(w1667), .D(w1910), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1702 (.Q(w1692), .D(w1706), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1703 (.Q(w1644), .D(w1912), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1704 (.Q(w1839), .D(w1914), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1705 (.Q(w1721), .D(w1908), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1706 (.Q(w1840), .D(w1904), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1707 (.Q(w1706), .D(w1961), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1708 (.Q(w1858), .D(w1866), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1709 (.Q(w1701), .D(w1678), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1710 (.Q(w1720), .D(w1867), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1711 (.Q(w1995), .D(w1999), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1712 (.Q(w1753), .D(w1749), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1713 (.Q(w1703), .D(w1861), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1714 (.Q(w9), .D(w1860), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1715 (.Q(w1718), .D(w1763), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1716 (.Q(w1715), .D(w1911), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1717 (.Q(w1734), .D(w1865), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1718 (.Q(w1726), .D(w1740), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1719 (.Q(w1784), .D(w1730), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1720 (.Q(w29), .D(w1755), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1721 (.Q(w22), .D(w1664), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1722 (.Q(w1748), .D(w1762), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1723 (.Q(w1963), .D(w1790), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1724 (.Q(w1786), .D(w1862), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1725 (.Q(w1744), .D(w1902), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1726 (.Q(w1770), .D(w1793), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1727 (.Q(w30), .D(w1933), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1728 (.Q(w1772), .D(w1864), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1729 (.Q(w1773), .D(w1863), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1730 (.Q(w1799), .D(w1742), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1731 (.Q(w1745), .D(w1905), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1732 (.Q(w1658), .D(w1989), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1733 (.Q(w1732), .D(w1988), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1734 (.Q(w1785), .D(w1741), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1735 (.Q(w1746), .D(w1743), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1736 (.Q(w1789), .D(w1906), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1737 (.Q(w1767), .D(w1903), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1738 (.Q(w25), .D(w1665), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1739 (.Q(w1768), .D(w1658), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1740 (.Q(w1800), .D(w1754), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1741 (.Q(w1852), .D(w1901), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_not g1742 (.nZ(w1687), .A(M5) );
	vdp_not g1743 (.nZ(w6), .A(w1936) );
	vdp_not g1744 (.nZ(w7), .A(w1667) );
	vdp_not g1745 (.nZ(w1859), .A(w1662) );
	vdp_not g1746 (.nZ(w1671), .A(w53) );
	vdp_not g1747 (.nZ(w1673), .A(w1932) );
	vdp_not g1748 (.nZ(w1759), .A(w1) );
	vdp_not g1749 (.nZ(w1711), .A(w1679) );
	vdp_not g1750 (.nZ(w1693), .A(w1692) );
	vdp_not g1751 (.nZ(w1704), .A(w1667) );
	vdp_not g1752 (.nZ(w1705), .A(w44) );
	vdp_not g1753 (.nZ(w8), .A(w1699) );
	vdp_not g1754 (.nZ(w1689), .A(w39) );
	vdp_not g1755 (.nZ(w1994), .A(w53) );
	vdp_not g1756 (.nZ(w13), .A(w1957) );
	vdp_not g1757 (.nZ(w1958), .A(w1715) );
	vdp_not g1758 (.nZ(w1961), .A(w1725) );
	vdp_not g1759 (.nZ(w1758), .A(w1684) );
	vdp_not g1760 (.nZ(w1980), .A(w1683) );
	vdp_not g1761 (.nZ(w1709), .A(H40) );
	vdp_not g1762 (.nZ(w14), .A(w1756) );
	vdp_not g1763 (.nZ(w1950), .A(w1670) );
	vdp_not g1764 (.nZ(w1796), .A(w1728) );
	vdp_not g1765 (.nZ(w1774), .A(w1760) );
	vdp_not g1766 (.nZ(w1791), .A(w52) );
	vdp_not g1767 (.nZ(w1736), .A(w1907) );
	vdp_not g1768 (.nZ(w12), .A(w1937) );
	vdp_not g1769 (.nZ(w1802), .A(w1800) );
	vdp_not g1770 (.nZ(w1702), .A(w42) );
	vdp_not g1771 (.nZ(w1719), .A(w51) );
	vdp_not g1772 (.nZ(w1668), .A(w41) );
	vdp_not g1773 (.nZ(w1923), .A(w19) );
	vdp_not g1774 (.nZ(w1981), .A(w45) );
	vdp_not g1775 (.nZ(w1983), .A(M5) );
	vdp_not g1776 (.nZ(w1976), .A(w1737) );
	vdp_not g1777 (.nZ(w1816), .A(w1765) );
	vdp_not g1778 (.nZ(w1954), .A(w1930) );
	vdp_not g1779 (.nZ(w1818), .A(w1086) );
	vdp_not g1780 (.nZ(w1835), .A(w1833) );
	vdp_not g1781 (.nZ(w1829), .A(w1487) );
	vdp_not g1782 (.nZ(w1830), .A(PAL) );
	vdp_aon22 g1783 (.Z(w2004), .B1(w1820), .A1(w1819), .A2(DB[4]), .B2(w1818) );
	vdp_aon22 g1784 (.Z(w1943), .B1(w1820), .A1(w1819), .A2(DB[5]), .B2(w1806) );
	vdp_aon22 g1785 (.Z(w1944), .B1(w1820), .A1(w1819), .B2(w1954), .A2(DB[6]) );
	vdp_aon22 g1786 (.Z(w1940), .B2(1'b1), .A2(DB[7]), .B1(w1820), .A1(w1819) );
	vdp_aon22 g1787 (.Z(w1939), .B2(1'b1), .A2(DB[8]), .B1(w1820), .A1(w1819) );
	vdp_aon22 g1788 (.Z(w1809), .B2(1'b1), .B1(w1669), .A2(DB[8]), .A1(w1998) );
	vdp_aon22 g1789 (.Z(w1953), .B2(w1805), .A2(DB[3]), .B1(w1820), .A1(w1819) );
	vdp_aon22 g1790 (.Z(w1827), .A2(DB[2]), .B2(w1830), .B1(w1820), .A1(w1819) );
	vdp_aon22 g1791 (.Z(w1828), .A2(DB[1]), .B2(w1804), .B1(w1820), .A1(w1819) );
	vdp_aon22 g1792 (.Z(w1945), .A1(w1998), .B1(w1669), .B2(1'b1), .A2(DB[7]) );
	vdp_aon22 g1793 (.Z(w21), .A1(w1983), .B2(w1807), .B1(M5), .A2(w1784) );
	vdp_aon22 g1794 (.Z(w1777), .B1(w1669), .A1(w1998), .A2(DB[6]), .B2(1'b1) );
	vdp_aon22 g1795 (.Z(w1752), .B1(w1768), .B2(w1769), .A2(w1853), .A1(w1766) );
	vdp_not g1796 (.nZ(w1769), .A(w1766) );
	vdp_aon22 g1797 (.Z(w1946), .B1(w1669), .A1(w1998), .B2(1'b0), .A2(DB[5]) );
	vdp_not g1798 (.nZ(w1797), .A(w1794) );
	vdp_aon22 g1799 (.Z(w1990), .B1(w1669), .A1(w1998), .B2(w1950), .A2(DB[4]) );
	vdp_aon22 g1800 (.Z(w1947), .B2(w1949), .B1(w1669), .A2(DB[3]), .A1(w1998) );
	vdp_aon22 g1801 (.Z(w1750), .A2(w1687), .B2(M5), .A1(w1752), .B1(w1751) );
	vdp_aon22 g1802 (.Z(w1948), .A2(DB[2]), .B2(w1722), .A1(w1998), .B1(w1669) );
	vdp_aon22 g1803 (.Z(w1959), .B2(w1858), .B1(w44), .A2(w1705), .A1(w1704) );
	vdp_aon22 g1804 (.Z(w1696), .B1(w1935), .A1(HCLK2), .B2(w1689), .A2(w39) );
	vdp_aon22 g1805 (.Z(w1974), .A1(w1998), .B1(w1669), .B2(w1707), .A2(DB[1]) );
	vdp_aon22 g1806 (.Z(w1674), .A2(DB[0]), .B1(w1669), .B2(w1670), .A1(w1998) );
	vdp_not g1807 (.nZ(w4), .A(w1839) );
	vdp_not g1808 (.nZ(w3), .A(w1703) );
	vdp_rs_ff g1809 (.Q(w1747), .S(w1798), .R(w1926) );
	vdp_rs_ff g1810 (.Q(w1795), .R(w1786), .S(w1788) );
	vdp_rs_ff g1811 (.Q(w1730), .S(w1964), .R(w1746) );
	vdp_rs_ff g1812 (.Q(w1925), .R(w1993), .S(w1726) );
	vdp_rs_ff g1813 (.Q(w1731), .R(w1721), .S(w1987) );
	vdp_aon22 g1814 (.Z(w1832), .A2(DB[0]), .B2(w1803), .B1(w1820), .A1(w1819) );
	vdp_notif0 g1815 (.nZ(DB[1]), .A(VRAM_REFRESH), .nE(w1685) );
	vdp_notif0 g1816 (.nZ(DB[0]), .A(w32), .nE(w1685) );
	vdp_notif0 g1817 (.nZ(DB[7]), .A(w27), .nE(w1686) );
	vdp_notif0 g1818 (.A(w7), .nZ(DB[6]), .nE(w1686) );
	vdp_notif0 g1819 (.A(w6), .nZ(DB[2]), .nE(w1685) );
	vdp_notif0 g1820 (.A(w8), .nZ(DB[3]), .nE(w1685) );
	vdp_notif0 g1821 (.nZ(DB[5]), .A(w14), .nE(w1685) );
	vdp_notif0 g1822 (.A(w13), .nZ(DB[4]), .nE(w1685) );
	vdp_notif0 g1823 (.A(w16), .nZ(DB[5]), .nE(w1686) );
	vdp_notif0 g1824 (.nZ(DB[7]), .A(w9), .nE(w1685) );
	vdp_notif0 g1825 (.nZ(DB[6]), .A(w3), .nE(w1685) );
	vdp_notif0 g1826 (.nZ(DB[4]), .A(w17), .nE(w1686) );
	vdp_notif0 g1827 (.nZ(DB[9]), .A(w29), .nE(w1685) );
	vdp_notif0 g1828 (.nZ(DB[8]), .A(w22), .nE(w1685) );
	vdp_notif0 g1829 (.nZ(DB[3]), .A(w11), .nE(w1686) );
	vdp_notif0 g1830 (.nZ(DB[2]), .A(w28), .nE(w1686) );
	vdp_notif0 g1831 (.nZ(DB[10]), .A(w30), .nE(w1685) );
	vdp_notif0 g1832 (.nZ(DB[11]), .A(w12), .nE(w1685) );
	vdp_notif0 g1833 (.nZ(DB[12]), .A(w24), .nE(w1685) );
	vdp_notif0 g1834 (.nZ(DB[13]), .A(w25), .nE(w1685) );
	vdp_notif0 g1835 (.nZ(DB[1]), .A(w15), .nE(w1686) );
	vdp_notif0 g1836 (.nZ(DB[0]), .A(w10), .nE(w1686) );
	vdp_not g1837 (.nZ(VPOS[9]), .A(w1942) );
	vdp_not g1838 (.nZ(VPOS[8]), .A(w1941) );
	vdp_not g1839 (.nZ(VPOS[7]), .A(w1738) );
	vdp_not g1840 (.nZ(HPOS[7]), .A(w1976) );
	vdp_not g1841 (.nZ(HPOS[8]), .A(w1816) );
	vdp_not g1842 (.nZ(HPOS[6]), .A(w1736) );
	vdp_not g1843 (.nZ(VPOS[6]), .A(w1977) );
	vdp_not g1844 (.nZ(VPOS[5]), .A(w1978) );
	vdp_not g1845 (.nZ(HPOS[5]), .A(w1774) );
	vdp_not g1846 (.nZ(HPOS[4]), .A(w1796) );
	vdp_not g1847 (.nZ(VPOS[4]), .A(w1979) );
	vdp_not g1848 (.nZ(HPOS[3]), .A(w1980) );
	vdp_not g1849 (.nZ(VPOS[3]), .A(w1723) );
	vdp_not g1850 (.nZ(HPOS[2]), .A(w1758) );
	vdp_not g1851 (.nZ(VPOS[2]), .A(w1712) );
	vdp_not g1852 (.nZ(HPOS[1]), .A(w1711) );
	vdp_not g1853 (.nZ(VPOS[1]), .A(w1672) );
	vdp_not g1854 (.nZ(HPOS[0]), .A(w1673) );
	vdp_not g1855 (.nZ(VPOS[0]), .A(w1666) );
	vdp_aoi22 g1856 (.Z(w1935), .A1(w1659), .B1(w1688), .B2(M5), .A2(w1687) );
	vdp_aon22 g1857 (.Z(w1713), .A2(w1687), .B1(w1714), .B2(M5), .A1(w1754) );
	vdp_aoi22 g1858 (.Z(w1666), .B2(w1759), .B1(w1695), .A1(ODD_EVEN), .A2(w1) );
	vdp_aoi22 g1859 (.Z(w1672), .B2(w1759), .B1(w1837), .A1(w1695), .A2(w1) );
	vdp_aoi22 g1860 (.Z(w1712), .A2(w1), .A1(w1837), .B2(w1759), .B1(w1929) );
	vdp_aoi22 g1861 (.Z(w1723), .A1(w1929), .B2(w1759), .A2(w1), .B1(w1822) );
	vdp_aoi22 g1862 (.Z(w1979), .B1(w1928), .A1(w1822), .A2(w1), .B2(w1759) );
	vdp_aoi22 g1863 (.Z(w1978), .B1(w1776), .A1(w1928), .A2(w1), .B2(w1759) );
	vdp_aoi22 g1864 (.Z(w1977), .A2(w1), .B2(w1759), .B1(w1739), .A1(w1776) );
	vdp_aoi22 g1865 (.Z(w1738), .B2(w1759), .A1(w1739), .B1(w1811), .A2(w1) );
	vdp_aoi22 g1866 (.Z(w1941), .B2(w1759), .A2(w1), .A1(w1811), .B1(w1838) );
	vdp_aoi22 g1867 (.Z(w1942), .B1(1'b0), .A2(w1), .B2(w1759), .A1(w1838) );
	vdp_comp_dff g1868 (.Q(w1645), .D(w1690), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_comp_dff g1869 (.Q(w1792), .D(w1965), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_cnt_bit g1870 (.CI(w1967), .Q(w1853), .nEN(SYSRES), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g1871 (.nZ(w1938), .A(w55) );
	vdp_and g1872 (.Z(w1779), .A(w1794), .B(w1731) );
	vdp_and g1873 (.Z(w1780), .A(w1794), .B(w1731) );
	vdp_and g1874 (.Z(w1782), .A(w1992), .B(w1795) );
	vdp_and g1875 (.Z(w1783), .A(w1795), .B(w1797) );
	vdp_and g1876 (.Z(w1781), .A(w1842), .B(w1747) );
	vdp_and g1877 (.Z(w1992), .A(w1841), .B(w1729) );
	vdp_and g1878 (.Z(w1722), .A(w53), .B(w1709) );
	vdp_and g1879 (.Z(w16), .A(w1959), .B(w1700) );
	vdp_and g1880 (.Z(w1707), .A(w1671), .B(w1709) );
	vdp_and g1881 (.Z(w26), .A(w1630), .B(w1925) );
	vdp_and g1882 (.Z(w1708), .A(w52), .B(w1792) );
	vdp_and g1883 (.Z(w1733), .A(w1923), .B(w53) );
	vdp_and g1884 (.Z(w15), .A(w1700), .B(w1789) );
	vdp_and g1885 (.Z(w1764), .A(w1981), .B(w1733) );
	vdp_and g1886 (.Z(w10), .A(w1852), .B(w1700) );
	vdp_and g1887 (.Z(w1952), .A(w1801), .B(w4) );
	vdp_or g1888 (.Z(w1806), .A(w1927), .B(w1930) );
	vdp_or g1889 (.Z(w1805), .A(w1955), .B(w1930) );
	vdp_and g1890 (.Z(w1766), .A(M5), .B(w23) );
	vdp_and g1891 (.Z(w1967), .A(w1802), .B(w1754) );
	vdp_or g1892 (.Z(w1788), .A(SYSRES), .B(w1787) );
	vdp_or g1893 (.Z(w28), .A(w1773), .B(w1772) );
	vdp_or g1894 (.Z(w24), .A(w1767), .B(w1773) );
	vdp_or g1895 (.Z(w1989), .A(w1779), .B(w1783) );
	vdp_or g1896 (.Z(w1798), .A(w1785), .B(w1744) );
	vdp_or g1897 (.Z(w1926), .A(SYSRES), .B(w1787) );
	vdp_or g1898 (.Z(w1787), .A(w1734), .B(w1799) );
	vdp_or g1899 (.Z(w1964), .A(w1745), .B(SYSRES) );
	vdp_or g1900 (.Z(w1949), .A(w1670), .B(w1991) );
	vdp_or g1901 (.Z(w1993), .A(SYSRES), .B(w1744) );
	vdp_or g1902 (.Z(w1962), .A(w1708), .B(w1645) );
	vdp_or g1903 (.Z(w1911), .A(w1963), .B(w1790) );
	vdp_and g1904 (.Z(w11), .A(w1748), .B(w1700) );
	vdp_and g1905 (.Z(w1790), .A(w1660), .B(w1733) );
	vdp_or g1906 (.Z(w1987), .A(SYSRES), .B(w1734) );
	vdp_not g1907 (.nZ(w1686), .A(w54) );
	vdp_not g1908 (.nZ(w1685), .A(w48) );
	vdp_aon33 g1909 (.Z(w1834), .A3(w1833), .A2(w1938), .A1(w4), .B1(w55), .B3(1'b1), .B2(w1234) );
	vdp_aoi21 g1910 (.Z(w1936), .A1(w1691), .A2(w1700), .B(w1661) );
	vdp_aoi21 g1911 (.Z(w1699), .A1(w1697), .B(w1698), .A2(w1700) );
	vdp_aoi21 g1912 (.Z(w1662), .A1(w40), .A2(w50), .B(w1694) );
	vdp_aoi21 g1913 (.Z(w1725), .A1(w1706), .B(w1960), .A2(w1962) );
	vdp_aoi21 g1914 (.Z(w1957), .A1(w1700), .B(w1956), .A2(w1701) );
	vdp_aoi21 g1915 (.Z(w1756), .B(w1966), .A1(w1700), .A2(w1720) );
	vdp_aoi21 g1916 (.Z(w1937), .A1(w1700), .A2(w1770), .B(w1771) );
	vdp_xor g1917 (.Z(w1754), .B(w1659), .A(w1732) );
	vdp_xor g1918 (.Z(w1803), .A(ODD_EVEN), .B(w1830) );
	vdp_and3 g1919 (.Z(w1661), .A(w1719), .B(w42), .C(w1668) );
	vdp_and3 g1920 (.Z(w1997), .A(w1996), .B(w1857), .C(w1716) );
	vdp_and3 g1921 (.Z(w1698), .A(w1702), .B(w51), .C(w1668) );
	vdp_and3 g1922 (.Z(w1956), .A(w51), .B(w1668), .C(w42) );
	vdp_and3 g1923 (.Z(w1966), .A(w1702), .B(w1719), .C(w1773) );
	vdp_and3 g1924 (.Z(w1771), .A(w42), .B(w1719), .C(w41) );
	vdp_or3 g1925 (.Z(w1988), .A(w1781), .B(w1782), .C(w1780) );
	vdp_and3 g1926 (.Z(w1991), .A(w53), .B(w1709), .C(M5) );
	vdp_and3 g1927 (.Z(w1868), .A(w1706), .B(w53), .C(w1693) );
	vdp_and3 g1928 (.Z(w1670), .A(H40), .B(M5), .C(w1671) );
	vdp_nor4 g1929 (.Z(w1716), .A(w1757), .B(w1793), .C(w1664), .D(w1755) );
	vdp_nor4 g1930 (.Z(w1833), .A(w56), .B(w1836), .D(w1952), .C(SYSRES) );
	vdp_comp_we g1931 (.Z(w1817), .nZ(w1951), .A(w1835) );
	vdp_comp_we g1932 (.Z(w1819), .nZ(w1820), .A(w56) );
	vdp_comp_we g1933 (.Z(w1998), .nZ(w1669), .A(w57) );
	vdp_comp_we g1934 (.Z(w1676), .nZ(w1675), .A(w1660) );
	vdp_and3 g1935 (.Z(w18), .A(w1110), .B(w1925), .C(w31) );
	vdp_or4 g1936 (.Z(w1660), .A(w57), .B(SYSRES), .C(w1868), .D(w1982) );
	vdp_nor3 g1937 (.Z(w1857), .A(w1860), .B(w1717), .C(w1867) );
	vdp_nor3 g1938 (.Z(w1794), .A(w1729), .B(w1842), .C(w1841) );
	vdp_nand g1939 (.Z(w1749), .A(w1750), .B(w1791) );
	vdp_nand g1940 (.Z(w1999), .A(w1713), .B(w1994) );
	vdp_nand g1941 (.Z(w1861), .A(w1958), .B(w1717) );
	vdp_nor3 g1942 (.Z(w1700), .A(w42), .B(w51), .C(w41) );
	vdp_nor g1943 (.Z(w1930), .A(w1830), .B(M5) );
	vdp_nor g1944 (.Z(w1804), .A(ODD_EVEN), .B(w1830) );
	vdp_nor g1945 (.Z(w1927), .A(w1818), .B(PAL) );
	vdp_nor g1946 (.Z(w1955), .A(w1818), .B(w1830) );
	vdp_nor g1947 (.Z(w1960), .A(w1644), .B(SYSRES) );
	vdp_SDELAY8 g1948 (.Q(w1807), .D(w1784), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2), .nC3(nHCLK1), .C3(HCLK1), .nC4(nHCLK2), .C4(HCLK2), .nC5(nHCLK1), .C5(HCLK1), .nC6(nHCLK2), .C6(HCLK2), .nC7(nHCLK1), .C7(HCLK1), .nC8(nHCLK2), .C8(HCLK2), .nC9(nHCLK1), .C9(HCLK1), .nC10(nHCLK2), .C10(HCLK2), .nC11(nHCLK1), .C11(HCLK1), .nC12(nHCLK2), .C12(HCLK2), .nC13(nHCLK1), .C13(HCLK1), .nC14(nHCLK2), .C14(HCLK2), .nC15(nHCLK1), .C15(HCLK1), .nC16(nHCLK2), .C16(HCLK2) );
	vdp_SDELAY7 g1949 (.Q(w1751), .D(w1752), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .nC4(nHCLK2), .C5(HCLK1), .nC5(nHCLK1), .C6(HCLK2), .nC6(nHCLK2), .C7(HCLK1), .nC7(nHCLK1), .C8(HCLK2), .nC8(nHCLK2), .C9(HCLK1), .nC9(nHCLK1), .C10(HCLK2), .nC10(nHCLK2), .C11(HCLK1), .nC11(nHCLK1), .C12(HCLK2), .nC12(nHCLK2), .C13(HCLK1), .nC13(nHCLK1), .C14(HCLK2), .nC14(nHCLK2), .C3(HCLK1) );
	vdp_SDELAY8 g1950 (.Q(w1714), .D(w1754), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2), .C3(HCLK1), .nC4(nHCLK2), .C4(HCLK2), .nC5(nHCLK1), .C5(HCLK1), .nC6(nHCLK2), .C6(HCLK2), .nC7(nHCLK1), .C7(HCLK1), .nC8(nHCLK2), .C8(HCLK2), .nC9(nHCLK1), .C9(HCLK1), .nC10(nHCLK2), .C10(HCLK2), .C11(HCLK1), .nC12(nHCLK2), .C12(HCLK2), .nC13(nHCLK1), .C13(HCLK1), .nC14(nHCLK2), .C14(HCLK2), .nC15(nHCLK1), .C15(HCLK1), .nC16(nHCLK2), .C16(HCLK2), .nC3(nHCLK1), .nC11(nHCLK1) );
	vdp_SDELAY8 g1951 (.Q(w1688), .D(w1659), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2), .C3(HCLK1), .nC4(nHCLK2), .C4(HCLK2), .nC5(nHCLK1), .C5(HCLK1), .nC6(nHCLK2), .C6(HCLK2), .nC7(nHCLK1), .C7(HCLK1), .nC8(nHCLK2), .C8(HCLK2), .nC9(nHCLK1), .C9(HCLK1), .nC10(nHCLK2), .C10(HCLK2), .nC11(nHCLK1), .C11(HCLK1), .nC12(nHCLK2), .C12(HCLK2), .nC13(nHCLK1), .C13(HCLK1), .nC14(nHCLK2), .C14(HCLK2), .nC15(nHCLK1), .C15(HCLK1), .nC16(nHCLK2), .C16(HCLK2), .nC3(nHCLK1) );
	vdp_cnt_bit_load g1952 (.D(w1828), .Q(w1837), .nL(w1951), .L(w1817), .CI(w1922), .nC1(nHCLK1), .CO(w2001), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1953 (.D(w1827), .Q(w1929), .nL(w1951), .L(w1817), .CI(w2001), .nC1(nHCLK1), .CO(w2002), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1954 (.D(w1953), .Q(w1822), .nL(w1951), .L(w1817), .CI(w2002), .nC1(nHCLK1), .CO(w2003), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1955 (.D(w2004), .Q(w1928), .nL(w1951), .L(w1817), .CI(w2003), .nC1(nHCLK1), .CO(w1856), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1956 (.D(w1943), .Q(w1776), .nL(w1951), .L(w1817), .CI(w1856), .nC1(nHCLK1), .CO(w1855), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1957 (.D(w1944), .Q(w1739), .nL(w1951), .L(w1817), .CI(w1855), .nC1(nHCLK1), .CO(w2005), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1958 (.D(w1940), .Q(w1811), .nL(w1951), .L(w1817), .CI(w2005), .nC1(nHCLK1), .CO(w1854), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1959 (.D(w1939), .Q(w1838), .nL(w1951), .L(w1817), .CI(w1854), .nC1(nHCLK1), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1960 (.D(w1809), .Q(w1765), .nL(w1675), .L(w1676), .CI(w1810), .nC1(nHCLK1), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1961 (.D(w1945), .Q(w1737), .nL(w1675), .L(w1676), .CI(w1735), .nC1(nHCLK1), .CO(w1810), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1962 (.D(w1777), .Q(w1907), .nL(w1675), .L(w1676), .CI(w1775), .nC1(nHCLK1), .CO(w1735), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1963 (.D(w1946), .Q(w1760), .nL(w1675), .L(w1676), .CI(w1761), .nC1(nHCLK1), .CO(w1775), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1964 (.D(w1990), .Q(w1728), .nL(w1675), .L(w1676), .CI(w1727), .nC1(nHCLK1), .CO(w1761), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1965 (.D(w1947), .Q(w1683), .nL(w1675), .L(w1676), .CI(w1724), .nC1(nHCLK1), .CO(w1727), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1966 (.D(w1948), .Q(w1684), .nL(w1675), .L(w1676), .CI(w1710), .nC1(nHCLK1), .CO(w1724), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1967 (.D(w1974), .Q(w1679), .nL(w1675), .L(w1676), .CI(w2000), .nC1(nHCLK1), .CO(w1710), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1968 (.D(w1674), .Q(w1932), .nL(w1675), .L(w1676), .CI(w1859), .nC1(nHCLK1), .CO(w2000), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_or8 g1969 (.Z(w1823), .A(w1869), .B(w1870), .C(w1871), .D(w1872), .E(w1919), .F(w1920), .G(w1921), .H(w1874) );
	vdp_or8 g1970 (.Z(w1824), .A(w1875), .B(w1918), .C(w1917), .D(w1900), .E(w1916), .F(w1876), .G(w1877), .H(w1915) );
	vdp_or8 g1971 (.Z(w1825), .A(w2006), .B(w1985), .C(w1986), .D(w1972), .E(w1899), .F(w1898), .G(w1971), .H(w1897) );
	vdp_or5 g1972 (.Z(w1826), .A(w1893), .B(w1894), .C(w1895), .D(w1896), .E(w6780) );
	vdp_or7 g1973 (.Z(w1815), .A(w1889), .B(w1890), .C(w1891), .D(w1892), .E(w6777), .F(w6778), .G(w6779) );
	vdp_or7 g1974 (.Z(w1813), .A(w1878), .B(w1879), .C(w1880), .D(w1881), .E(w1882), .F(w1883), .G(w1884) );
	vdp_nor g1975 (.Z(w1694), .A(w1660), .B(w40) );
	vdp_and g1976 (.Z(w17), .A(w1700), .B(w1718) );
	vdp_not g1977 (.nZ(w1643), .A(w1885) );
	vdp_nor3 g1978 (.Z(w1814), .A(w1888), .B(w1887), .C(w1886) );
	vdp_rs_ff g1979 (.S(w1924), .R(w1626), .Q(w1624) );
	vdp_rs_ff g1980 (.S(w1638), .R(w1634), .Q(w1622) );
	vdp_and g1981 (.Z(w1841), .A(w1613), .B(M5) );
	vdp_nor4 g1982 (.Z(w1996), .A(w1682), .B(w1681), .C(w1680), .D(w1678) );
	vdp_nand3 g1983 (.A(w2127), .B(w2126), .C(w2124), .Z(w2120) );
	vdp_nand3 g1984 (.A(w2124), .B(w2126), .C(w2129), .Z(w2115) );
	vdp_nand3 g1985 (.A(w2124), .B(w2127), .C(w2128), .Z(w2116) );
	vdp_nand3 g1986 (.A(w2128), .B(w2124), .C(w2129), .Z(w2117) );
	vdp_nand3 g1987 (.A(w2128), .B(w2125), .C(w2129), .Z(w2112) );
	vdp_nand3 g1988 (.A(w2125), .B(w2127), .C(w2128), .Z(w2111) );
	vdp_nand3 g1989 (.A(w2126), .B(w2125), .C(w2129), .Z(w2119) );
	vdp_nand3 g1990 (.A(w2127), .B(w2126), .C(w2125), .Z(w2118) );
	vdp_nand3 g1991 (.A(w2100), .B(w2101), .C(w2096), .Z(w2110) );
	vdp_nand3 g1992 (.A(w2096), .B(w2101), .C(w2099), .Z(w2109) );
	vdp_nand3 g1993 (.A(w2098), .B(w2097), .C(w2099), .Z(w2103) );
	vdp_nand3 g1994 (.A(w2097), .B(w2100), .C(w2098), .Z(w2104) );
	vdp_nand3 g1995 (.A(w2101), .B(w2097), .C(w2099), .Z(w2105) );
	vdp_nand3 g1996 (.A(w2100), .B(w2101), .C(w2097), .Z(w2106) );
	vdp_nand3 g1997 (.A(w2098), .B(w2096), .C(w2099), .Z(w2107) );
	vdp_nand3 g1998 (.A(w2096), .B(w2100), .C(w2098), .Z(w2108) );
	vdp_nand3 g1999 (.A(w2088), .B(w2086), .C(w2084), .Z(w2081) );
	vdp_nand3 g2000 (.A(w2084), .B(w2086), .C(w2089), .Z(w2080) );
	vdp_nand3 g2001 (.A(w2087), .B(w2085), .C(w2089), .Z(w2074) );
	vdp_nand3 g2002 (.A(w2085), .B(w2088), .C(w2087), .Z(w2075) );
	vdp_nand3 g2003 (.A(w2086), .B(w2085), .C(w2089), .Z(w2076) );
	vdp_nand3 g2004 (.A(w2088), .B(w2086), .C(w2085), .Z(w2077) );
	vdp_nand3 g2005 (.A(w2087), .B(w2084), .C(w2089), .Z(w2078) );
	vdp_nand3 g2006 (.A(w2084), .B(w2088), .C(w2087), .Z(w2079) );
	vdp_nand3 g2007 (.A(w2027), .B(w2024), .C(w2028), .Z(w2021) );
	vdp_nand3 g2008 (.A(w2028), .B(w2024), .C(w2026), .Z(w2020) );
	vdp_nand3 g2009 (.A(w2025), .B(w2023), .C(w2026), .Z(w2014) );
	vdp_nand3 g2010 (.A(w2023), .B(w2027), .C(w2025), .Z(w2015) );
	vdp_nand3 g2011 (.A(w2024), .B(w2023), .C(w2026), .Z(w2016) );
	vdp_nand3 g2012 (.A(w2027), .B(w2024), .C(w2023), .Z(w2017) );
	vdp_nand3 g2013 (.A(w2025), .B(w2028), .C(w2026), .Z(w2018) );
	vdp_nand3 g2014 (.A(w2028), .B(w2027), .C(w2025), .Z(w2019) );
	vdp_not g2015 (.nZ(w2022), .A(w2009) );
	vdp_not g2016 (.nZ(w2082), .A(w2010) );
	vdp_not g2017 (.nZ(w2090), .A(w2007) );
	vdp_not g2018 (.nZ(w2121), .A(w2008) );
	vdp_nand g2019 (.Z(w2012), .B(w2013), .A(w2022) );
	vdp_nand g2020 (.Z(w2013), .B(w2022), .A(w2029) );
	vdp_nand g2021 (.Z(w2072), .B(w2073), .A(w2082) );
	vdp_nand g2022 (.Z(w2073), .B(w2082), .A(w2033) );
	vdp_comp_we g2023 (.A(w2083), .Z(w2085), .nZ(w2084) );
	vdp_comp_we g2024 (.A(w2143), .Z(w2087), .nZ(w2086) );
	vdp_comp_we g2025 (.A(w2142), .Z(w2089), .nZ(w2088) );
	vdp_comp_we g2026 (.A(w2030), .Z(w2023), .nZ(w2028) );
	vdp_comp_we g2027 (.A(w2031), .Z(w2025), .nZ(w2024) );
	vdp_comp_we g2028 (.A(w2032), .Z(w2026), .nZ(w2027) );
	vdp_nand g2029 (.Z(w2091), .B(w2090), .A(w2094) );
	vdp_comp_we g2030 (.A(w2093), .Z(w2097), .nZ(w2096) );
	vdp_comp_we g2031 (.A(w2095), .Z(w2098), .nZ(w2101) );
	vdp_comp_we g2032 (.A(w2102), .Z(w2099), .nZ(w2100) );
	vdp_nand g2033 (.Z(w2092), .B(w2091), .A(w2090) );
	vdp_nand g2034 (.Z(w2113), .B(w2121), .A(w2122) );
	vdp_comp_we g2035 (.A(w2123), .Z(w2125), .nZ(w2124) );
	vdp_comp_we g2036 (.A(w2130), .Z(w2128), .nZ(w2126) );
	vdp_comp_we g2037 (.A(w2131), .Z(w2129), .nZ(w2127) );
	vdp_nand g2038 (.Z(w2114), .B(w2113), .A(w2121) );
	vdp_comp_str g2039 (.A(w2154), .Z(w2155), .nZ(w2153) );
	vdp_comp_str g2040 (.A(w2171), .Z(w2144), .nZ(w2145) );
	vdp_comp_str g2041 (.A(w2180), .Z(w2135), .nZ(w2134) );
	vdp_comp_str g2042 (.A(w2181), .Z(w2036), .nZ(w2035) );
	vdp_comp_str g2043 (.A(w2044), .Z(w2045), .nZ(w2046) );
	vdp_comp_str g2044 (.A(w2218), .Z(w2404), .nZ(w2281) );
	vdp_comp_str g2045 (.A(w2430), .Z(w2397), .nZ(w2396) );
	vdp_comp_str g2046 (.A(w2400), .Z(w2411), .nZ(w2398) );
	vdp_comp_str g2047 (.A(w2189), .Z(w2401), .nZ(w2399) );
	vdp_comp_str g2048 (.A(w2309), .Z(w2052), .nZ(w2056) );
	vdp_comp_str g2049 (.A(w2431), .Z(w2053), .nZ(w2057) );
	vdp_comp_str g2050 (.A(w2187), .Z(w2055), .nZ(w2058) );
	vdp_slatch g2051 (.Q(w2415), .C(w2055), .D(w2182), .nC(w2058) );
	vdp_slatch g2052 (.Q(w2414), .C(w2053), .D(w2182), .nC(w2057) );
	vdp_slatch g2053 (.Q(w2376), .C(w2055), .D(w2316), .nC(w2058) );
	vdp_slatch g2054 (.Q(w2413), .C(w2052), .D(w2182), .nC(w2056) );
	vdp_slatch g2055 (.Q(w2418), .C(w2055), .D(w2317), .nC(w2058) );
	vdp_slatch g2056 (.Q(w2375), .C(w2052), .D(w2316), .nC(w2056) );
	vdp_slatch g2057 (.Q(w2377), .C(w2053), .D(w2316), .nC(w2057) );
	vdp_slatch g2058 (.Q(w2311), .C(w2055), .D(w2319), .nC(w2058) );
	vdp_slatch g2059 (.Q(w2416), .C(w2052), .D(w2317), .nC(w2056) );
	vdp_slatch g2060 (.Q(w2417), .C(w2053), .D(w2317), .nC(w2057) );
	vdp_slatch g2061 (.Q(w2065), .C(w2055), .D(w2054), .nC(w2058) );
	vdp_slatch g2062 (.Q(w2310), .C(w2052), .D(w2319), .nC(w2056) );
	vdp_slatch g2063 (.Q(w2312), .C(w2053), .D(w2319), .nC(w2057) );
	vdp_slatch g2064 (.Q(w2062), .C(w2052), .D(w2054), .nC(w2056) );
	vdp_slatch g2065 (.Q(w2064), .C(w2053), .D(w2054), .nC(w2057) );
	vdp_slatch g2066 (.Q(w2059), .C(w2055), .D(w2051), .nC(w2058) );
	vdp_slatch g2067 (.Q(w2071), .C(w2052), .D(w2051), .nC(w2056) );
	vdp_slatch g2068 (.Q(w2060), .C(w2053), .D(w2051), .nC(w2057) );
	vdp_slatch g2069 (.Q(w2390), .C(w2401), .D(w2182), .nC(w2399) );
	vdp_slatch g2070 (.Q(w2389), .C(w2411), .D(w2182), .nC(w2398) );
	vdp_slatch g2071 (.Q(w2395), .C(w2401), .D(w2316), .nC(w2399) );
	vdp_slatch g2072 (.Q(w2391), .C(w2397), .D(w2182), .nC(w2396) );
	vdp_slatch g2073 (.Q(w2383), .C(w2401), .D(w2409), .nC(w2399) );
	vdp_slatch g2074 (.Q(w2393), .C(w2397), .D(w2316), .nC(w2396) );
	vdp_slatch g2075 (.Q(w2394), .C(w2411), .D(w2316), .nC(w2398) );
	vdp_slatch g2076 (.Q(w2380), .C(w2401), .D(w2319), .nC(w2399) );
	vdp_slatch g2077 (.Q(w2381), .C(w2397), .D(w2409), .nC(w2396) );
	vdp_slatch g2078 (.Q(w2382), .C(w2411), .D(w2409), .nC(w2398) );
	vdp_slatch g2079 (.Q(w2378), .C(w2397), .D(w2319), .nC(w2396) );
	vdp_slatch g2080 (.Q(w2379), .C(w2411), .D(w2319), .nC(w2398) );
	vdp_slatch g2081 (.Q(w2265), .C(w2404), .D(w2409), .nC(w2281) );
	vdp_slatch g2082 (.Q(w2407), .C(w2404), .D(w2316), .nC(w2281) );
	vdp_slatch g2083 (.Q(w2408), .C(w2404), .D(w2182), .nC(w2281) );
	vdp_and g2084 (.Z(w2225), .A(w2408), .B(w2407) );
	vdp_and g2085 (.Z(w2392), .A(w2407), .B(w2405) );
	vdp_and g2086 (.Z(w2374), .A(w2408), .B(w2406) );
	vdp_and g2087 (.Z(w2320), .A(w2405), .B(w2406) );
	vdp_slatch g2088 (.Q(w2157), .C(w2155), .D(w2151), .nC(w2153) );
	vdp_or g2089 (.Z(w2131), .A(w2156), .B(w2157) );
	vdp_notif0 g2090 (.A(w2131), .nZ(DB[0]), .nE(w2037) );
	vdp_slatch g2091 (.Q(w2441), .C(w2155), .D(w2148), .nC(w2153) );
	vdp_or g2092 (.Z(w2130), .A(w2156), .B(w2441) );
	vdp_notif0 g2093 (.A(w2130), .nZ(DB[1]), .nE(w2037) );
	vdp_slatch g2094 (.Q(w2442), .C(w2155), .D(w2150), .nC(w2153) );
	vdp_or g2095 (.Z(w2123), .A(w2156), .B(w2442) );
	vdp_notif0 g2096 (.A(w2123), .nZ(DB[2]), .nE(w2037) );
	vdp_slatch g2097 (.Q(w2161), .C(w2155), .D(w2162), .nC(w2153) );
	vdp_or g2098 (.Z(w2122), .A(w2156), .B(w2161) );
	vdp_notif0 g2099 (.A(w2122), .nZ(DB[3]), .nE(w2037) );
	vdp_slatch g2100 (.Q(w2152), .C(w2144), .D(w2151), .nC(w2145) );
	vdp_or g2101 (.Z(w2102), .A(w2149), .B(w2152) );
	vdp_notif0 g2102 (.A(w2102), .nZ(DB[4]), .nE(w2037) );
	vdp_slatch g2103 (.Q(w2147), .C(w2144), .D(w2148), .nC(w2145) );
	vdp_or g2104 (.Z(w2095), .A(w2149), .B(w2147) );
	vdp_notif0 g2105 (.A(w2095), .nZ(DB[5]), .nE(w2037) );
	vdp_slatch g2106 (.Q(w2146), .C(w2144), .D(w2150), .nC(w2145) );
	vdp_or g2107 (.Z(w2093), .A(w2149), .B(w2146) );
	vdp_notif0 g2108 (.A(w2093), .nZ(DB[6]), .nE(w2037) );
	vdp_slatch g2109 (.Q(w2141), .C(w2144), .D(w2162), .nC(w2145) );
	vdp_or g2110 (.Z(w2094), .A(w2149), .B(w2141) );
	vdp_notif0 g2111 (.A(w2094), .nZ(DB[7]), .nE(w2037) );
	vdp_slatch g2112 (.Q(w2440), .C(w2135), .D(w2151), .nC(w2134) );
	vdp_or g2113 (.Z(w2142), .A(w2136), .B(w2440) );
	vdp_notif0 g2114 (.A(w2142), .nZ(DB[8]), .nE(w2037) );
	vdp_slatch g2115 (.Q(w2140), .C(w2135), .D(w2148), .nC(w2134) );
	vdp_or g2116 (.Z(w2143), .A(w2136), .B(w2140) );
	vdp_notif0 g2117 (.A(w2143), .nZ(DB[9]), .nE(w2037) );
	vdp_slatch g2118 (.Q(w2133), .C(w2135), .D(w2150), .nC(w2134) );
	vdp_or g2119 (.Z(w2083), .A(w2136), .B(w2133) );
	vdp_notif0 g2120 (.A(w2083), .nZ(DB[10]), .nE(w2037) );
	vdp_slatch g2121 (.Q(w2132), .C(w2135), .D(w2162), .nC(w2134) );
	vdp_or g2122 (.Z(w2033), .A(w2136), .B(w2132) );
	vdp_notif0 g2123 (.A(w2033), .nZ(DB[11]), .nE(w2037) );
	vdp_slatch g2124 (.Q(w2038), .C(w2036), .D(w2151), .nC(w2035) );
	vdp_or g2125 (.Z(w2032), .A(w2034), .B(w2038) );
	vdp_notif0 g2126 (.A(w2032), .nZ(DB[12]), .nE(w2037) );
	vdp_slatch g2127 (.Q(w2039), .C(w2036), .D(w2148), .nC(w2035) );
	vdp_or g2128 (.Z(w2031), .A(w2034), .B(w2039) );
	vdp_notif0 g2129 (.A(w2031), .nZ(DB[13]), .nE(w2037) );
	vdp_slatch g2130 (.Q(w2040), .C(w2036), .D(w2150), .nC(w2035) );
	vdp_or g2131 (.Z(w2030), .A(w2034), .B(w2040) );
	vdp_notif0 g2132 (.A(w2030), .nZ(DB[14]), .nE(w2037) );
	vdp_slatch g2133 (.Q(w2041), .C(w2036), .D(w2162), .nC(w2035) );
	vdp_or g2134 (.Z(w2029), .A(w2034), .B(w2041) );
	vdp_notif0 g2135 (.A(w2029), .nZ(DB[15]), .nE(w2037) );
	vdp_not g2136 (.A(PSG_TEST_OE), .nZ(w2037) );
	vdp_not g2137 (.nZ(w2210), .A(PSG_Z80_CLK) );
	vdp_clkgen g2138 (.PH(w2210), .CLK1(w2211), .nCLK1(w2212), .CLK2(w2213), .nCLK2(w2214) );
	vdp_comp_dff g2139 (.D(SYSRES), .nC1(w2212), .C1(w2211), .C2(w2213), .nC2(w2214), .Q(w2242) );
	vdp_sr_bit g2140 (.D(w2242), .nC1(w2212), .nC2(w2214), .C1(w2211), .C2(w2213), .Q(w2244) );
	vdp_sr_bit g2141 (.D(w2217), .nC1(w2212), .nC2(w2214), .C1(w2211), .C2(w2213), .Q(w2216) );
	vdp_not g2142 (.nZ(w2243), .A(w2244) );
	vdp_and g2143 (.Z(w2215), .A(w2242), .B(w2243) );
	vdp_nor g2144 (.Z(w2217), .A(w2216), .B(w2215) );
	vdp_cnt_bit g2145 (.CI(w2216), .R(w2215), .C1(w2211), .nC1(w2212), .nC2(w2214), .C2(w2213), .Q(w2241) );
	vdp_dlatch_inv g2146 (.nQ(w2240), .D(w2241), .nC(w2212), .C(w2211) );
	vdp_not g2147 (.nZ(w2239), .A(w2240) );
	vdp_nand g2148 (.Z(w2238), .A(w2216), .B(w2240) );
	vdp_not g2149 (.nZ(w2237), .A(w2238) );
	vdp_not g2150 (.nZ(w2236), .A(w2235) );
	vdp_not g2151 (.nZ(PSG_CLK1), .A(w2238) );
	vdp_not g2152 (.nZ(PSG_nCLK1), .A(w2237) );
	vdp_not g2153 (.nZ(PSG_nCLK2), .A(w2236) );
	vdp_not g2154 (.nZ(PSG_CLK2), .A(w2235) );
	vdp_nand g2155 (.Z(w2235), .A(w2216), .B(w2239) );
	vdp_sr_bit g2156 (.D(w2345), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2201) );
	vdp_sr_bit g2157 (.D(w2346), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2345) );
	vdp_sr_bit g2158 (.D(w2344), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2346) );
	vdp_sr_bit g2159 (.D(w2205), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2344) );
	vdp_sr_bit g2160 (.D(w2343), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2204) );
	vdp_sr_bit g2161 (.D(w2342), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2343) );
	vdp_sr_bit g2162 (.D(w2341), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2342) );
	vdp_sr_bit g2163 (.D(w2209), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2341) );
	vdp_sr_bit g2164 (.D(w2340), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2208) );
	vdp_sr_bit g2165 (.D(w2339), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2340) );
	vdp_sr_bit g2166 (.D(w2338), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2339) );
	vdp_sr_bit g2167 (.D(w2271), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2338) );
	vdp_sr_bit g2168 (.D(w2336), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2270) );
	vdp_sr_bit g2169 (.D(w2337), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2336) );
	vdp_sr_bit g2170 (.D(w2335), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2337) );
	vdp_sr_bit g2171 (.D(w2269), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2335) );
	vdp_sr_bit g2172 (.D(w2334), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2268) );
	vdp_sr_bit g2173 (.D(w2333), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2334) );
	vdp_sr_bit g2174 (.D(w2332), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2333) );
	vdp_sr_bit g2175 (.D(w2257), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2332) );
	vdp_sr_bit g2176 (.D(w2331), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2256) );
	vdp_sr_bit g2177 (.D(w2330), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2331) );
	vdp_sr_bit g2178 (.D(w2327), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2330) );
	vdp_sr_bit g2179 (.D(w2254), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2327) );
	vdp_sr_bit g2180 (.D(w2328), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2255) );
	vdp_sr_bit g2181 (.D(w2329), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2328) );
	vdp_sr_bit g2182 (.D(w2355), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2329) );
	vdp_sr_bit g2183 (.D(w2323), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2355) );
	vdp_sr_bit g2184 (.D(w2354), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2324) );
	vdp_sr_bit g2185 (.D(w2356), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2354) );
	vdp_sr_bit g2186 (.D(w2357), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2356) );
	vdp_sr_bit g2187 (.D(w2292), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2357) );
	vdp_sr_bit g2188 (.D(w2282), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2291) );
	vdp_sr_bit g2189 (.D(w2283), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2282) );
	vdp_sr_bit g2190 (.D(w2284), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2283) );
	vdp_sr_bit g2191 (.D(w2293), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2284) );
	vdp_sr_bit g2192 (.D(w2199), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2289) );
	vdp_sr_bit g2193 (.D(w2198), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2199) );
	vdp_sr_bit g2194 (.D(w2197), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2198) );
	vdp_sr_bit g2195 (.D(w2195), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2197) );
	vdp_aon2222 g2196 (.Z(w2067), .D2(1'b0), .C2(w2071), .C1(w2063), .D1(w2070), .B1(w2060), .A2(w2059), .A1(w2061), .B2(w2069) );
	vdp_cgi2a g2197 (.Z(w2410), .A(w2067), .C(w2422), .B(w2201) );
	vdp_aon2222 g2198 (.Z(w2068), .D2(1'b0), .C2(w2062), .C1(w2063), .D1(w2070), .B1(w2064), .A2(w2065), .A1(w2061), .B2(w2069) );
	vdp_cgi2a g2199 (.Z(w2422), .A(w2068), .C(w2421), .B(w2204) );
	vdp_aon2222 g2200 (.Z(w2315), .D2(1'b0), .C2(w2310), .C1(w2063), .D1(w2070), .B1(w2312), .A2(w2311), .A1(w2061), .B2(w2069) );
	vdp_cgi2a g2201 (.Z(w2421), .A(w2315), .C(w2420), .B(w2208) );
	vdp_aon2222 g2202 (.Z(w2314), .D2(w2392), .C2(w2416), .C1(w2063), .D1(w2070), .B1(w2417), .A2(w2418), .A1(w2061), .B2(w2069) );
	vdp_cgi2a g2203 (.Z(w2420), .A(w2314), .C(w2321), .B(w2270) );
	vdp_aon2222 g2204 (.Z(w2313), .D2(w2374), .C2(w2375), .C1(w2063), .D1(w2070), .B1(w2377), .A2(w2376), .A1(w2061), .B2(w2069) );
	vdp_cgi2a g2205 (.Z(w2321), .A(w2313), .C(w2322), .B(w2268) );
	vdp_aon2222 g2206 (.Z(w2385), .D2(w2320), .C2(w2413), .C1(w2063), .D1(w2070), .B1(w2414), .A2(w2415), .A1(w2061), .B2(w2069) );
	vdp_cgi2a g2207 (.Z(w2322), .A(w2385), .C(w2419), .B(w2256) );
	vdp_aon2222 g2208 (.Z(w2384), .D2(1'b0), .C2(w2378), .C1(w2063), .D1(w2070), .B1(w2379), .A2(w2380), .A1(w2061), .B2(w2069) );
	vdp_cgi2a g2209 (.Z(w2419), .A(w2384), .C(w2412), .B(w2255) );
	vdp_aon2222 g2210 (.Z(w2386), .D2(1'b0), .C2(w2381), .C1(w2063), .D1(w2070), .B1(w2382), .A2(w2383), .A1(w2061), .B2(w2069) );
	vdp_cgi2a g2211 (.Z(w2412), .A(w2386), .C(w2285), .B(w2324) );
	vdp_aon2222 g2212 (.Z(w2387), .D2(1'b0), .C2(w2393), .C1(w2063), .D1(w2070), .B1(w2394), .A2(w2395), .A1(w2061), .B2(w2069) );
	vdp_cgi2a g2213 (.Z(w2285), .A(w2387), .C(w2286), .B(w2291) );
	vdp_aon2222 g2214 (.Z(w2288), .D2(1'b0), .C2(w2391), .C1(w2063), .D1(w2070), .B1(w2389), .A2(w2390), .A1(w2061), .B2(w2069) );
	vdp_cgi2a g2215 (.Z(w2286), .A(w2288), .C(1'b1), .B(w2289) );
	vdp_not g2216 (.nZ(w2070), .A(w2388) );
	vdp_sr_bit g2217 (.D(w2369), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .Q(w2290) );
	vdp_nand g2218 (.Z(w2388), .A(w2364), .B(w2290) );
	vdp_not g2219 (.nZ(w2063), .A(w2370) );
	vdp_sr_bit g2220 (.D(w2365), .Q(w2369), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_nand g2221 (.Z(w2370), .A(w2364), .B(w2369) );
	vdp_not g2222 (.nZ(w2069), .A(w2368) );
	vdp_sr_bit g2223 (.D(w2301), .Q(w2365), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_nand g2224 (.Z(w2368), .A(w2364), .B(w2365) );
	vdp_not g2225 (.nZ(w2061), .A(w2366) );
	vdp_sr_bit g2226 (.D(w2367), .Q(w2301), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_nand g2227 (.Z(w2366), .A(w2364), .B(w2301) );
	vdp_sr_bit g2228 (.D(w2191), .Q(w2272), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_sr_bit g2229 (.D(w2373), .Q(w2371), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_sr_bit g2230 (.D(w2372), .Q(w2373), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_sr_bit g2231 (.D(w2300), .Q(w2372), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_sr_bit g2232 (.D(w2410), .Q(w2300), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_not g2233 (.nZ(w2364), .A(w2272) );
	vdp_nor4 g2234 (.Z(w2367), .A(w2369), .B(w2365), .D(w2301), .C(w2191) );
	vdp_nor4 g2235 (.Z(w2262), .A(w2304), .B(w2305), .D(w2302), .C(w2303) );
	vdp_nor4 g2236 (.Z(w2264), .A(w2297), .B(w2298), .D(w2277), .C(w2278) );
	vdp_nor3 g2237 (.Z(w2263), .A(w2273), .B(w2274), .C(w2275) );
	vdp_not g2238 (.nZ(w2049), .A(w2272) );
	vdp_nand4 g2239 (.Z(w2261), .A(w2262), .B(w2264), .D(w2232), .C(w2263) );
	vdp_nand g2240 (.Z(w2266), .A(w2200), .B(w2265) );
	vdp_nand g2241 (.Z(w2267), .A(w2261), .B(w2266) );
	vdp_lfsr_bit g2242 (.Q(w2297), .A(w2267), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2295), .B(w2296) );
	vdp_lfsr_bit g2243 (.Q(w2298), .A(w2297), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2295), .B(w2296) );
	vdp_lfsr_bit g2244 (.Q(w2278), .A(w2298), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2295), .B(w2296) );
	vdp_lfsr_bit g2245 (.Q(w2277), .A(w2278), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2295), .B(w2296) );
	vdp_lfsr_bit g2246 (.Q(w2273), .A(w2277), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2295), .B(w2296) );
	vdp_lfsr_bit g2247 (.Q(w2274), .A(w2273), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2295), .B(w2296) );
	vdp_lfsr_bit g2248 (.Q(w2275), .A(w2274), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2295), .B(w2296) );
	vdp_lfsr_bit g2249 (.Q(w2302), .A(w2275), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2295), .B(w2296) );
	vdp_lfsr_bit g2250 (.Q(w2303), .A(w2302), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2295), .B(w2296) );
	vdp_lfsr_bit g2251 (.Q(w2304), .A(w2303), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2295), .B(w2296) );
	vdp_lfsr_bit g2252 (.Q(w2305), .A(w2304), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2295), .B(w2296) );
	vdp_lfsr_bit g2253 (.Q(w2306), .A(w2305), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2295), .B(w2296) );
	vdp_lfsr_bit g2254 (.Q(w2307), .A(w2306), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2295), .B(w2296) );
	vdp_lfsr_bit g2255 (.Q(w2294), .A(w2307), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2295), .B(w2296) );
	vdp_lfsr_bit g2256 (.Q(w2194), .A(w2294), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2295), .B(w2296) );
	vdp_lfsr_bit g2257 (.Q(w2308), .A(w2194), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2295), .B(w2296) );
	vdp_xor g2258 (.Z(w2200), .A(w2307), .B(w2308) );
	vdp_and g2259 (.Z(w2353), .A(w2196), .B(w2289) );
	vdp_ha g2260 (.SUM(w2195), .CO(w2251), .B(w2353), .A(1'b1) );
	vdp_and g2261 (.Z(w2326), .A(w2196), .B(w2291) );
	vdp_ha g2262 (.SUM(w2293), .CO(w2250), .B(w2326), .A(w2251) );
	vdp_and g2263 (.Z(w2325), .A(w2196), .B(w2324) );
	vdp_ha g2264 (.SUM(w2292), .CO(w2249), .B(w2325), .A(w2250) );
	vdp_and g2265 (.Z(w2253), .A(w2196), .B(w2255) );
	vdp_ha g2266 (.SUM(w2323), .CO(w2248), .B(w2253), .A(w2249) );
	vdp_and g2267 (.Z(w2352), .A(w2196), .B(w2256) );
	vdp_ha g2268 (.SUM(w2254), .CO(w2247), .B(w2352), .A(w2248) );
	vdp_and g2269 (.Z(w2351), .A(w2196), .B(w2268) );
	vdp_ha g2270 (.SUM(w2257), .CO(w2246), .B(w2351), .A(w2247) );
	vdp_and g2271 (.Z(w2350), .A(w2196), .B(w2270) );
	vdp_ha g2272 (.SUM(w2269), .CO(w2245), .B(w2350), .A(w2246) );
	vdp_and g2273 (.Z(w2349), .A(w2196), .B(w2208) );
	vdp_ha g2274 (.SUM(w2271), .CO(w2207), .B(w2349), .A(w2245) );
	vdp_and g2275 (.Z(w2348), .A(w2196), .B(w2204) );
	vdp_ha g2276 (.SUM(w2209), .CO(w2206), .B(w2348), .A(w2207) );
	vdp_and g2277 (.Z(w2347), .A(w2196), .B(w2201) );
	vdp_ha g2278 (.SUM(w2205), .B(w2347), .A(w2206) );
	vdp_and g2279 (.Z(w2276), .A(w2301), .B(w2371) );
	vdp_cnt_bit g2280 (.CI(w2276), .R(w2272), .C1(PSG_CLK1), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C2(PSG_CLK2), .Q(w2402) );
	vdp_and g2281 (.Z(w2280), .A(w2301), .B(w2373) );
	vdp_cnt_bit g2282 (.CI(w2280), .R(w2272), .C1(PSG_CLK1), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C2(PSG_CLK2), .Q(w2403) );
	vdp_and g2283 (.Z(w2279), .A(w2301), .B(w2372) );
	vdp_cnt_bit g2284 (.CI(w2279), .R(w2272), .C1(PSG_CLK1), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C2(PSG_CLK2), .Q(w2226) );
	vdp_and g2285 (.Z(w2299), .A(w2301), .B(w2300) );
	vdp_cnt_bit g2286 (.CI(w2299), .R(w2272), .C1(PSG_CLK1), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C2(PSG_CLK2), .Q(w2219) );
	vdp_nor g2287 (.Z(w2196), .A(w2410), .B(w2272) );
	vdp_slatch g2288 (.Q(w2050), .C(w2047), .D(DB[7]), .nC(w2048) );
	vdp_comp_str g2289 (.A(w1060), .Z(w2047), .nZ(w2048) );
	vdp_and g2290 (.Z(w2042), .A(w2049), .B(w2050) );
	vdp_and g2291 (.Z(w2044), .A(w2043), .B(w2042) );
	vdp_and g2292 (.Z(w2429), .A(w2049), .B(w2428) );
	vdp_slatch g2293 (.Q(w2428), .C(w2047), .D(DB[6]), .nC(w2048) );
	vdp_slatch g2294 (.Q(w2170), .C(w2045), .D(w2429), .nC(w2046) );
	vdp_and g2295 (.Z(w2051), .A(w2049), .B(w2138) );
	vdp_slatch g2296 (.Q(w2138), .C(w2047), .D(DB[5]), .nC(w2048) );
	vdp_slatch g2297 (.Q(w2139), .C(w2045), .D(w2051), .nC(w2046) );
	vdp_and g2298 (.Z(w2054), .A(w2049), .B(w2137) );
	vdp_slatch g2299 (.Q(w2137), .C(w2047), .D(DB[4]), .nC(w2048) );
	vdp_slatch g2300 (.Q(w2169), .C(w2045), .D(w2054), .nC(w2046) );
	vdp_and g2301 (.Z(w2319), .A(w2049), .B(w2176) );
	vdp_slatch g2302 (.Q(w2176), .C(w2047), .D(DB[3]), .nC(w2048) );
	vdp_or g2303 (.Z(w2162), .A(w2177), .B(w2319) );
	vdp_and g2304 (.Z(w2317), .A(w2049), .B(w2427) );
	vdp_or g2305 (.Z(w2150), .A(w2177), .B(w2317) );
	vdp_slatch g2306 (.Q(w2427), .C(w2047), .D(DB[2]), .nC(w2048) );
	vdp_not g2307 (.nZ(w2177), .A(w2049) );
	vdp_and g2308 (.Z(w2316), .A(w2049), .B(w2318) );
	vdp_or g2309 (.Z(w2148), .A(w2177), .B(w2316) );
	vdp_slatch g2310 (.Q(w2318), .C(w2047), .D(DB[1]), .nC(w2048) );
	vdp_and g2311 (.Z(w2182), .A(w2049), .B(w2183) );
	vdp_or g2312 (.Z(w2151), .A(w2177), .B(w2182) );
	vdp_slatch g2313 (.Q(w2183), .C(w2047), .D(DB[0]), .nC(w2048) );
	vdp_not g2314 (.nZ(w2181), .A(w2179) );
	vdp_aoi21 g2315 (.Z(w2179), .B(w2191), .A1(w2184), .A2(w2178) );
	vdp_and3 g2316 (.Z(w2178), .A(w2159), .B(w2158), .C(w2169) );
	vdp_not g2317 (.nZ(w2180), .A(w2425) );
	vdp_aoi21 g2318 (.Z(w2425), .B(w2191), .A1(w2184), .A2(w2426) );
	vdp_and3 g2319 (.Z(w2426), .A(w2159), .B(w2139), .C(w2169) );
	vdp_not g2320 (.nZ(w2443), .A(w2424) );
	vdp_aoi21 g2321 (.Z(w2424), .B(w2191), .A1(w2184), .A2(w2423) );
	vdp_and3 g2322 (.Z(w2423), .A(w2170), .B(w2158), .C(w2160) );
	vdp_not g2323 (.nZ(w2188), .A(w2042) );
	vdp_or g2324 (.Z(w2190), .A(w2042), .B(w2191) );
	vdp_and g2325 (.Z(w2430), .A(w2190), .B(w2443) );
	vdp_and g2326 (.Z(w2309), .A(w2188), .B(w2443) );
	vdp_and g2327 (.Z(w2400), .A(w2190), .B(w2175) );
	vdp_and g2328 (.Z(w2431), .A(w2188), .B(w2175) );
	vdp_not g2329 (.nZ(w2175), .A(w2174) );
	vdp_aoi21 g2330 (.Z(w2174), .B(w2191), .A1(w2184), .A2(w2173) );
	vdp_and3 g2331 (.Z(w2173), .A(w2159), .B(w2139), .C(w2160) );
	vdp_not g2332 (.nZ(w2171), .A(w2172) );
	vdp_aoi21 g2333 (.Z(w2172), .B(w2191), .A1(w2184), .A2(w2186) );
	vdp_and3 g2334 (.Z(w2186), .A(w2170), .B(w2158), .C(w2169) );
	vdp_and g2335 (.Z(w2189), .A(w2190), .B(w2185) );
	vdp_and g2336 (.Z(w2187), .A(w2188), .B(w2185) );
	vdp_not g2337 (.nZ(w2185), .A(w2168) );
	vdp_aoi21 g2338 (.Z(w2168), .B(w2191), .A1(w2184), .A2(w2167) );
	vdp_and3 g2339 (.Z(w2167), .A(w2159), .B(w2158), .C(w2160) );
	vdp_and3 g2340 (.Z(w2166), .A(w2170), .B(w2139), .C(w2169) );
	vdp_not g2341 (.nZ(w2154), .A(w2165) );
	vdp_aoi21 g2342 (.Z(w2165), .B(w2191), .A1(w2184), .A2(w2166) );
	vdp_and3 g2343 (.Z(w2163), .A(w2170), .B(w2139), .C(w2160) );
	vdp_not g2344 (.nZ(w2218), .A(w2164) );
	vdp_aoi21 g2345 (.Z(w2164), .B(w2191), .A1(w2184), .A2(w2163) );
	vdp_not g2346 (.nZ(w2405), .A(w2408) );
	vdp_not g2347 (.nZ(w2406), .A(w2407) );
	vdp_not g2348 (.nZ(w2160), .A(w2169) );
	vdp_not g2349 (.nZ(w2158), .A(w2139) );
	vdp_not g2350 (.nZ(w2159), .A(w2170) );
	vdp_nor g2351 (.Z(w2034), .A(w2402), .B(w1156) );
	vdp_nor g2352 (.Z(w2136), .A(w2403), .B(w1156) );
	vdp_nor g2353 (.Z(w2149), .A(w2226), .B(w1156) );
	vdp_nor g2354 (.Z(w2156), .A(w2194), .B(w1156) );
	vdp_aon22 g2355 (.Z(w2221), .A2(w2226), .A1(w2225), .B2(w2220), .B1(w2219) );
	vdp_sr_bit g2356 (.D(w2221), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2222) );
	vdp_not g2357 (.nZ(w2220), .A(w2225) );
	vdp_not g2358 (.nZ(w2223), .A(w2222) );
	vdp_not g2359 (.nZ(w2359), .A(w1157) );
	vdp_not g2360 (.nZ(w2358), .A(w1158) );
	vdp_not g2361 (.nZ(w2259), .A(w2258) );
	vdp_sr_bit g2362 (.D(w2043), .nC1(w2212), .nC2(w2214), .C1(w2211), .C2(w2213), .Q(w2184) );
	vdp_nand g2363 (.Z(w2360), .A(w1157), .B(w2358) );
	vdp_nand g2364 (.Z(w2224), .A(w1158), .B(w1157) );
	vdp_nand g2365 (.Z(w2361), .A(w2358), .B(w2359) );
	vdp_nand g2366 (.Z(w2362), .A(w1158), .B(w2359) );
	vdp_and g2367 (.Z(w2228), .A(w2221), .B(w2223) );
	vdp_and g2368 (.Z(w2008), .A(w1156), .B(w2224) );
	vdp_and g2369 (.Z(w2010), .A(w1156), .B(w2360) );
	vdp_and g2370 (.Z(w2009), .A(w1156), .B(w2361) );
	vdp_and g2371 (.Z(w2007), .A(w1156), .B(w2362) );
	vdp_nor4 g2372 (.Z(w2232), .A(w2294), .B(w2307), .D(w2306), .C(w2194) );
	vdp_not g2373 (.nZ(w2229), .A(w2228) );
	vdp_not g2374 (.nZ(w2296), .A(w2230) );
	vdp_not g2375 (.nZ(w2295), .A(w2363) );
	vdp_not g2376 (.nZ(w2191), .A(w2259) );
	vdp_nand g2377 (.Z(w2230), .A(w2227), .B(w2229) );
	vdp_nand g2378 (.Z(w2363), .A(w2227), .B(w2228) );
	vdp_nor g2379 (.Z(w2227), .A(w2191), .B(w2231) );
	vdp_rs_ff g2380 (.S(w2218), .R(w2231), .Q(w2260) );
	vdp_rs_ff g2381 (.S(w2043), .R(w1060), .Q(w2233) );
	vdp_nor g2382 (.Z(w2234), .A(w1060), .B(w2233) );
	vdp_comp_dff g2383 (.D(w2234), .nC1(w2212), .C1(w2211), .C2(w2213), .nC2(w2214), .Q(w2043) );
	vdp_comp_dff g2384 (.D(SYSRES), .nC1(PSG_nCLK1), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC2(PSG_nCLK2), .Q(w2258) );
	vdp_comp_dff g2385 (.D(w2260), .nC1(PSG_nCLK1), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC2(PSG_nCLK2), .Q(w2231) );
	vdp_sr_bit g2386 (.Q(w2616), .D(w2610), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2387 (.nZ(AD_RD_DIR), .A(w2609) );
	vdp_sr_bit g2388 (.Q(w2617), .D(w2478), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2389 (.Q(w2544), .D(w2491), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2390 (.Q(w2600), .D(w33), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2391 (.Q(w2470), .D(w35), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2392 (.nZ(w2612), .A(w2468) );
	vdp_or g2393 (.Z(w2478), .A(w35), .B(w2470) );
	vdp_sr_bit g2394 (.Q(w2487), .D(w2489), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_sr_bit g2395 (.Q(w2613), .D(w2602), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2396 (.nZ(w2543), .A(w2613) );
	vdp_or g2397 (.Z(w2466), .A(w2470), .B(w2469) );
	vdp_sr_bit g2398 (.Q(w2469), .D(w551), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2399 (.Q(w2467), .D(w32), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2400 (.Q(w2604), .D(w2467), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2401 (.Q(w2603), .D(w2479), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2402 (.Q(w2598), .D(w2600), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2403 (.Q(w2615), .D(w2620), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_not g2404 (.nZ(w2594), .A(w2675) );
	vdp_not g2405 (.nZ(w2490), .A(128k) );
	vdp_sr_bit g2406 (.Q(w2479), .D(VRAM_REFRESH), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2407 (.nZ(w2551), .A(w2465) );
	vdp_not g2408 (.nZ(w2618), .A(w2605) );
	vdp_not g2409 (.nZ(w2485), .A(w2477) );
	vdp_oai21 g2410 (.Z(w2465), .B(w2485), .A1(w2618), .A2(w2606) );
	vdp_or g2411 (.Z(w2477), .A(w2612), .B(w2611) );
	vdp_or g2412 (.Z(w2610), .A(w2469), .B(w551) );
	vdp_not g2413 (.nZ(w2619), .A(w2471) );
	vdp_not g2414 (.nZ(w2667), .A(w2620) );
	vdp_dlatch_inv g2415 (.nQ(w2620), .D(w3), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2416 (.nQ(w2614), .D(w2486), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g2417 (.nQ(w2486), .D(w2615), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g2418 (.nQ(w2468), .D(w2466), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2419 (.nQ(w2611), .D(w2468), .C(HCLK2), .nC(nHCLK2) );
	vdp_dlatch_inv g2420 (.nQ(w2608), .D(w2607), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2421 (.nQ(w2605), .D(w2604), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2422 (.nQ(w2606), .D(w2605), .C(HCLK2), .nC(nHCLK2) );
	vdp_aon22 g2423 (.Z(nCAS1), .A1(w2486), .B1(w2475), .B2(1'b1), .A2(w2613) );
	vdp_and3 g2424 (.Z(nWE1), .A(w2474), .B(w2617), .C(w2475) );
	vdp_and3 g2425 (.Z(nWE0), .A(w2475), .B(w2474), .C(w2616) );
	vdp_aoi222 g2426 (.Z(w2609), .A1(1'b1), .B1(w2472), .B2(1'b1), .A2(w95), .C1(w2477), .C2(w2475) );
	vdp_aon333 g2427 (.Z(nOE1), .A1(w2551), .A2(w2615), .A3(w2475), .B1(w2608), .B2(w2608), .B3(w2619), .C1(w2608), .C2(w2608), .C3(w2472) );
	vdp_or3 g2428 (.Z(w2607), .A(w2602), .B(w2604), .C(w2467) );
	vdp_sr_bit g2429 (.Q(w2472), .D(w2667), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_dlatch_inv g2430 (.nQ(w2474), .D(w2472), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g2431 (.nQ(w2601), .D(w2474), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g2432 (.nQ(w2475), .D(w2473), .C(DCLK1), .nC(nDCLK1) );
	vdp_not g2433 (.nZ(w2473), .A(w2601) );
	vdp_nand g2434 (.Z(w2695), .A(w2601), .B(w2472) );
	vdp_nand g2435 (.Z(w2694), .A(w2472), .B(w2614) );
	vdp_nand g2436 (.Z(w2481), .A(w2615), .B(1'b1) );
	vdp_aoi33 g2437 (.Z(w2681), .A1(w2598), .A2(w34), .A3(w34), .B1(w2492), .B2(w2493), .B3(w3) );
	vdp_and g2438 (.Z(w2488), .A(w2475), .B(w2474) );
	vdp_not g2439 (.nZ(w2482), .A(w2544) );
	vdp_comp_strong g2440 (.nZ(w2499), .Z(w2498), .A(w2505) );
	vdp_comp_strong g2441 (.nZ(w2566), .Z(w2589), .A(w2590) );
	vdp_comp_strong g2442 (.nZ(w2500), .Z(w2545), .A(w2590) );
	vdp_comp_strong g2443 (.nZ(w2549), .Z(w2548), .A(w2505) );
	vdp_comp_strong g2444 (.nZ(w2506), .Z(w2550), .A(w2502) );
	vdp_comp_strong g2445 (.nZ(w2553), .Z(w2595), .A(w2502) );
	vdp_not g2446 (.nZ(w2508), .A(w2472) );
	vdp_not g2447 (.nZ(w2493), .A(w34) );
	vdp_not g2448 (.nZ(w2492), .A(w36) );
	vdp_comp_strong g2449 (.nZ(w2547), .Z(w6776), .A(w2488) );
	vdp_comp_strong g2450 (.nZ(w2483), .Z(w2591), .A(w2488) );
	vdp_or g2451 (.Z(w2602), .A(w2479), .B(w2603) );
	vdp_and g2452 (.Z(w2489), .A(128k), .B(HCLK1) );
	vdp_comp_we g2453 (.nZ(w2592), .Z(w2593), .A(w95) );
	vdp_comp_we g2454 (.nZ(w2501), .Z(w2679), .A(w2509) );
	vdp_not g2455 (.nZ(w2680), .A(w2544) );
	vdp_not g2456 (.nZ(w2504), .A(w2695) );
	vdp_not g2457 (.nZ(w6781), .A(w2694) );
	vdp_not g2458 (.nZ(w6782), .A(w2481) );
	vdp_comp_we g2459 (.nZ(w6783), .Z(w2597), .A(M5) );
	vdp_comp_we g2460 (.nZ(w2552), .Z(w2507), .A(128k) );
	vdp_and g2461 (.Z(w2491), .A(w105), .B(w3) );
	vdp_and g2462 (.Z(w2502), .A(w3), .B(HCLK1) );
	vdp_and g2463 (.Z(w2505), .A(HCLK2), .B(w2599) );
	vdp_and g2464 (.Z(w2590), .A(w3), .B(HCLK1) );
	vdp_oai21 g2465 (.Z(w2675), .A1(HCLK2), .A2(w2490), .B(DCLK1) );
	vdp_notif0 g2466 (.nZ(AD_DATA[0]), .A(w2496), .nE(w2482) );
	vdp_aon22 g2467 (.Z(nYS), .A1(VRAMA[16]), .A2(w2593), .B1(w2592), .B2(w2659) );
	vdp_aon22 g2468 (.Z(w2635), .A1(VRAMA[15]), .B1(w2592), .A2(w2593), .B2(w2573) );
	vdp_aon22 g2469 (.Z(w2633), .A1(VRAMA[14]), .B1(w2592), .A2(w2593), .B2(w2456) );
	vdp_aon22 g2470 (.Z(w2455), .A1(VRAMA[6]), .B1(w2592), .A2(w2593), .B2(w2634) );
	vdp_aon22 g2471 (.Z(w2447), .A1(VRAMA[7]), .B1(w2592), .A2(w2593), .B2(w2446) );
	vdp_aon22 g2472 (.Z(w2663), .A1(VRAMA[13]), .B1(w2592), .A2(w2593), .B2(w2464) );
	vdp_aon22 g2473 (.Z(w2632), .A1(VRAMA[5]), .B1(w2592), .A2(w2593), .B2(w2683) );
	vdp_aon22 g2474 (.Z(w2638), .A1(VRAMA[12]), .B1(w2592), .A2(w2593), .B2(w2533) );
	vdp_aon22 g2475 (.Z(w2462), .A1(VRAMA[4]), .B1(w2592), .A2(w2593), .B2(w2540) );
	vdp_aon22 g2476 (.Z(w2637), .A1(VRAMA[11]), .B1(w2592), .A2(w2593), .B2(w2688) );
	vdp_aon22 g2477 (.Z(w2572), .A1(VRAMA[3]), .B1(w2592), .A2(w2593), .B2(w2684) );
	vdp_aon22 g2478 (.Z(w2665), .A1(VRAMA[10]), .B1(w2592), .A2(w2593), .B2(w2585) );
	vdp_aon22 g2479 (.Z(w2571), .A1(VRAMA[2]), .B1(w2592), .A2(w2593), .B2(w2529) );
	vdp_aon22 g2480 (.Z(w2494), .A1(VRAMA[8]), .B1(w2592), .A2(w2593), .B2(w2497) );
	vdp_aon22 g2481 (.Z(w2686), .A1(VRAMA[0]), .B1(w2592), .A2(w2593), .B2(w2520) );
	vdp_aon22 g2482 (.Z(w2687), .A1(VRAMA[9]), .B1(w2592), .A2(w2593), .B2(w2567) );
	vdp_aon22 g2483 (.Z(w2523), .A1(VRAMA[1]), .B1(w2592), .A2(w2593), .B2(w2525) );
	vdp_notif0 g2484 (.nZ(AD_DATA[1]), .A(w2515), .nE(w2482) );
	vdp_notif0 g2485 (.nZ(AD_DATA[2]), .A(w2569), .nE(w2482) );
	vdp_notif0 g2486 (.nZ(AD_DATA[3]), .A(w2526), .nE(w2482) );
	vdp_notif0 g2487 (.nZ(AD_DATA[5]), .A(w2463), .nE(w2482) );
	vdp_notif0 g2488 (.nZ(AD_DATA[4]), .A(w2546), .nE(w2482) );
	vdp_notif0 g2489 (.nZ(AD_DATA[6]), .A(w2457), .nE(w2482) );
	vdp_notif0 g2490 (.nZ(AD_DATA[7]), .A(w2454), .nE(w2482) );
	vdp_slatch g2491 (.nQ(w2496), .D(w2495), .nC(w2483), .C(w2591) );
	vdp_slatch g2492 (.nQ(w2515), .D(w2514), .nC(w2483), .C(w2591) );
	vdp_slatch g2493 (.nQ(w2569), .D(w2522), .nC(w2483), .C(w2591) );
	vdp_slatch g2494 (.nQ(w2526), .D(w2527), .nC(w2483), .C(w2591) );
	vdp_slatch g2495 (.nQ(w2546), .D(w2480), .nC(w2483), .C(w2591) );
	vdp_slatch g2496 (.nQ(w2463), .D(w2664), .nC(w2483), .C(w2591) );
	vdp_slatch g2497 (.nQ(w2457), .D(w2535), .nC(w2483), .C(w2591) );
	vdp_slatch g2498 (.nQ(w2454), .D(w2636), .nC(w2483), .C(w2591) );
	vdp_slatch g2499 (.nQ(w2449), .D(w2448), .nC(w2547), .C(w6776) );
	vdp_slatch g2500 (.nQ(w2538), .D(w2534), .nC(w2547), .C(w6776) );
	vdp_slatch g2501 (.nQ(w2576), .D(w2676), .nC(w2547), .C(w6776) );
	vdp_slatch g2502 (.nQ(w2577), .D(w2461), .nC(w2547), .C(w6776) );
	vdp_slatch g2503 (.nQ(w2639), .D(w2536), .nC(w2547), .C(w6776) );
	vdp_slatch g2504 (.nQ(w2530), .D(w2528), .nC(w2547), .C(w6776) );
	vdp_slatch g2505 (.nQ(w2524), .D(w2570), .nC(w2547), .C(w6776) );
	vdp_slatch g2506 (.nQ(w2554), .D(w2666), .nC(w2547), .C(w6776) );
	vdp_slatch g2507 (.Q(w2497), .D(w2557), .nC(w2499), .C(w2498) );
	vdp_slatch g2508 (.Q(w2567), .D(w2690), .nC(w2499), .C(w2498) );
	vdp_slatch g2509 (.Q(w2688), .D(w2642), .nC(w2499), .C(w2498) );
	vdp_slatch g2510 (.Q(w2585), .D(w2568), .nC(w2499), .C(w2498) );
	vdp_slatch g2511 (.Q(w2464), .D(w2556), .nC(w2499), .C(w2498) );
	vdp_slatch g2512 (.Q(w2533), .D(w2643), .nC(w2499), .C(w2498) );
	vdp_slatch g2513 (.Q(w2573), .D(w2646), .nC(w2499), .C(w2498) );
	vdp_slatch g2514 (.Q(w2456), .D(w2555), .nC(w2499), .C(w2498) );
	vdp_slatch g2515 (.nQ(w2645), .D(w355), .nC(w2566), .C(w2589) );
	vdp_slatch g2516 (.nQ(w2647), .D(RD_DATA[6]), .nC(w2566), .C(w2589) );
	vdp_slatch g2517 (.nQ(w2644), .D(RD_DATA[5]), .nC(w2566), .C(w2589) );
	vdp_slatch g2518 (.nQ(w2692), .D(RD_DATA[4]), .nC(w2566), .C(w2589) );
	vdp_slatch g2519 (.nQ(w2641), .D(w321), .nC(w2566), .C(w2589) );
	vdp_slatch g2520 (.nQ(w2693), .D(RD_DATA[2]), .nC(w2566), .C(w2589) );
	vdp_slatch g2521 (.nQ(w2691), .D(RD_DATA[0]), .nC(w2566), .C(w2589) );
	vdp_slatch g2522 (.nQ(w2640), .D(RD_DATA[1]), .nC(w2566), .C(w2589) );
	vdp_notif0 g2523 (.nZ(w355), .A(w2449), .nE(w2680) );
	vdp_notif0 g2524 (.nZ(RD_DATA[6]), .A(w2538), .nE(w2680) );
	vdp_notif0 g2525 (.nZ(RD_DATA[5]), .A(w2576), .nE(w2680) );
	vdp_notif0 g2526 (.nZ(RD_DATA[4]), .A(w2577), .nE(w2680) );
	vdp_notif0 g2527 (.nZ(w321), .A(w2639), .nE(w2680) );
	vdp_notif0 g2528 (.nZ(RD_DATA[2]), .A(w2530), .nE(w2680) );
	vdp_notif0 g2529 (.nZ(RD_DATA[1]), .A(w2524), .nE(w2680) );
	vdp_notif0 g2530 (.nZ(RD_DATA[0]), .A(w2554), .nE(w2680) );
	vdp_slatch g2531 (.nQ(w2669), .D(AD_DATA[7]), .nC(w2500), .C(w2545) );
	vdp_slatch g2532 (.nQ(w2668), .D(AD_DATA[6]), .nC(w2500), .C(w2545) );
	vdp_slatch g2533 (.nQ(w2689), .D(AD_DATA[5]), .nC(w2500), .C(w2545) );
	vdp_slatch g2534 (.nQ(w2671), .D(AD_DATA[3]), .nC(w2500), .C(w2545) );
	vdp_slatch g2535 (.nQ(w2672), .D(AD_DATA[2]), .nC(w2500), .C(w2545) );
	vdp_slatch g2536 (.nQ(w2674), .D(AD_DATA[1]), .nC(w2500), .C(w2545) );
	vdp_slatch g2537 (.nQ(w2673), .D(AD_DATA[0]), .nC(w2500), .C(w2545) );
	vdp_slatch g2538 (.Q(w2453), .D(w2565), .nC(w2549), .C(w2548) );
	vdp_slatch g2539 (.Q(w2460), .D(w2564), .nC(w2549), .C(w2548) );
	vdp_slatch g2540 (.Q(w2537), .D(w2563), .nC(w2549), .C(w2548) );
	vdp_slatch g2541 (.Q(w2677), .D(w2560), .nC(w2549), .C(w2548) );
	vdp_slatch g2542 (.Q(w2588), .D(w2561), .nC(w2549), .C(w2548) );
	vdp_slatch g2543 (.Q(w2521), .D(w2559), .nC(w2549), .C(w2548) );
	vdp_slatch g2544 (.Q(w2575), .D(w2452), .nC(w2506), .C(w2550) );
	vdp_slatch g2545 (.Q(w2682), .D(w2459), .nC(w2506), .C(w2550) );
	vdp_slatch g2546 (.Q(w2649), .D(w2513), .nC(w2506), .C(w2550) );
	vdp_slatch g2547 (.Q(w2579), .D(w2512), .nC(w2506), .C(w2550) );
	vdp_slatch g2548 (.Q(w2586), .D(w2587), .nC(w2506), .C(w2550) );
	vdp_slatch g2549 (.Q(w2678), .D(w2518), .nC(w2506), .C(w2550) );
	vdp_slatch g2550 (.Q(w2584), .D(w2484), .nC(w2506), .C(w2550) );
	vdp_slatch g2551 (.Q(w2685), .D(w2519), .nC(w2506), .C(w2550) );
	vdp_slatch g2552 (.Q(w2596), .D(w2517), .nC(w2553), .C(w2595) );
	vdp_slatch g2553 (.Q(w2583), .D(w2700), .nC(w2553), .C(w2595) );
	vdp_slatch g2554 (.Q(w2531), .D(w2511), .nC(w2553), .C(w2595) );
	vdp_slatch g2555 (.Q(w2580), .D(w2696), .nC(w2553), .C(w2595) );
	vdp_slatch g2556 (.Q(w2541), .D(w2458), .nC(w2553), .C(w2595) );
	vdp_slatch g2557 (.Q(w2578), .D(w2510), .nC(w2553), .C(w2595) );
	vdp_slatch g2558 (.Q(w2539), .D(w2451), .nC(w2553), .C(w2595) );
	vdp_slatch g2559 (.Q(w2574), .D(w2450), .nC(w2553), .C(w2595) );
	vdp_sr_bit g2560 (.Q(w2509), .D(w34), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2561 (.nZ(w2707), .A(w106) );
	vdp_not g2562 (.nZ(w2581), .A(w2582) );
	vdp_not g2563 (.nZ(w6784), .A(M5) );
	vdp_not g2564 (.nZ(w2516), .A(w2508) );
	vdp_not g2565 (.nZ(w2471), .A(w2516) );
	vdp_aoi21 g2566 (.Z(w2582), .B(w2650), .A2(VRAMA[9]), .A1(w6784) );
	vdp_aoi22 g2567 (.Z(w2690), .A1(w2524), .B1(w2501), .B2(w2640), .A2(w2679) );
	vdp_aoi22 g2568 (.Z(w2642), .A1(w2639), .B1(w2501), .B2(w2641), .A2(w2679) );
	vdp_aoi22 g2569 (.Z(w2568), .A1(w2530), .B1(w2501), .B2(w2693), .A2(w2679) );
	vdp_aoi22 g2570 (.Z(w2556), .A1(w2576), .B1(w2501), .B2(w2644), .A2(w2679) );
	vdp_aoi22 g2571 (.Z(w2643), .A1(w2577), .B1(w2501), .B2(w2692), .A2(w2679) );
	vdp_aoi22 g2572 (.Z(w2646), .A1(w2449), .B1(w2501), .B2(w2645), .A2(w2679) );
	vdp_aoi22 g2573 (.Z(w2555), .A1(w2538), .B1(w2501), .B2(w2647), .A2(w2679) );
	vdp_slatch g2574 (.Q(w2503), .D(w2558), .nC(w2549), .C(w2548) );
	vdp_slatch g2575 (.nQ(w2670), .D(AD_DATA[4]), .nC(w2500), .C(w2545) );
	vdp_slatch g2576 (.Q(w2532), .D(w2562), .nC(w2549), .C(w2548) );
	vdp_aoi22 g2577 (.Z(w2558), .A1(w2496), .B1(w2501), .B2(w2673), .A2(w2679) );
	vdp_aoi22 g2578 (.Z(w2559), .A1(w2515), .B1(w2501), .B2(w2674), .A2(w2679) );
	vdp_aoi22 g2579 (.Z(w2560), .A1(w2569), .B1(w2501), .B2(w2672), .A2(w2679) );
	vdp_aoi22 g2580 (.Z(w2561), .A1(w2526), .B1(w2501), .B2(w2671), .A2(w2679) );
	vdp_aoi22 g2581 (.Z(w2562), .A1(w2546), .B1(w2501), .B2(w2670), .A2(w2679) );
	vdp_aoi22 g2582 (.Z(w2563), .A1(w2463), .B1(w2501), .B2(w2689), .A2(w2679) );
	vdp_aoi22 g2583 (.Z(w2565), .A1(w2454), .B1(w2501), .B2(w2669), .A2(w2679) );
	vdp_aoi22 g2584 (.Z(w2564), .A1(w2457), .B1(w2501), .B2(w2668), .A2(w2679) );
	vdp_aon22 g2585 (.Z(w2519), .A1(VRAMA[2]), .B1(w6783), .B2(VRAMA[1]), .A2(w2597) );
	vdp_aon22 g2586 (.Z(w2518), .A1(VRAMA[3]), .B1(w6783), .B2(VRAMA[2]), .A2(w2597) );
	vdp_aon22 g2587 (.Z(w2484), .A1(VRAMA[4]), .B1(w6783), .B2(VRAMA[3]), .A2(w2597) );
	vdp_aon22 g2588 (.Z(w2587), .A1(VRAMA[5]), .B1(w6783), .B2(VRAMA[4]), .A2(w2597) );
	vdp_aon22 g2589 (.Z(w2512), .A1(VRAMA[6]), .B1(w6783), .B2(VRAMA[5]), .A2(w2597) );
	vdp_aon22 g2590 (.Z(w2513), .A1(VRAMA[7]), .B1(w6783), .B2(VRAMA[6]), .A2(w2597) );
	vdp_aon22 g2591 (.Z(w2459), .A1(VRAMA[8]), .B1(w6783), .B2(VRAMA[7]), .A2(w2597) );
	vdp_aon22 g2592 (.Z(w2452), .A1(VRAMA[9]), .B1(w6783), .B2(VRAMA[8]), .A2(w2597) );
	vdp_and g2593 (.Z(w2650), .A(VRAMA[1]), .B(M5) );
	vdp_aon22 g2594 (.Z(w2450), .A1(w2648), .B1(w2552), .B2(VRAMA[15]), .A2(w2507) );
	vdp_aon22 g2595 (.Z(w2451), .A1(VRAMA[15]), .B1(w2552), .B2(VRAMA[14]), .A2(w2507) );
	vdp_aon22 g2596 (.Z(w2458), .A1(VRAMA[14]), .B1(w2552), .B2(VRAMA[13]), .A2(w2507) );
	vdp_aon22 g2597 (.Z(w2696), .A1(VRAMA[12]), .B1(w2552), .B2(VRAMA[11]), .A2(w2507) );
	vdp_aon22 g2598 (.Z(w2510), .A1(VRAMA[13]), .B1(w2552), .B2(VRAMA[12]), .A2(w2507) );
	vdp_aon22 g2599 (.Z(w2511), .A1(VRAMA[11]), .B1(w2552), .B2(VRAMA[10]), .A2(w2507) );
	vdp_aon22 g2600 (.Z(w2700), .A1(VRAMA[10]), .B1(w2552), .B2(w2581), .A2(w2507) );
	vdp_aon22 g2601 (.Z(w2517), .A1(w2650), .B1(w2552), .B2(VRAMA[0]), .A2(w2507) );
	vdp_aon22 g2602 (.Z(w2648), .A1(w2707), .B1(w106), .B2(w89), .A2(VRAMA[16]) );
	vdp_aon222 g2603 (.Z(w2520), .A1(w2504), .A2(w2503), .B1(w6781), .B2(w2685), .C1(w6782), .C2(w2596) );
	vdp_aon222 g2604 (.Z(w2525), .A1(w2504), .A2(w2521), .B1(w6781), .B2(w2678), .C1(w6782), .C2(w2583) );
	vdp_aon222 g2605 (.Z(w2529), .A1(w2504), .A2(w2677), .B1(w6781), .B2(w2584), .C1(w6782), .C2(w2531) );
	vdp_aon222 g2606 (.Z(w2684), .A1(w2504), .A2(w2588), .B1(w6781), .B2(w2586), .C1(w6782), .C2(w2580) );
	vdp_aon222 g2607 (.Z(w2540), .A1(w2504), .A2(w2532), .B1(w6781), .B2(w2579), .C1(w6782), .C2(w2578) );
	vdp_aon222 g2608 (.Z(w2683), .A1(w2504), .A2(w2537), .B1(w6781), .B2(w2649), .C1(w6782), .C2(w2541) );
	vdp_aon222 g2609 (.Z(w2634), .A1(w2504), .A2(w2460), .B1(w6781), .B2(w2682), .C1(w6782), .C2(w2539) );
	vdp_aon222 g2610 (.Z(w2446), .A1(w2504), .A2(w2453), .B1(w6781), .B2(w2575), .C1(w6782), .C2(w2574) );
	vdp_dlatch_inv g2611 (.nQ(w2599), .D(w2681), .C(HCLK1), .nC(nHCLK1) );
	vdp_comp_we g2612 (.Z(w2542), .A(w2601) );
	vdp_aon22 g2613 (.Z(nRAS1), .A1(1'b1), .B1(w2543), .B2(w2486), .A2(w2542) );
	vdp_aoi22 g2614 (.Z(w2557), .A1(w2554), .B1(w2501), .B2(w2691), .A2(w2679) );
	vdp_and g2615 (.Z(w2621), .B(w2705), .A(DCLK2) );
	vdp_nor g2616 (.Z(w2701), .A(w2623), .B(RES) );
	vdp_sr_bit g2617 (.Q(w2623), .D(w2701), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_dlatch_inv g2618 (.nQ(w2702), .D(w2624), .C(DCLK1), .nC(nDCLK1) );
	vdp_and g2619 (.Z(w2703), .A(DCLK2), .B(w2702) );
	vdp_dlatch_inv g2620 (.nQ(w2705), .D(w2623), .C(DCLK1), .nC(nDCLK1) );
	vdp_not g2621 (.nZ(w2627), .A(w2629) );
	vdp_not g2622 (.nZ(w2626), .A(w2704) );
	vdp_neg_dff g2623 (.Q(w2629), .C(DCLK1), .D(1'b1), .R(w2621) );
	vdp_not g2624 (.A(w2623), .nZ(w2624) );
	vdp_neg_dff g2625 (.Q(w2704), .R(w2703), .C(DCLK1), .D(1'b1) );
	vdp_sr_bit g2626 (.Q(w2782), .D(w2774), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2627 (.Q(w2778), .D(w2777), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2628 (.Q(w2973), .D(w2778), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2629 (.Q(w2796), .D(w2973), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2630 (.Q(w2751), .D(RD_DATA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2631 (.Q(w2752), .D(RD_DATA[2]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2632 (.Q(w2753), .D(w321), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2633 (.Q(w2954), .D(w2976), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2634 (.Q(w2976), .D(w2977), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2635 (.Q(w2977), .D(w2978), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2636 (.Q(w2978), .D(w2979), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2637 (.Q(w2979), .D(w2980), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2638 (.Q(w2980), .D(w2981), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2639 (.Q(w2981), .D(w2982), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2640 (.Q(w2982), .D(w18), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2641 (.Q(w2760), .D(w2788), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2642 (.Q(w2758), .D(w2985), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2643 (.Q(w3013), .D(w2987), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2644 (.Q(w2987), .D(w2734), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2645 (.Q(w2734), .D(w103), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2646 (.Q(w2709), .D(w2708), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2647 (.Q(w2714), .D(w2857), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2648 (.Q(w2772), .D(w2969), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2649 (.Q(w2776), .D(w2984), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2650 (.Q(w2792), .D(w2784), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2651 (.Q(w2708), .D(w2787), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2652 (.Q(w2813), .D(w2790), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2653 (.Q(w2812), .D(w2858), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2654 (.Q(PLANE_A_PRIO), .D(w2804), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2655 (.Q(PLANE_B_PRIO), .D(w2805), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2656 (.Q(w2768), .D(w2806), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2657 (.Q(w2811), .D(w2810), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2658 (.Q(w2730), .D(w2809), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2659 (.Q(w2809), .D(w125), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2660 (.Q(w2731), .D(w3015), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2661 (.Q(w3015), .D(w124), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2662 (.Q(w2822), .D(w2795), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2663 (.Q(w2808), .D(w2807), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2664 (.Q(SPR_PRIO), .D(w2961), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2665 (.Q(w2819), .D(w173), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2666 (.Q(w2818), .D(w172), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2667 (.Q(w2723), .D(w2739), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2668 (.Q(w2728), .D(w2740), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2669 (.Q(w2725), .D(w2750), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2670 (.Q(w2716), .D(w2741), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2671 (.Q(w2735), .D(w2748), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2672 (.Q(w2715), .D(w2742), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2673 (.Q(w2710), .D(w2845), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2674 (.Q(w2720), .D(w2743), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2675 (.Q(w2726), .D(w2737), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_slatch g2676 (.nQ(w3011), .D(w2739), .C(w2736), .nC(w2733) );
	vdp_slatch g2677 (.nQ(w3012), .D(w2737), .C(w2736), .nC(w2733) );
	vdp_slatch g2678 (.nQ(w3010), .D(w2740), .C(w2736), .nC(w2733) );
	vdp_slatch g2679 (.nQ(w3009), .D(w2750), .C(w2736), .nC(w2733) );
	vdp_slatch g2680 (.nQ(w3008), .D(w2741), .C(w2736), .nC(w2733) );
	vdp_slatch g2681 (.nQ(w3007), .D(w2748), .C(w2736), .nC(w2733) );
	vdp_slatch g2682 (.nQ(w3006), .D(w2742), .C(w2736), .nC(w2733) );
	vdp_slatch g2683 (.nQ(w3005), .D(w2845), .C(w2736), .nC(w2733) );
	vdp_slatch g2684 (.nQ(w3004), .D(w2743), .C(w2736), .nC(w2733) );
	vdp_slatch g2685 (.Q(w2794), .D(REG_BUS[7]), .nC(w2771), .C(w2781) );
	vdp_slatch g2686 (.Q(w2791), .D(REG_BUS[5]), .nC(w2771), .C(w2781) );
	vdp_slatch g2687 (.Q(w2783), .D(REG_BUS[4]), .nC(w2771), .C(w2781) );
	vdp_slatch g2688 (.Q(w2779), .D(REG_BUS[3]), .nC(w2771), .C(w2781) );
	vdp_slatch g2689 (.Q(w2775), .D(REG_BUS[2]), .nC(w2771), .C(w2781) );
	vdp_slatch g2690 (.Q(w2972), .D(REG_BUS[1]), .nC(w2771), .C(w2781) );
	vdp_slatch g2691 (.Q(w2773), .D(REG_BUS[0]), .nC(w2771), .C(w2781) );
	vdp_slatch g2692 (.Q(w2947), .D(REG_BUS[6]), .nC(w2771), .C(w2781) );
	vdp_aon2222 g2693 (.Z(w2924), .B2(w2863), .B1(w2868), .A2(w2999), .A1(w2863), .D2(w2859), .D1(w2868), .C2(w2868), .C1(w2860) );
	vdp_aon22 g2694 (.Z(w2889), .B2(w2859), .B1(w2873), .A2(w3000), .A1(w2864) );
	vdp_aon22 g2695 (.Z(w2894), .B2(w2859), .B1(w2869), .A2(w2999), .A1(w2864) );
	vdp_not g2696 (.nZ(w2877), .A(w2923) );
	vdp_not g2697 (.nZ(w2871), .A(w2872) );
	vdp_not g2698 (.nZ(w2876), .A(w2875) );
	vdp_not g2699 (.nZ(w2895), .A(w2924) );
	vdp_not g2700 (.nZ(w2888), .A(w2881) );
	vdp_buf g2701 (.Z(w2863), .A(w2758) );
	vdp_not g2702 (.nZ(w2958), .A(w2916) );
	vdp_not g2703 (.nZ(w2919), .A(w2917) );
	vdp_not g2704 (.nZ(w2920), .A(w2921) );
	vdp_not g2705 (.nZ(w2884), .A(w2860) );
	vdp_sr_bit g2706 (.Q(w2883), .D(w2731), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2707 (.Q(w2921), .D(w2729), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2708 (.Q(w2860), .D(w2730), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2709 (.Q(w2916), .D(w2918), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2710 (.Q(w2917), .D(w2754), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g2711 (.Z(w2995), .A(w2920), .B(w2958), .C(w2917) );
	vdp_and3 g2712 (.Z(w2997), .A(w2919), .B(w2921), .C(w2958) );
	vdp_and3 g2713 (.Z(w2996), .A(w2920), .B(w2958), .C(w2919) );
	vdp_and3 g2714 (.Z(w2882), .A(w2958), .B(w2917), .C(w2921) );
	vdp_and3 g2715 (.Z(w2880), .A(w2920), .B(w2916), .C(w2919) );
	vdp_and3 g2716 (.Z(w2878), .A(w2916), .B(w2917), .C(w2921) );
	vdp_and3 g2717 (.Z(w2998), .A(w2920), .B(w2917), .C(w2916) );
	vdp_and3 g2718 (.Z(w2879), .A(w2919), .B(w2921), .C(w2916) );
	vdp_sr_bit g2719 (.Q(w2875), .D(w2922), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2720 (.Q(w2872), .D(w2719), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2721 (.Q(w2923), .D(w2755), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g2722 (.Z(w2874), .A(w2876), .B(w2877), .C(w2871) );
	vdp_and3 g2723 (.Z(w2873), .A(w2871), .B(w2875), .C(w2877) );
	vdp_and3 g2724 (.Z(w3000), .A(w2876), .B(w2877), .C(w2872) );
	vdp_and3 g2725 (.Z(w2869), .A(w2877), .B(w2872), .C(w2875) );
	vdp_and3 g2726 (.Z(w2870), .A(w2871), .B(w2875), .C(w2923) );
	vdp_and3 g2727 (.Z(w2867), .A(w2876), .B(w2923), .C(w2871) );
	vdp_and3 g2728 (.Z(w2999), .A(w2876), .B(w2872), .C(w2923) );
	vdp_and3 g2729 (.Z(w2868), .A(w2923), .B(w2872), .C(w2875) );
	vdp_not g2730 (.nZ(w2957), .A(w3014) );
	vdp_not g2731 (.nZ(w2912), .A(w2914) );
	vdp_not g2732 (.nZ(w2913), .A(w2915) );
	vdp_sr_bit g2733 (.Q(w2914), .D(w2953), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2734 (.Q(w2915), .D(w2951), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2735 (.Q(w3014), .D(w2717), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g2736 (.Z(w2866), .A(w2913), .B(w2957), .C(w2912) );
	vdp_and3 g2737 (.Z(w2865), .A(w2912), .B(w2915), .C(w2957) );
	vdp_and3 g2738 (.A(w2913), .B(w2957), .C(w2914), .Z(w2862) );
	vdp_and3 g2739 (.Z(w3001), .A(w2957), .B(w2914), .C(w2915) );
	vdp_and3 g2740 (.Z(w2861), .A(w2913), .B(w3014), .C(w2912) );
	vdp_and3 g2741 (.Z(w3003), .A(w2912), .B(w2915), .C(w3014) );
	vdp_and3 g2742 (.Z(w2956), .A(w3014), .B(w2914), .C(w2915) );
	vdp_and3 g2743 (.Z(w3002), .A(w2913), .B(w2914), .C(w3014) );
	vdp_aon22 g2744 (.nZ(w2946), .B2(w2859), .B1(w3002), .A2(w3003), .A1(w2860) );
	vdp_aon22 g2745 (.nZ(w2911), .B2(w2859), .B1(w2861), .A2(w2865), .A1(w2860) );
	vdp_aon22 g2746 (.nZ(w2945), .B2(w2860), .B1(w2866), .A2(w2956), .A1(w2864) );
	vdp_and g2747 (.nZ(w2910), .B(w2860), .A(w2861) );
	vdp_and g2748 (.nZ(w2944), .B(w2860), .A(w3002) );
	vdp_and g2749 (.nZ(w2943), .B(w2860), .A(w2862) );
	vdp_aon22 g2750 (.nZ(w2942), .B2(w2863), .B1(w3003), .A2(w2861), .A1(w2863) );
	vdp_aon22 g2751 (.nZ(w2941), .B2(w2859), .B1(w3003), .A2(w3001), .A1(w2860) );
	vdp_aon2222 g2752 (.Z(w2925), .B2(w2863), .B1(w2956), .A2(w3002), .A1(w2863), .D2(w2859), .D1(w2956), .C2(w2956), .C1(w2860) );
	vdp_aon22 g2753 (.Z(w2908), .B2(w2859), .B1(w2865), .A2(w2862), .A1(w2864) );
	vdp_aon22 g2754 (.Z(w2905), .B2(w2859), .B1(w3001), .A2(w3002), .A1(w2864) );
	vdp_and g2755 (.Z(w2909), .B(w3003), .A(w2864) );
	vdp_and g2756 (.Z(w2904), .B(w2864), .A(w3001) );
	vdp_and g2757 (.Z(w2906), .B(w2865), .A(w2864) );
	vdp_aon22 g2758 (.Z(w2903), .B2(w2863), .B1(w3001), .A2(w2862), .A1(w2863) );
	vdp_aon22 g2759 (.Z(w2902), .B2(w2859), .B1(w2862), .A2(w2861), .A1(w2864) );
	vdp_aon2222 g2760 (.Z(w2940), .B2(w2863), .B1(w2865), .A2(w2866), .A1(w2863), .D2(w2859), .D1(w2866), .C2(w2866), .C1(w2864) );
	vdp_not g2761 (.nZ(w2907), .A(w2925) );
	vdp_aon22 g2762 (.nZ(w2939), .B2(w2859), .B1(w2999), .A2(w2870), .A1(w2860) );
	vdp_aon22 g2763 (.nZ(w2938), .B2(w2859), .B1(w2867), .A2(w2873), .A1(w2860) );
	vdp_aon22 g2764 (.nZ(w2901), .B2(w2860), .B1(w2874), .A2(w2868), .A1(w2864) );
	vdp_and g2765 (.nZ(w2900), .B(w2860), .A(w2867) );
	vdp_and g2766 (.nZ(w2899), .B(w2860), .A(w2999) );
	vdp_and g2767 (.nZ(w2898), .B(w2860), .A(w3000) );
	vdp_aon22 g2768 (.nZ(w2897), .B2(w2863), .B1(w2870), .A2(w2867), .A1(w2863) );
	vdp_aon22 g2769 (.nZ(w2896), .B2(w2859), .B1(w2870), .A2(w2869), .A1(w2860) );
	vdp_and g2770 (.Z(w2893), .B(w2870), .A(w2864) );
	vdp_and g2771 (.Z(w2992), .B(w2864), .A(w2869) );
	vdp_and g2772 (.Z(w2892), .B(w2873), .A(w2864) );
	vdp_aon22 g2773 (.Z(w2891), .B2(w2863), .B1(w2869), .A2(w3000), .A1(w2863) );
	vdp_aon22 g2774 (.Z(w2890), .B2(w2859), .B1(w3000), .A2(w2867), .A1(w2864) );
	vdp_aon2222 g2775 (.Z(w2993), .B2(w2863), .B1(w2873), .A2(w2874), .A1(w2863), .D2(w2859), .D1(w2874), .C2(w2874), .C1(w2864) );
	vdp_aon22 g2776 (.nZ(w2887), .B2(w2859), .B1(w2998), .A2(w2879), .A1(w2860) );
	vdp_aon22 g2777 (.nZ(w2937), .B2(w2859), .B1(w2880), .A2(w2997), .A1(w2860) );
	vdp_aon22 g2778 (.nZ(w2933), .B2(w2860), .B1(w2996), .A2(w2878), .A1(w2864) );
	vdp_and g2779 (.nZ(w2934), .B(w2860), .A(w2880) );
	vdp_and g2780 (.nZ(w2935), .B(w2860), .A(w2998) );
	vdp_and g2781 (.nZ(w2932), .B(w2860), .A(w2995) );
	vdp_aon22 g2782 (.nZ(w2936), .B2(w2863), .B1(w2879), .A2(w2880), .A1(w2863) );
	vdp_aon22 g2783 (.nZ(w2994), .B2(w2859), .B1(w2879), .A2(w2882), .A1(w2860) );
	vdp_aon2222 g2784 (.Z(w2881), .B2(w2863), .B1(w2878), .A2(w2998), .A1(w2863), .D2(w2859), .D1(w2878), .C2(w2878), .C1(w2860) );
	vdp_aon22 g2785 (.Z(w2885), .B2(w2859), .B1(w2997), .A2(w2995), .A1(w2864) );
	vdp_aon22 g2786 (.Z(w2886), .B2(w2863), .B1(w2882), .A2(w2995), .A1(w2863) );
	vdp_aon22 g2787 (.Z(w2931), .B2(w2859), .B1(w2882), .A2(w2998), .A1(w2864) );
	vdp_and g2788 (.Z(w2930), .B(w2864), .A(w2882) );
	vdp_and g2789 (.Z(w2929), .B(w2997), .A(w2864) );
	vdp_and g2790 (.Z(w2928), .B(w2864), .A(w2879) );
	vdp_aon22 g2791 (.Z(w2926), .B2(w2859), .B1(w2995), .A2(w2880), .A1(w2864) );
	vdp_aon2222 g2792 (.Z(w2927), .B2(w2863), .B1(w2997), .A2(w2996), .A1(w2863), .D2(w2859), .D1(w2996), .C2(w2996), .C1(w2864) );
	vdp_nor3 g2793 (.Z(w2859), .A(w2863), .B(w2883), .C(w2860) );
	vdp_and g2794 (.Z(w2864), .A(w2883), .B(w2884) );
	vdp_bufif0 g2795 (.A(w2773), .nE(w2780), .Z(COL[0]) );
	vdp_bufif0 g2796 (.A(w2972), .nE(w2780), .Z(COL[1]) );
	vdp_bufif0 g2797 (.A(w2775), .nE(w2780), .Z(COL[2]) );
	vdp_bufif0 g2798 (.A(w2779), .nE(w2780), .Z(COL[3]) );
	vdp_bufif0 g2799 (.A(w2793), .nE(w2780), .Z(COL[4]) );
	vdp_bufif0 g2800 (.A(w2971), .nE(w2780), .Z(COL[5]) );
	vdp_and g2801 (.Z(w2971), .A(M5), .B(w2791) );
	vdp_or g2802 (.Z(w2793), .A(w2763), .B(w2783) );
	vdp_not g2803 (.nZ(w2659), .A(M5) );
	vdp_not g2804 (.nZ(w2761), .A(w2970) );
	vdp_not g2805 (.nZ(w2762), .A(w2764) );
	vdp_not g2806 (.nZ(w2763), .A(M5) );
	vdp_not g2807 (.nZ(w2759), .A(w2765) );
	vdp_not g2808 (.nZ(w2780), .A(w2768) );
	vdp_comp_strong g2809 (.nZ(w2771), .Z(w2781), .A(w73) );
	vdp_not g2810 (.nZ(w2769), .A(w96) );
	vdp_not g2811 (.nZ(w2983), .A(w19) );
	vdp_aon222 g2812 (.Z(w2969), .B2(w2761), .A2(w2762), .A1(VRAMA[0]), .B1(VRAMA[1]), .C2(w2759), .C1(COL[0]) );
	vdp_aon222 g2813 (.Z(w2984), .B2(w2761), .A2(w2762), .A1(VRAMA[1]), .B1(VRAMA[2]), .C2(w2759), .C1(COL[1]) );
	vdp_aon222 g2814 (.Z(w2774), .B2(w2761), .A2(w2762), .A1(VRAMA[2]), .B1(VRAMA[3]), .C2(w2759), .C1(COL[2]) );
	vdp_aon222 g2815 (.Z(w2784), .B2(w2761), .A2(w2762), .A1(VRAMA[3]), .B1(VRAMA[4]), .C2(w2759), .C1(COL[3]) );
	vdp_aon222 g2816 (.Z(w2790), .B2(w2761), .A2(w2762), .A1(VRAMA[4]), .B1(VRAMA[5]), .C2(w2759), .C1(COL[4]) );
	vdp_aon222 g2817 (.Z(w2858), .B2(w2761), .A2(w2762), .A1(1'b0), .B1(VRAMA[6]), .C2(w2759), .C1(COL[5]) );
	vdp_nand g2818 (.Z(w2970), .A(w2765), .B(M5) );
	vdp_nand g2819 (.Z(w2764), .A(w2765), .B(w2763) );
	vdp_and g2820 (.Z(w2795), .A(w2796), .B(w3022) );
	vdp_aon222 g2821 (.Z(w3022), .B2(w3017), .A2(w2801), .A1(w2756), .B1(w2803), .C2(w3016), .C1(w2824) );
	vdp_not g2822 (.nZ(w3017), .A(w2968) );
	vdp_not g2823 (.nZ(w3016), .A(w2757) );
	vdp_not g2824 (.nZ(w2829), .A(w2814) );
	vdp_nor g2825 (.Z(w2803), .A(w2757), .B(w2961) );
	vdp_nor g2826 (.Z(w2968), .A(w2824), .B(w2823) );
	vdp_and g2827 (.Z(w2802), .A(w2797), .B(w2837) );
	vdp_and g2828 (.Z(w2801), .A(w2814), .B(w2828) );
	vdp_and g2829 (.Z(w2831), .A(w2828), .B(w2829) );
	vdp_or g2830 (.Z(w2961), .A(w2832), .B(w2831) );
	vdp_or g2831 (.Z(w2800), .A(w2756), .B(w2757) );
	vdp_and g2832 (.Z(w2770), .A(w2796), .B(w2769) );
	vdp_and g2833 (.Z(w2950), .A(w2797), .B(w2834) );
	vdp_and g2834 (.Z(w2960), .A(w2798), .B(w2836) );
	vdp_not g2835 (.nZ(w2842), .A(w96) );
	vdp_or g2836 (.Z(w2804), .A(w2835), .B(w2821) );
	vdp_not g2837 (.nZ(w3020), .A(w2798) );
	vdp_not g2838 (.nZ(w2948), .A(w2698) );
	vdp_not g2839 (.nZ(w2826), .A(w2815) );
	vdp_not g2840 (.nZ(w2825), .A(w2816) );
	vdp_not g2841 (.nZ(w2830), .A(w2699) );
	vdp_and g2842 (.Z(w2849), .A(w2798), .B(w2833) );
	vdp_and g2843 (.Z(w2827), .A(w2799), .B(w2839) );
	vdp_not g2844 (.nZ(w2959), .A(w93) );
	vdp_not g2845 (.nZ(w2966), .A(w94) );
	vdp_and g2846 (.Z(w2832), .A(w2966), .B(w93) );
	vdp_and g2847 (.Z(w2835), .A(w2959), .B(w94) );
	vdp_and g2848 (.Z(w2848), .A(w93), .B(w94) );
	vdp_or3 g2849 (.Z(w2765), .A(w103), .B(w172), .C(w173) );
	vdp_and3 g2850 (.Z(w2965), .A(w2799), .B(w2798), .C(w2836) );
	vdp_and3 g2851 (.Z(w2834), .A(w2825), .B(w2815), .C(w2699) );
	vdp_and3 g2852 (.Z(w2833), .A(w2826), .B(w2816), .C(w2830) );
	vdp_and3 g2853 (.Z(w2839), .A(w2825), .B(w2815), .C(w2830) );
	vdp_and3 g2854 (.Z(w2836), .A(w2815), .B(w2816), .C(w2830) );
	vdp_and g2855 (.Z(w2955), .A(M5), .B(w84) );
	vdp_or g2856 (.Z(w2797), .A(w2948), .B(w2814) );
	vdp_and3 g2857 (.Z(w2807), .A(w2801), .B(w2757), .C(w2968) );
	vdp_and3 g2858 (.Z(w2964), .A(w2799), .B(w2797), .C(w2834) );
	vdp_and3 g2859 (.Z(w2963), .A(w2799), .B(w2797), .C(w2839) );
	vdp_and3 g2860 (.Z(w2821), .A(w2820), .B(w2770), .C(w3020) );
	vdp_and3 g2861 (.Z(w2814), .A(w2800), .B(w2817), .C(w2955) );
	vdp_and3 g2862 (.Z(w2843), .A(w2798), .B(w2797), .C(w2837) );
	vdp_and3 g2863 (.Z(w3019), .A(w2798), .B(w2797), .C(w2833) );
	vdp_and3 g2864 (.Z(w2840), .A(w2799), .B(w2798), .C(w2797) );
	vdp_and3 g2865 (.Z(w2841), .A(w2770), .B(w2838), .C(w3018) );
	vdp_and g2866 (.Z(w2806), .A(w2949), .B(w2962) );
	vdp_not g2867 (.nZ(w2844), .A(w2770) );
	vdp_not g2868 (.nZ(w3018), .A(w2799) );
	vdp_or g2869 (.Z(w2805), .A(w2848), .B(w2841) );
	vdp_or g2870 (.Z(w2962), .A(w2844), .B(w2840) );
	vdp_not g2871 (.nZ(w2975), .A(M5) );
	vdp_notif0 g2872 (.A(w3012), .nE(w2738), .nZ(w321) );
	vdp_notif0 g2873 (.nZ(RD_DATA[2]), .A(w3011), .nE(w2738) );
	vdp_notif0 g2874 (.nZ(RD_DATA[1]), .A(w3010), .nE(w2738) );
	vdp_notif0 g2875 (.nZ(AD_DATA[7]), .A(w3009), .nE(w2738) );
	vdp_notif0 g2876 (.nZ(AD_DATA[6]), .A(w3008), .nE(w2738) );
	vdp_notif0 g2877 (.nZ(AD_DATA[5]), .A(w3007), .nE(w2738) );
	vdp_notif0 g2878 (.nZ(AD_DATA[3]), .A(w3006), .nE(w2738) );
	vdp_notif0 g2879 (.nZ(AD_DATA[2]), .A(w3005), .nE(w2738) );
	vdp_notif0 g2880 (.nZ(AD_DATA[1]), .A(w3004), .nE(w2738) );
	vdp_notif0 g2881 (.nZ(DB[1]), .A(w2731), .nE(w2722) );
	vdp_notif0 g2882 (.A(w2730), .nE(w2722) );
	vdp_notif0 g2883 (.nZ(DB[2]), .A(w2951), .nE(w2722) );
	vdp_notif0 g2884 (.nZ(DB[5]), .A(w2922), .nE(w2722) );
	vdp_notif0 g2885 (.nZ(DB[8]), .A(w2729), .nE(w2722) );
	vdp_notif0 g2886 (.nZ(DB[10]), .A(w2918), .nE(w2722) );
	vdp_notif0 g2887 (.nZ(DB[9]), .A(w2754), .nE(w2722) );
	vdp_notif0 g2888 (.nZ(DB[7]), .A(w2755), .nE(w2722) );
	vdp_notif0 g2889 (.nZ(DB[6]), .A(w2719), .nE(w2722) );
	vdp_notif0 g2890 (.nZ(DB[4]), .A(w2717), .nE(w2722) );
	vdp_comp_we g2891 (.A(M5), .nZ(w2712), .Z(w2711) );
	vdp_notif0 g2892 (.nZ(DB[3]), .A(w2953), .nE(w2722) );
	vdp_not g2893 (.A(w83), .nZ(w2722) );
	vdp_and g2894 (.Z(w2713), .A(w2714), .B(w2709) );
	vdp_and3 g2895 (.Z(w2953), .A(w92), .B(w2714), .C(w2952) );
	vdp_and3 g2896 (.Z(w2717), .A(w92), .B(w2714), .C(w2986) );
	vdp_and3 g2897 (.Z(w2719), .A(w92), .B(w2714), .C(w2718) );
	vdp_and3 g2898 (.Z(w2755), .A(w92), .B(w2714), .C(w2721) );
	vdp_and3 g2899 (.Z(w2754), .A(w92), .B(w2714), .C(w2724) );
	vdp_and3 g2900 (.Z(w2918), .A(w92), .B(w2714), .C(w2727) );
	vdp_and3 g2901 (.Z(w2729), .A(M5), .B(w2714), .C(w2728) );
	vdp_and3 g2902 (.Z(w2922), .A(M5), .B(w2714), .C(w2735) );
	vdp_and3 g2903 (.Z(w2951), .A(M5), .B(w2714), .C(w2720) );
	vdp_comp_strong g2904 (.nZ(w2733), .A(w2732), .Z(w2736) );
	vdp_and g2905 (.Z(w2732), .A(w2734), .B(HCLK1) );
	vdp_not g2906 (.nZ(w2738), .A(w3013) );
	vdp_aon22 g2907 (.Z(w2974), .B2(FIFOo[5]), .A2(FIFOo[7]), .A1(w2786), .B1(w2785) );
	vdp_aon22 g2908 (.Z(w2749), .B2(FIFOo[4]), .A2(FIFOo[6]), .A1(w2786), .B1(w2785) );
	vdp_aon22 g2909 (.Z(w2747), .B2(FIFOo[3]), .A2(FIFOo[5]), .A1(w2786), .B1(w2785) );
	vdp_aon22 g2910 (.Z(w2746), .B2(FIFOo[2]), .A2(FIFOo[3]), .A1(w2786), .B1(w2785) );
	vdp_aon22 g2911 (.Z(w2745), .B2(FIFOo[1]), .A2(FIFOo[2]), .A1(w2786), .B1(w2785) );
	vdp_aon22 g2912 (.Z(w2744), .B2(FIFOo[0]), .A2(FIFOo[1]), .A1(w2786), .B1(w2785) );
	vdp_comp_we g2913 (.Z(w2786), .nZ(w2785), .A(M5) );
	vdp_aon22 g2914 (.Z(w2777), .B2(w2975), .A2(M5), .A1(w2954), .B1(w18) );
	vdp_aon22 g2915 (.Z(w125), .B2(w2808), .A2(w2794), .A1(w96), .B1(w2842) );
	vdp_aon22 g2916 (.Z(w124), .B2(w2822), .A2(w2947), .A1(w96), .B1(w2842) );
	vdp_and3 g2917 (.Z(w2828), .A(w2770), .B(w2698), .C(w3021) );
	vdp_aon22 g2918 (.Z(w2837), .B2(w2825), .A2(w2816), .A1(w2699), .B1(w2826) );
	vdp_aon22 g2919 (.Z(w2721), .B2(w2735), .A2(w2725), .A1(w2711), .B1(w2712) );
	vdp_aon22 g2920 (.Z(w2718), .B2(w2715), .A2(w2716), .A1(w2711), .B1(w2712) );
	vdp_aon22 g2921 (.Z(w2952), .B2(w2720), .A2(w2710), .A1(w2711), .B1(w2712) );
	vdp_aon22 g2922 (.Z(w2986), .B2(w2710), .A2(w2715), .A1(w2711), .B1(w2712) );
	vdp_aon22 g2923 (.Z(w2724), .B2(w2716), .A2(w2723), .A1(w2711), .B1(w2712) );
	vdp_aon22 g2924 (.Z(w2727), .B2(w2725), .A2(w2726), .A1(w2711), .B1(w2712) );
	vdp_and4 g2925 (.Z(w2823), .A(w2826), .B(w2699), .C(w2955), .D(w2825) );
	vdp_or5 g2926 (.Z(w2820), .A(w2802), .B(w2833), .C(w2836), .D(w2964), .E(w2963) );
	vdp_or5 g2927 (.Z(w2838), .A(w2843), .B(w2839), .C(w2950), .D(w2960), .E(w3019) );
	vdp_or5 g2928 (.Z(w3021), .A(w2834), .B(w2837), .C(w2849), .D(w2827), .E(w2965) );
	vdp_nor4 g2929 (.Z(w2787), .A(COL[2]), .B(COL[3]), .C(COL[1]), .D(COL[0]) );
	vdp_nor g2930 (.Z(w2949), .A(w93), .B(w94) );
	vdp_nor g2931 (.Z(w2798), .A(w2967), .B(w2847) );
	vdp_nor g2932 (.Z(w2967), .A(w2698), .B(M5) );
	vdp_nand g2933 (.Z(w2799), .A(M5), .B(w2846) );
	vdp_nand g2934 (.Z(w2810), .A(SPR_PRIO), .B(w19) );
	vdp_and4 g2935 (.Z(w2824), .A(w2825), .B(w2955), .C(w2826), .D(w2830) );
	vdp_aoi21 g2936 (.Z(w2985), .B(w2713), .A2(w2983), .A1(w2760) );
	vdp_nor g2937 (.Z(w2857), .A(w21), .B(w20) );
	vdp_n_fet g2938 (.A(w2768), .Z(COL[6]) );
	vdp_slatch g2939 (.Q(w4128), .D(S[3]), .C(w3149), .nC(w3139) );
	vdp_slatch g2940 (.Q(w4130), .D(S[3]), .C(w3130), .nC(w3129) );
	vdp_slatch g2941 (.Q(w4132), .D(S[3]), .C(w3131), .nC(w3127) );
	vdp_slatch g2942 (.Q(w4134), .D(S[3]), .C(w3148), .nC(w3140) );
	vdp_slatch g2943 (.Q(w4136), .D(S[7]), .C(w3149), .nC(w3139) );
	vdp_slatch g2944 (.Q(w4139), .D(S[7]), .C(w3130), .nC(w3129) );
	vdp_slatch g2945 (.Q(w4138), .D(S[7]), .C(w3131), .nC(w3127) );
	vdp_slatch g2946 (.Q(w4143), .D(S[7]), .C(w3148), .nC(w3140) );
	vdp_slatch g2947 (.Q(w4142), .D(S[2]), .C(w3149), .nC(w3139) );
	vdp_slatch g2948 (.Q(w4149), .D(S[2]), .C(w3130), .nC(w3129) );
	vdp_slatch g2949 (.Q(w4148), .D(S[2]), .C(w3131), .nC(w3127) );
	vdp_slatch g2950 (.Q(w4151), .D(S[2]), .C(w3148), .nC(w3140) );
	vdp_slatch g2951 (.Q(w4150), .D(S[6]), .C(w3149), .nC(w3139) );
	vdp_slatch g2952 (.Q(w4155), .D(S[6]), .C(w3130), .nC(w3129) );
	vdp_slatch g2953 (.Q(w4154), .D(S[6]), .C(w3131), .nC(w3127) );
	vdp_slatch g2954 (.Q(w4159), .D(S[6]), .C(w3148), .nC(w3140) );
	vdp_slatch g2955 (.Q(w4158), .D(S[1]), .C(w3149), .nC(w3139) );
	vdp_slatch g2956 (.Q(w4163), .D(S[1]), .C(w3130), .nC(w3129) );
	vdp_slatch g2957 (.Q(w4162), .D(S[1]), .C(w3131), .nC(w3127) );
	vdp_slatch g2958 (.Q(w4167), .D(S[1]), .C(w3148), .nC(w3140) );
	vdp_slatch g2959 (.Q(w4166), .D(S[5]), .C(w3149), .nC(w3139) );
	vdp_slatch g2960 (.Q(w4171), .D(S[5]), .C(w3130), .nC(w3129) );
	vdp_slatch g2961 (.Q(w4170), .D(S[5]), .C(w3131), .nC(w3127) );
	vdp_slatch g2962 (.Q(w4175), .D(S[5]), .C(w3148), .nC(w3140) );
	vdp_slatch g2963 (.Q(w4174), .D(S[0]), .C(w3149), .nC(w3139) );
	vdp_slatch g2964 (.Q(w4179), .D(S[0]), .C(w3130), .nC(w3129) );
	vdp_slatch g2965 (.Q(w4178), .D(S[0]), .C(w3131), .nC(w3127) );
	vdp_slatch g2966 (.Q(w4183), .D(S[0]), .C(w3148), .nC(w3140) );
	vdp_slatch g2967 (.Q(w4182), .D(S[4]), .C(w3149), .nC(w3139) );
	vdp_slatch g2968 (.Q(w4187), .D(S[4]), .C(w3130), .nC(w3129) );
	vdp_slatch g2969 (.Q(w4186), .D(S[4]), .C(w3131), .nC(w3127) );
	vdp_slatch g2970 (.Q(w4190), .D(S[4]), .C(w3148), .nC(w3140) );
	vdp_slatch g2971 (.Q(w4129), .D(w4128), .C(w3119), .nC(w3136) );
	vdp_slatch g2972 (.Q(w4131), .D(w4130), .C(w3137), .nC(w3128) );
	vdp_slatch g2973 (.Q(w4133), .D(w4132), .C(w3138), .nC(w3126) );
	vdp_slatch g2974 (.Q(w4135), .D(w4134), .C(w3134), .nC(w3135) );
	vdp_slatch g2975 (.Q(w4137), .D(w4136), .C(w3119), .nC(w3136) );
	vdp_slatch g2976 (.Q(w4141), .D(w4139), .C(w3137), .nC(w3128) );
	vdp_slatch g2977 (.Q(w4140), .D(w4138), .C(w3138), .nC(w3126) );
	vdp_slatch g2978 (.Q(w4145), .D(w4143), .C(w3134), .nC(w3135) );
	vdp_slatch g2979 (.Q(w4144), .D(w4142), .C(w3119), .nC(w3136) );
	vdp_slatch g2980 (.Q(w4147), .D(w4149), .C(w3137), .nC(w3128) );
	vdp_slatch g2981 (.Q(w4146), .D(w4148), .C(w3138), .nC(w3126) );
	vdp_slatch g2982 (.Q(w4153), .D(w4151), .C(w3134), .nC(w3135) );
	vdp_slatch g2983 (.Q(w4152), .D(w4150), .C(w3119), .nC(w3136) );
	vdp_slatch g2984 (.Q(w4157), .D(w4155), .C(w3137), .nC(w3128) );
	vdp_slatch g2985 (.Q(w4156), .D(w4154), .C(w3138), .nC(w3126) );
	vdp_slatch g2986 (.Q(w4161), .D(w4159), .C(w3134), .nC(w3135) );
	vdp_slatch g2987 (.Q(w4160), .D(w4158), .C(w3119), .nC(w3136) );
	vdp_slatch g2988 (.Q(w4165), .D(w4163), .C(w3137), .nC(w3128) );
	vdp_slatch g2989 (.Q(w4164), .D(w4162), .C(w3138), .nC(w3126) );
	vdp_slatch g2990 (.Q(w4169), .D(w4167), .C(w3134), .nC(w3135) );
	vdp_slatch g2991 (.Q(w4168), .D(w4166), .C(w3119), .nC(w3136) );
	vdp_slatch g2992 (.Q(w4173), .D(w4171), .C(w3137), .nC(w3128) );
	vdp_slatch g2993 (.Q(w4172), .D(w4170), .C(w3138), .nC(w3126) );
	vdp_slatch g2994 (.Q(w4177), .D(w4175), .C(w3134), .nC(w3135) );
	vdp_slatch g2995 (.Q(w4176), .D(w4174), .C(w3119), .nC(w3136) );
	vdp_slatch g2996 (.Q(w4181), .D(w4179), .C(w3137), .nC(w3128) );
	vdp_slatch g2997 (.Q(w4180), .D(w4178), .C(w3138), .nC(w3126) );
	vdp_slatch g2998 (.Q(w4185), .D(w4183), .C(w3134), .nC(w3135) );
	vdp_slatch g2999 (.Q(w4184), .D(w4182), .C(w3119), .nC(w3136) );
	vdp_slatch g3000 (.Q(w4189), .D(w4187), .C(w3137), .nC(w3128) );
	vdp_slatch g3001 (.Q(w4188), .D(w4186), .C(w3138), .nC(w3126) );
	vdp_slatch g3002 (.Q(w4191), .D(w4190), .C(w3134), .nC(w3135) );
	vdp_slatch g3003 (.Q(w3176), .D(w4129), .C(w3141), .nC(w3167) );
	vdp_slatch g3004 (.Q(w3175), .D(w4131), .C(w3120), .nC(w3177) );
	vdp_slatch g3005 (.Q(w3174), .D(w4133), .C(w3132), .nC(w3178) );
	vdp_slatch g3006 (.Q(w3173), .D(w4135), .C(w3133), .nC(w3107) );
	vdp_slatch g3007 (.Q(w3172), .D(w4137), .C(w3141), .nC(w3167) );
	vdp_slatch g3008 (.Q(w3171), .D(w4141), .C(w3120), .nC(w3177) );
	vdp_slatch g3009 (.Q(w3170), .D(w4140), .C(w3132), .nC(w3178) );
	vdp_slatch g3010 (.Q(w3169), .D(w4145), .C(w3133), .nC(w3107) );
	vdp_slatch g3011 (.Q(w3168), .D(w4144), .C(w3141), .nC(w3167) );
	vdp_slatch g3012 (.Q(w3181), .D(w4147), .C(w3120), .nC(w3177) );
	vdp_slatch g3013 (.Q(w3185), .D(w4146), .C(w3132), .nC(w3178) );
	vdp_slatch g3014 (.Q(w3184), .D(w4153), .C(w3133), .nC(w3107) );
	vdp_slatch g3015 (.Q(w3183), .D(w4152), .C(w3141), .nC(w3167) );
	vdp_slatch g3016 (.Q(w3179), .D(w4157), .C(w3120), .nC(w3177) );
	vdp_slatch g3017 (.Q(w3180), .D(w4156), .C(w3132), .nC(w3178) );
	vdp_slatch g3018 (.D(w4161), .Q(w3182), .C(w3133), .nC(w3107) );
	vdp_slatch g3019 (.Q(w3186), .D(w4160), .C(w3141), .nC(w3167) );
	vdp_slatch g3020 (.Q(w3187), .D(w4165), .C(w3120), .nC(w3177) );
	vdp_slatch g3021 (.Q(w3189), .D(w4164), .C(w3132), .nC(w3178) );
	vdp_slatch g3022 (.Q(w3188), .D(w4169), .C(w3133), .nC(w3107) );
	vdp_slatch g3023 (.Q(w3230), .D(w4168), .C(w3141), .nC(w3167) );
	vdp_slatch g3024 (.Q(w3231), .D(w4173), .C(w3120), .nC(w3177) );
	vdp_slatch g3025 (.Q(w3227), .D(w4172), .C(w3132), .nC(w3178) );
	vdp_slatch g3026 (.Q(w3222), .D(w4177), .C(w3133), .nC(w3107) );
	vdp_slatch g3027 (.Q(w3234), .D(w4176), .C(w3141), .nC(w3167) );
	vdp_slatch g3028 (.Q(w3233), .D(w4181), .C(w3120), .nC(w3177) );
	vdp_slatch g3029 (.Q(w3232), .D(w4180), .C(w3132), .nC(w3178) );
	vdp_slatch g3030 (.Q(w3229), .D(w4185), .C(w3133), .nC(w3107) );
	vdp_slatch g3031 (.Q(w3215), .D(w4184), .C(w3141), .nC(w3167) );
	vdp_slatch g3032 (.Q(w3214), .D(w4189), .C(w3120), .nC(w3177) );
	vdp_slatch g3033 (.Q(w3216), .D(w4188), .C(w3132), .nC(w3178) );
	vdp_slatch g3034 (.Q(w3217), .D(w4191), .C(w3133), .nC(w3107) );
	vdp_slatch g3035 (.Q(w3294), .D(w4413), .C(w3290), .nC(w3292) );
	vdp_slatch g3036 (.Q(w3295), .D(w4414), .C(w3289), .nC(w3300) );
	vdp_slatch g3037 (.Q(w3296), .D(w4416), .C(w3288), .nC(w3301) );
	vdp_slatch g3038 (.Q(w3297), .D(w4415), .C(w3287), .nC(w3293) );
	vdp_slatch g3039 (.Q(w3298), .D(w4247), .C(w3290), .nC(w3292) );
	vdp_slatch g3040 (.Q(w3299), .D(w4246), .C(w3289), .nC(w3300) );
	vdp_slatch g3041 (.Q(w3305), .D(w4241), .C(w3288), .nC(w3301) );
	vdp_slatch g3042 (.Q(w3306), .D(w4240), .C(w3287), .nC(w3293) );
	vdp_slatch g3043 (.Q(w3307), .D(w4237), .C(w3290), .nC(w3292) );
	vdp_slatch g3044 (.Q(w3308), .D(w4236), .C(w3289), .nC(w3300) );
	vdp_slatch g3045 (.Q(w3309), .D(w4235), .C(w3288), .nC(w3301) );
	vdp_slatch g3046 (.Q(w3304), .D(w4232), .C(w3287), .nC(w3293) );
	vdp_slatch g3047 (.Q(w3310), .D(w4229), .C(w3290), .nC(w3292) );
	vdp_slatch g3048 (.Q(w3311), .D(w4230), .C(w3289), .nC(w3300) );
	vdp_slatch g3049 (.Q(w3312), .D(w4225), .C(w3288), .nC(w3301) );
	vdp_slatch g3050 (.Q(w3313), .D(w4226), .C(w3287), .nC(w3293) );
	vdp_slatch g3051 (.Q(w3238), .D(w4223), .C(w3290), .nC(w3292) );
	vdp_slatch g3052 (.Q(w4014), .D(w4222), .C(w3289), .nC(w3300) );
	vdp_slatch g3053 (.Q(w3240), .D(w4219), .C(w3288), .nC(w3301) );
	vdp_slatch g3054 (.Q(w3241), .D(w4218), .C(w3287), .nC(w3293) );
	vdp_slatch g3055 (.Q(w3314), .D(w4215), .C(w3290), .nC(w3292) );
	vdp_slatch g3056 (.Q(w3239), .D(w4214), .C(w3289), .nC(w3300) );
	vdp_slatch g3057 (.Q(w3219), .D(w4211), .C(w3288), .nC(w3301) );
	vdp_slatch g3058 (.Q(w3242), .D(w4210), .C(w3287), .nC(w3293) );
	vdp_slatch g3059 (.Q(w3245), .D(w4207), .C(w3290), .nC(w3292) );
	vdp_slatch g3060 (.Q(w3253), .D(w4206), .C(w3289), .nC(w3300) );
	vdp_slatch g3061 (.Q(w3252), .D(w4203), .C(w3288), .nC(w3301) );
	vdp_slatch g3062 (.Q(w3251), .D(w4202), .C(w3287), .nC(w3293) );
	vdp_slatch g3063 (.Q(w3249), .D(w4199), .C(w3290), .nC(w3292) );
	vdp_slatch g3064 (.Q(w3243), .D(w4198), .C(w3289), .nC(w3300) );
	vdp_slatch g3065 (.Q(w3250), .D(w4195), .C(w3288), .nC(w3301) );
	vdp_slatch g3066 (.Q(w3244), .D(w4194), .C(w3287), .nC(w3293) );
	vdp_slatch g3067 (.Q(w4413), .D(w4250), .C(w3291), .nC(w3278) );
	vdp_slatch g3068 (.Q(w4414), .D(w4251), .C(w3099), .nC(w3279) );
	vdp_slatch g3069 (.Q(w4416), .D(w4249), .C(w3285), .nC(w3087) );
	vdp_slatch g3070 (.Q(w4415), .D(w4248), .C(w3286), .nC(w3088) );
	vdp_slatch g3071 (.Q(w4247), .D(w4245), .C(w3291), .nC(w3278) );
	vdp_slatch g3072 (.Q(w4246), .D(w4244), .C(w3099), .nC(w3279) );
	vdp_slatch g3073 (.Q(w4241), .D(w4243), .C(w3285), .nC(w3087) );
	vdp_slatch g3074 (.Q(w4240), .D(w4242), .C(w3286), .nC(w3088) );
	vdp_slatch g3075 (.Q(w4237), .D(w4239), .C(w3291), .nC(w3278) );
	vdp_slatch g3076 (.Q(w4236), .D(w4238), .C(w3099), .nC(w3279) );
	vdp_slatch g3077 (.Q(w4235), .D(w4233), .C(w3285), .nC(w3087) );
	vdp_slatch g3078 (.Q(w4232), .D(w4234), .C(w3286), .nC(w3088) );
	vdp_slatch g3079 (.Q(w4229), .D(w4231), .C(w3291), .nC(w3278) );
	vdp_slatch g3080 (.Q(w4230), .D(w4228), .C(w3099), .nC(w3279) );
	vdp_slatch g3081 (.Q(w4225), .D(w4227), .C(w3285), .nC(w3087) );
	vdp_slatch g3082 (.Q(w4226), .D(w4224), .C(w3286), .nC(w3088) );
	vdp_slatch g3083 (.Q(w4223), .D(w4221), .C(w3291), .nC(w3278) );
	vdp_slatch g3084 (.Q(w4222), .D(w4220), .C(w3099), .nC(w3279) );
	vdp_slatch g3085 (.Q(w4219), .D(w4217), .C(w3285), .nC(w3087) );
	vdp_slatch g3086 (.Q(w4218), .D(w4216), .C(w3286), .nC(w3088) );
	vdp_slatch g3087 (.Q(w4215), .D(w4213), .C(w3291), .nC(w3278) );
	vdp_slatch g3088 (.Q(w4214), .D(w4212), .C(w3099), .nC(w3279) );
	vdp_slatch g3089 (.Q(w4211), .D(w4209), .C(w3285), .nC(w3087) );
	vdp_slatch g3090 (.Q(w4210), .D(w4208), .C(w3286), .nC(w3088) );
	vdp_slatch g3091 (.Q(w4207), .D(w4205), .C(w3291), .nC(w3278) );
	vdp_slatch g3092 (.Q(w4206), .D(w4204), .C(w3099), .nC(w3279) );
	vdp_slatch g3093 (.Q(w4203), .D(w4201), .C(w3285), .nC(w3087) );
	vdp_slatch g3094 (.Q(w4202), .D(w4200), .C(w3286), .nC(w3088) );
	vdp_slatch g3095 (.Q(w4199), .D(w4197), .C(w3291), .nC(w3278) );
	vdp_slatch g3096 (.Q(w4198), .D(w4196), .C(w3099), .nC(w3279) );
	vdp_slatch g3097 (.Q(w4195), .D(w4193), .C(w3285), .nC(w3087) );
	vdp_slatch g3098 (.Q(w4194), .D(w4192), .C(w3286), .nC(w3088) );
	vdp_slatch g3099 (.Q(w4250), .D(S[3]), .C(w3051), .nC(w3085) );
	vdp_slatch g3100 (.Q(w4251), .D(S[3]), .C(w3055), .nC(w3089) );
	vdp_slatch g3101 (.Q(w4249), .D(S[3]), .C(w3058), .nC(w3086) );
	vdp_slatch g3102 (.Q(w4248), .D(S[3]), .C(w3060), .nC(w3084) );
	vdp_slatch g3103 (.Q(w4245), .D(S[7]), .C(w3051), .nC(w3085) );
	vdp_slatch g3104 (.Q(w4244), .D(S[7]), .C(w3055), .nC(w3089) );
	vdp_slatch g3105 (.Q(w4243), .D(S[7]), .C(w3058), .nC(w3086) );
	vdp_slatch g3106 (.Q(w4242), .D(S[7]), .C(w3060), .nC(w3084) );
	vdp_slatch g3107 (.Q(w4239), .D(S[2]), .C(w3051), .nC(w3085) );
	vdp_slatch g3108 (.Q(w4238), .D(S[2]), .C(w3055), .nC(w3089) );
	vdp_slatch g3109 (.Q(w4233), .D(S[2]), .C(w3058), .nC(w3086) );
	vdp_slatch g3110 (.Q(w4234), .D(S[2]), .C(w3060), .nC(w3084) );
	vdp_slatch g3111 (.Q(w4231), .D(S[6]), .C(w3051), .nC(w3085) );
	vdp_slatch g3112 (.Q(w4228), .D(S[6]), .C(w3055), .nC(w3089) );
	vdp_slatch g3113 (.Q(w4227), .D(S[6]), .C(w3058), .nC(w3086) );
	vdp_slatch g3114 (.Q(w4224), .D(S[6]), .C(w3060), .nC(w3084) );
	vdp_slatch g3115 (.Q(w4221), .D(S[1]), .C(w3051), .nC(w3085) );
	vdp_slatch g3116 (.Q(w4220), .D(S[1]), .C(w3055), .nC(w3089) );
	vdp_slatch g3117 (.Q(w4217), .D(S[1]), .C(w3058), .nC(w3086) );
	vdp_slatch g3118 (.Q(w4216), .D(S[1]), .C(w3060), .nC(w3084) );
	vdp_slatch g3119 (.Q(w4213), .D(S[5]), .C(w3051), .nC(w3085) );
	vdp_slatch g3120 (.Q(w4212), .D(S[5]), .C(w3055), .nC(w3089) );
	vdp_slatch g3121 (.Q(w4209), .D(S[5]), .C(w3058), .nC(w3086) );
	vdp_slatch g3122 (.Q(w4208), .D(S[5]), .C(w3060), .nC(w3084) );
	vdp_slatch g3123 (.Q(w4205), .D(S[0]), .C(w3051), .nC(w3085) );
	vdp_slatch g3124 (.Q(w4204), .D(S[0]), .C(w3055), .nC(w3089) );
	vdp_slatch g3125 (.Q(w4201), .D(S[0]), .C(w3058), .nC(w3086) );
	vdp_slatch g3126 (.Q(w4200), .D(S[0]), .C(w3060), .nC(w3084) );
	vdp_slatch g3127 (.Q(w4197), .D(S[4]), .C(w3051), .nC(w3085) );
	vdp_slatch g3128 (.Q(w4196), .D(S[4]), .C(w3055), .nC(w3089) );
	vdp_slatch g3129 (.Q(w4193), .D(S[4]), .C(w3058), .nC(w3086) );
	vdp_slatch g3130 (.Q(w4192), .D(S[4]), .C(w3060), .nC(w3084) );
	vdp_slatch g3131 (.Q(w4255), .D(S[3]), .C(w3052), .nC(w3077) );
	vdp_slatch g3132 (.Q(w4254), .D(S[3]), .C(w3056), .nC(w3082) );
	vdp_slatch g3133 (.Q(w4259), .D(S[3]), .C(w3057), .nC(w3083) );
	vdp_slatch g3134 (.Q(w4258), .D(S[3]), .C(w3059), .nC(w3078) );
	vdp_slatch g3135 (.Q(w4263), .D(S[7]), .C(w3052), .nC(w3077) );
	vdp_slatch g3136 (.Q(w4262), .D(S[7]), .C(w3056), .nC(w3082) );
	vdp_slatch g3137 (.Q(w4267), .D(S[7]), .C(w3057), .nC(w3083) );
	vdp_slatch g3138 (.Q(w4266), .D(S[7]), .C(w3059), .nC(w3078) );
	vdp_slatch g3139 (.Q(w4271), .D(S[2]), .C(w3052), .nC(w3077) );
	vdp_slatch g3140 (.Q(w4270), .D(S[2]), .C(w3056), .nC(w3082) );
	vdp_slatch g3141 (.Q(w4275), .D(S[2]), .C(w3057), .nC(w3083) );
	vdp_slatch g3142 (.Q(w4274), .D(S[2]), .C(w3059), .nC(w3078) );
	vdp_slatch g3143 (.Q(w4277), .D(S[6]), .C(w3052), .nC(w3077) );
	vdp_slatch g3144 (.Q(w4278), .D(S[6]), .C(w3056), .nC(w3082) );
	vdp_slatch g3145 (.Q(w4314), .D(S[6]), .C(w3057), .nC(w3083) );
	vdp_slatch g3146 (.Q(w4313), .D(S[6]), .C(w3059), .nC(w3078) );
	vdp_slatch g3147 (.Q(w4310), .D(S[1]), .C(w3052), .nC(w3077) );
	vdp_slatch g3148 (.Q(w4309), .D(S[1]), .C(w3056), .nC(w3082) );
	vdp_slatch g3149 (.Q(w4306), .D(S[1]), .C(w3057), .nC(w3083) );
	vdp_slatch g3150 (.Q(w4305), .D(S[1]), .C(w3059), .nC(w3078) );
	vdp_slatch g3151 (.Q(w4302), .D(S[5]), .C(w3052), .nC(w3077) );
	vdp_slatch g3152 (.Q(w4301), .D(S[5]), .C(w3056), .nC(w3082) );
	vdp_slatch g3153 (.Q(w4298), .D(S[5]), .C(w3057), .nC(w3083) );
	vdp_slatch g3154 (.Q(w4297), .D(S[5]), .C(w3059), .nC(w3078) );
	vdp_slatch g3155 (.Q(w4294), .D(S[0]), .C(w3052), .nC(w3077) );
	vdp_slatch g3156 (.Q(w4293), .D(S[0]), .C(w3056), .nC(w3082) );
	vdp_slatch g3157 (.Q(w4290), .D(S[0]), .C(w3057), .nC(w3083) );
	vdp_slatch g3158 (.Q(w4289), .D(S[0]), .C(w3059), .nC(w3078) );
	vdp_slatch g3159 (.Q(w4286), .D(S[4]), .C(w3052), .nC(w3077) );
	vdp_slatch g3160 (.Q(w4285), .D(S[4]), .C(w3056), .nC(w3082) );
	vdp_slatch g3161 (.Q(w4282), .D(S[4]), .C(w3057), .nC(w3083) );
	vdp_slatch g3162 (.Q(w4281), .D(S[4]), .C(w3059), .nC(w3078) );
	vdp_slatch g3163 (.Q(w4253), .D(w4255), .C(w3039), .nC(w3079) );
	vdp_slatch g3164 (.Q(w4252), .D(w4254), .C(w3042), .nC(w3080) );
	vdp_slatch g3165 (.Q(w4257), .D(w4259), .C(w3047), .nC(w3081) );
	vdp_slatch g3166 (.Q(w4256), .D(w4258), .C(w3044), .nC(w3049) );
	vdp_slatch g3167 (.Q(w4261), .D(w4263), .C(w3039), .nC(w3079) );
	vdp_slatch g3168 (.Q(w4260), .D(w4262), .C(w3042), .nC(w3080) );
	vdp_slatch g3169 (.Q(w4265), .D(w4267), .C(w3047), .nC(w3081) );
	vdp_slatch g3170 (.Q(w4264), .D(w4266), .C(w3044), .nC(w3049) );
	vdp_slatch g3171 (.Q(w4269), .D(w4271), .C(w3039), .nC(w3079) );
	vdp_slatch g3172 (.Q(w4268), .D(w4270), .C(w3042), .nC(w3080) );
	vdp_slatch g3173 (.Q(w4379), .D(w4275), .C(w3047), .nC(w3081) );
	vdp_slatch g3174 (.Q(w4273), .D(w4274), .C(w3044), .nC(w3049) );
	vdp_slatch g3175 (.Q(w4272), .D(w4277), .C(w3039), .nC(w3079) );
	vdp_slatch g3176 (.Q(w4276), .D(w4278), .C(w3042), .nC(w3080) );
	vdp_slatch g3177 (.Q(w4312), .D(w4314), .C(w3047), .nC(w3081) );
	vdp_slatch g3178 (.Q(w4311), .D(w4313), .C(w3044), .nC(w3049) );
	vdp_slatch g3179 (.Q(w4308), .D(w4310), .C(w3039), .nC(w3079) );
	vdp_slatch g3180 (.Q(w4307), .D(w4309), .C(w3042), .nC(w3080) );
	vdp_slatch g3181 (.Q(w4304), .D(w4306), .C(w3047), .nC(w3081) );
	vdp_slatch g3182 (.Q(w4303), .D(w4305), .C(w3044), .nC(w3049) );
	vdp_slatch g3183 (.Q(w4300), .D(w4302), .C(w3039), .nC(w3079) );
	vdp_slatch g3184 (.Q(w4299), .D(w4301), .C(w3042), .nC(w3080) );
	vdp_slatch g3185 (.Q(w4296), .D(w4298), .C(w3047), .nC(w3081) );
	vdp_slatch g3186 (.Q(w4295), .D(w4297), .C(w3044), .nC(w3049) );
	vdp_slatch g3187 (.D(w4294), .Q(w4292), .C(w3039), .nC(w3079) );
	vdp_slatch g3188 (.Q(w4291), .D(w4293), .C(w3042), .nC(w3080) );
	vdp_slatch g3189 (.Q(w4288), .D(w4290), .C(w3047), .nC(w3081) );
	vdp_slatch g3190 (.Q(w4287), .D(w4289), .C(w3044), .nC(w3049) );
	vdp_slatch g3191 (.Q(w4284), .D(w4286), .C(w3039), .nC(w3079) );
	vdp_slatch g3192 (.Q(w4283), .D(w4285), .C(w3042), .nC(w3080) );
	vdp_slatch g3193 (.Q(w4280), .D(w4282), .C(w3047), .nC(w3081) );
	vdp_slatch g3194 (.Q(w4279), .D(w4281), .C(w3044), .nC(w3049) );
	vdp_slatch g3195 (.Q(w3360), .D(w4253), .C(w3040), .nC(w3041) );
	vdp_slatch g3196 (.Q(w3359), .D(w4252), .C(w3048), .nC(w3043) );
	vdp_slatch g3197 (.Q(w3347), .D(w4257), .C(w3045), .nC(w3046) );
	vdp_slatch g3198 (.Q(w3345), .D(w4256), .C(w3038), .nC(w3037) );
	vdp_slatch g3199 (.Q(w3358), .D(w4261), .C(w3040), .nC(w3041) );
	vdp_slatch g3200 (.Q(w3357), .D(w4260), .C(w3048), .nC(w3043) );
	vdp_slatch g3201 (.D(w4265), .C(w3045), .nC(w3046), .Q(w3356) );
	vdp_slatch g3202 (.Q(w3344), .D(w4264), .C(w3038), .nC(w3037) );
	vdp_slatch g3203 (.Q(w3355), .D(w4269), .C(w3040), .nC(w3041) );
	vdp_slatch g3204 (.Q(w3354), .D(w4268), .C(w3048), .nC(w3043) );
	vdp_slatch g3205 (.Q(w3353), .D(w4379), .C(w3045), .nC(w3046) );
	vdp_slatch g3206 (.Q(w3352), .D(w4273), .C(w3038), .nC(w3037) );
	vdp_slatch g3207 (.Q(w3351), .D(w4272), .C(w3040), .nC(w3041) );
	vdp_slatch g3208 (.Q(w3350), .D(w4276), .C(w3048), .nC(w3043) );
	vdp_slatch g3209 (.Q(w3349), .D(w4312), .C(w3045), .nC(w3046) );
	vdp_slatch g3210 (.Q(w3348), .D(w4311), .C(w3038), .nC(w3037) );
	vdp_slatch g3211 (.Q(w3340), .D(w4308), .C(w3040), .nC(w3041) );
	vdp_slatch g3212 (.Q(w3386), .D(w4307), .C(w3048), .nC(w3043) );
	vdp_slatch g3213 (.Q(w3341), .D(w4304), .C(w3045), .nC(w3046) );
	vdp_slatch g3214 (.Q(w3342), .D(w4303), .C(w3038), .nC(w3037) );
	vdp_slatch g3215 (.Q(w3390), .D(w4300), .C(w3040), .nC(w3041) );
	vdp_slatch g3216 (.Q(w3399), .D(w4299), .C(w3048), .nC(w3043) );
	vdp_slatch g3217 (.Q(w3391), .D(w4296), .C(w3045), .nC(w3046) );
	vdp_slatch g3218 (.Q(w3398), .D(w4295), .nC(w3037), .C(w3038) );
	vdp_slatch g3219 (.Q(w3397), .D(w4292), .C(w3040), .nC(w3041) );
	vdp_slatch g3220 (.Q(w3396), .D(w4291), .C(w3048), .nC(w3043) );
	vdp_slatch g3221 (.Q(w3392), .D(w4288), .C(w3045), .nC(w3046) );
	vdp_slatch g3222 (.Q(w3395), .D(w4287), .C(w3038), .nC(w3037) );
	vdp_slatch g3223 (.Q(w3394), .D(w4284), .C(w3040), .nC(w3041) );
	vdp_slatch g3224 (.Q(w3393), .D(w4283), .C(w3048), .nC(w3043) );
	vdp_slatch g3225 (.Q(w3346), .D(w4280), .C(w3045), .nC(w3046) );
	vdp_slatch g3226 (.Q(w3343), .D(w4279), .C(w3038), .nC(w3037) );
	vdp_slatch g3227 (.Q(w3378), .D(w4318), .nC(w3440), .C(w3439) );
	vdp_slatch g3228 (.Q(w3487), .D(w4317), .nC(w3443), .C(w3444) );
	vdp_slatch g3229 (.Q(w3380), .D(w4322), .nC(w3442), .C(w3441) );
	vdp_slatch g3230 (.Q(w3379), .D(w4321), .nC(w3446), .C(w3445) );
	vdp_slatch g3231 (.Q(w3486), .D(w4326), .nC(w3440), .C(w3439) );
	vdp_slatch g3232 (.Q(w3490), .D(w4325), .nC(w3443), .C(w3444) );
	vdp_slatch g3233 (.Q(w3489), .D(w4330), .nC(w3442), .C(w3441) );
	vdp_slatch g3234 (.Q(w3488), .D(w4329), .nC(w3446), .C(w3445) );
	vdp_slatch g3235 (.Q(w3381), .D(w4334), .nC(w3440), .C(w3439) );
	vdp_slatch g3236 (.Q(w3491), .D(w4333), .nC(w3443), .C(w3444) );
	vdp_slatch g3237 (.Q(w3485), .D(w4338), .nC(w3442), .C(w3441) );
	vdp_slatch g3238 (.Q(w3492), .D(w4337), .nC(w3446), .C(w3445) );
	vdp_slatch g3239 (.Q(w3493), .D(w4342), .nC(w3440), .C(w3439) );
	vdp_slatch g3240 (.Q(w3494), .D(w4341), .nC(w3443), .C(w3444) );
	vdp_slatch g3241 (.Q(w3382), .D(w4346), .nC(w3442), .C(w3441) );
	vdp_slatch g3242 (.Q(w3383), .D(w4345), .nC(w3446), .C(w3445) );
	vdp_slatch g3243 (.Q(w3477), .D(w4350), .nC(w3440), .C(w3439) );
	vdp_slatch g3244 (.Q(w3478), .D(w4349), .nC(w3443), .C(w3444) );
	vdp_slatch g3245 (.Q(w3479), .D(w4354), .nC(w3442), .C(w3441) );
	vdp_slatch g3246 (.Q(w3480), .D(w4353), .nC(w3446), .C(w3445) );
	vdp_slatch g3247 (.Q(w3481), .D(w4358), .nC(w3440), .C(w3439) );
	vdp_slatch g3248 (.Q(w3482), .D(w4357), .nC(w3443), .C(w3444) );
	vdp_slatch g3249 (.Q(w3483), .D(w4362), .nC(w3442), .C(w3441) );
	vdp_slatch g3250 (.Q(w3484), .D(w4361), .nC(w3446), .C(w3445) );
	vdp_slatch g3251 (.Q(w3476), .D(w4366), .nC(w3440), .C(w3439) );
	vdp_slatch g3252 (.Q(w3475), .D(w4365), .nC(w3443), .C(w3444) );
	vdp_slatch g3253 (.Q(w3474), .D(w4370), .nC(w3442), .C(w3441) );
	vdp_slatch g3254 (.Q(w3473), .D(w4369), .nC(w3446), .C(w3445) );
	vdp_slatch g3255 (.Q(w3472), .D(w4374), .nC(w3440), .C(w3439) );
	vdp_slatch g3256 (.Q(w3471), .D(w4373), .nC(w3443), .C(w3444) );
	vdp_slatch g3257 (.Q(w3469), .D(w4378), .nC(w3442), .C(w3441) );
	vdp_slatch g3258 (.Q(w3470), .D(w4377), .nC(w3446), .C(w3445) );
	vdp_slatch g3259 (.Q(w4318), .D(w4316), .C(w3404), .nC(w3438) );
	vdp_slatch g3260 (.Q(w4317), .D(w4315), .C(w3430), .nC(w3432) );
	vdp_slatch g3261 (.Q(w4322), .D(w4320), .C(w3405), .nC(w3433) );
	vdp_slatch g3262 (.Q(w4321), .D(w4319), .C(w3437), .nC(w3436) );
	vdp_slatch g3263 (.Q(w4326), .D(w4324), .C(w3404), .nC(w3438) );
	vdp_slatch g3264 (.Q(w4325), .D(w4323), .C(w3430), .nC(w3432) );
	vdp_slatch g3265 (.Q(w4330), .D(w4328), .C(w3405), .nC(w3433) );
	vdp_slatch g3266 (.Q(w4329), .D(w4327), .C(w3437), .nC(w3436) );
	vdp_slatch g3267 (.Q(w4334), .D(w4332), .C(w3404), .nC(w3438) );
	vdp_slatch g3268 (.Q(w4333), .D(w4331), .C(w3430), .nC(w3432) );
	vdp_slatch g3269 (.Q(w4338), .D(w4336), .C(w3405), .nC(w3433) );
	vdp_slatch g3270 (.Q(w4337), .D(w4335), .C(w3437), .nC(w3436) );
	vdp_slatch g3271 (.Q(w4342), .D(w4340), .C(w3404), .nC(w3438) );
	vdp_slatch g3272 (.Q(w4341), .D(w4339), .C(w3430), .nC(w3432) );
	vdp_slatch g3273 (.Q(w4346), .D(w4344), .C(w3405), .nC(w3433) );
	vdp_slatch g3274 (.Q(w4345), .D(w4343), .C(w3437), .nC(w3436) );
	vdp_slatch g3275 (.Q(w4350), .D(w4348), .C(w3404), .nC(w3438) );
	vdp_slatch g3276 (.Q(w4349), .D(w4347), .C(w3430), .nC(w3432) );
	vdp_slatch g3277 (.Q(w4354), .D(w4352), .C(w3405), .nC(w3433) );
	vdp_slatch g3278 (.Q(w4353), .D(w4351), .C(w3437), .nC(w3436) );
	vdp_slatch g3279 (.Q(w4358), .D(w4356), .C(w3404), .nC(w3438) );
	vdp_slatch g3280 (.Q(w4357), .D(w4355), .C(w3430), .nC(w3432) );
	vdp_slatch g3281 (.Q(w4362), .D(w4360), .C(w3405), .nC(w3433) );
	vdp_slatch g3282 (.Q(w4361), .D(w4359), .C(w3437), .nC(w3436) );
	vdp_slatch g3283 (.Q(w4366), .D(w4364), .C(w3404), .nC(w3438) );
	vdp_slatch g3284 (.Q(w4365), .D(w4363), .C(w3430), .nC(w3432) );
	vdp_slatch g3285 (.Q(w4370), .D(w4368), .C(w3405), .nC(w3433) );
	vdp_slatch g3286 (.Q(w4369), .D(w4367), .C(w3437), .nC(w3436) );
	vdp_slatch g3287 (.Q(w4374), .D(w4372), .C(w3404), .nC(w3438) );
	vdp_slatch g3288 (.Q(w4373), .D(w4371), .C(w3430), .nC(w3432) );
	vdp_slatch g3289 (.Q(w4378), .D(w4376), .C(w3405), .nC(w3433) );
	vdp_slatch g3290 (.Q(w4377), .D(w4375), .C(w3437), .nC(w3436) );
	vdp_slatch g3291 (.Q(w4316), .D(S[3]), .nC(w3431), .C(w3459) );
	vdp_slatch g3292 (.Q(w4315), .D(S[3]), .nC(w3447), .C(w3460) );
	vdp_slatch g3293 (.Q(w4320), .D(S[3]), .nC(w3434), .C(w3458) );
	vdp_slatch g3294 (.Q(w4319), .D(S[3]), .nC(w3435), .C(w3457) );
	vdp_slatch g3295 (.Q(w4324), .D(S[7]), .nC(w3431), .C(w3459) );
	vdp_slatch g3296 (.Q(w4323), .D(S[7]), .nC(w3447), .C(w3460) );
	vdp_slatch g3297 (.Q(w4328), .D(S[7]), .nC(w3434), .C(w3458) );
	vdp_slatch g3298 (.Q(w4327), .D(S[7]), .nC(w3435), .C(w3457) );
	vdp_slatch g3299 (.Q(w4332), .D(S[2]), .nC(w3431), .C(w3459) );
	vdp_slatch g3300 (.Q(w4331), .D(S[2]), .nC(w3447), .C(w3460) );
	vdp_slatch g3301 (.Q(w4336), .D(S[2]), .nC(w3434), .C(w3458) );
	vdp_slatch g3302 (.Q(w4335), .D(S[2]), .nC(w3435), .C(w3457) );
	vdp_slatch g3303 (.Q(w4340), .D(S[6]), .nC(w3431), .C(w3459) );
	vdp_slatch g3304 (.Q(w4339), .D(S[6]), .nC(w3447), .C(w3460) );
	vdp_slatch g3305 (.Q(w4344), .D(S[6]), .nC(w3434), .C(w3458) );
	vdp_slatch g3306 (.Q(w4343), .D(S[6]), .nC(w3435), .C(w3457) );
	vdp_slatch g3307 (.Q(w4348), .D(S[1]), .nC(w3431), .C(w3459) );
	vdp_slatch g3308 (.Q(w4347), .D(S[1]), .nC(w3447), .C(w3460) );
	vdp_slatch g3309 (.Q(w4352), .D(S[1]), .nC(w3434), .C(w3458) );
	vdp_slatch g3310 (.Q(w4351), .D(S[1]), .nC(w3435), .C(w3457) );
	vdp_slatch g3311 (.Q(w4356), .D(S[5]), .nC(w3431), .C(w3459) );
	vdp_slatch g3312 (.Q(w4355), .D(S[5]), .nC(w3447), .C(w3460) );
	vdp_slatch g3313 (.Q(w4360), .D(S[5]), .nC(w3434), .C(w3458) );
	vdp_slatch g3314 (.Q(w4359), .D(S[5]), .nC(w3435), .C(w3457) );
	vdp_slatch g3315 (.Q(w4364), .D(S[0]), .nC(w3431), .C(w3459) );
	vdp_slatch g3316 (.Q(w4363), .D(S[0]), .nC(w3447), .C(w3460) );
	vdp_slatch g3317 (.Q(w4368), .D(S[0]), .nC(w3434), .C(w3458) );
	vdp_slatch g3318 (.Q(w4367), .D(S[0]), .nC(w3435), .C(w3457) );
	vdp_slatch g3319 (.Q(w4372), .D(S[4]), .nC(w3431), .C(w3459) );
	vdp_slatch g3320 (.Q(w4371), .D(S[4]), .nC(w3447), .C(w3460) );
	vdp_slatch g3321 (.Q(w4376), .D(S[4]), .nC(w3434), .C(w3458) );
	vdp_slatch g3322 (.Q(w4375), .D(S[4]), .nC(w3435), .C(w3457) );
	vdp_aon2x8 g3323 (.Z(w4013), .A1(w3176), .B1(w3175), .C1(w3174), .D2(w3173), .A2(w3220), .B2(w3221), .C2(w3226), .D1(w3225), .E2(w3223), .F1(w3224), .E1(w3172), .F2(w3171), .G1(w3170), .H2(w3169), .G2(w3228), .H1(w3218) );
	vdp_aon2x8 g3324 (.Z(w3200), .A1(w3294), .B1(w3221), .C1(w3296), .D2(w3225), .A2(w3220), .B2(w3295), .C2(w3226), .D1(w3297), .E2(w3223), .F1(w3224), .E1(w3298), .F2(w3299), .G1(w3305), .H2(w3306), .G2(w3228), .H1(w3218) );
	vdp_aon2x8 g3325 (.Z(w3203), .A1(w3168), .B1(w3181), .C1(w3185), .D2(w3184), .A2(w3220), .B2(w3221), .C2(w3226), .D1(w3225), .E2(w3223), .F1(w3224), .E1(w3183), .F2(w3179), .G1(w3180), .H2(w3182), .G2(w3228), .H1(w3218) );
	vdp_aon2x8 g3326 (.Z(w3204), .A1(w3307), .B1(w3221), .C1(w3309), .D2(w3225), .A2(w3220), .B2(w3308), .C2(w3226), .D1(w3304), .E2(w3223), .F1(w3224), .E1(w3310), .F2(w3311), .G1(w3312), .H2(w3313), .G2(w3228), .H1(w3218) );
	vdp_aon2x8 g3327 (.Z(w3202), .A1(w3238), .B1(w3221), .C1(w3240), .D2(w3241), .A2(w3220), .B2(w4014), .C2(w3226), .D1(w3225), .E2(w3223), .F1(w3224), .E1(w3314), .F2(w3239), .G1(w3219), .H2(w3242), .G2(w3228), .H1(w3218) );
	vdp_aon2x8 g3328 (.Z(w3205), .A1(w3245), .B1(w3221), .C1(w3252), .D2(w3251), .A2(w3220), .B2(w3253), .C2(w3226), .D1(w3225), .E2(w3223), .F1(w3224), .E1(w3249), .F2(w3243), .G1(w3250), .G2(w3228), .H1(w3218), .H2(w3244) );
	vdp_aon2x8 g3329 (.Z(w3201), .A1(w3186), .B1(w3187), .C1(w3189), .D2(w3188), .A2(w3220), .B2(w3221), .C2(w3226), .D1(w3225), .E2(w3223), .F1(w3224), .E1(w3230), .F2(w3231), .G1(w3227), .H2(w3222), .G2(w3228), .H1(w3218) );
	vdp_aon2x8 g3330 (.Z(w3206), .A1(w3234), .B1(w3233), .C1(w3232), .D2(w3229), .A2(w3220), .B2(w3221), .C2(w3226), .D1(w3225), .E2(w3223), .F1(w3224), .E1(w3215), .F2(w3214), .G1(w3216), .H2(w3217), .G2(w3228), .H1(w3218) );
	vdp_aon2x8 g3331 (.A1(w3360), .B1(w3359), .C1(w3347), .D2(w3345), .A2(w3377), .B2(w3376), .C2(w3375), .D1(w3374), .E2(w3373), .F1(w3372), .E1(w3358), .F2(w3357), .G1(w3356), .H2(w3344), .G2(w3370), .H1(w3371), .Z(w3389) );
	vdp_aon2x8 g3332 (.Z(w3417), .A1(w3355), .B1(w3354), .C1(w3353), .D2(w3352), .A2(w3377), .B2(w3376), .C2(w3375), .D1(w3374), .E2(w3373), .F1(w3372), .E1(w3351), .F2(w3350), .G1(w3349), .H2(w3348), .G2(w3370), .H1(w3371) );
	vdp_aon2x8 g3333 (.Z(w3388), .A1(w3347), .B1(w3356), .C1(w3353), .D2(w3349), .A2(w3372), .B2(w3371), .C2(w3376), .D1(w3374), .E2(w3373), .F1(w3370), .E1(w3341), .F2(w3391), .G1(w3392), .H2(w3346), .G2(w3377), .H1(w3375) );
	vdp_aon2x8 g3334 (.Z(w3420), .A1(w3340), .B1(w3386), .C1(w3341), .D2(w3342), .A2(w3377), .B2(w3376), .C2(w3375), .D1(w3374), .E2(w3373), .F1(w3372), .E1(w3390), .F2(w3399), .G1(w3391), .H2(w3398), .G2(w3370), .H1(w3371) );
	vdp_aon2x8 g3335 (.Z(w3387), .A1(w3397), .B1(w3396), .C1(w3392), .D2(w3395), .A2(w3377), .B2(w3376), .C2(w3375), .D1(w3374), .E2(w3373), .F1(w3372), .E1(w3394), .F2(w3393), .G1(w3346), .H2(w3343), .G2(w3370), .H1(w3371) );
	vdp_aon2x8 g3336 (.Z(w3422), .A1(w3476), .B1(w3376), .C1(w3474), .D2(w3374), .A2(w3377), .B2(w3475), .C2(w3375), .D1(w3473), .E2(w3373), .F1(w3372), .E1(w3472), .F2(w3471), .G1(w3469), .H2(w3470), .G2(w3370), .H1(w3371) );
	vdp_aon2x8 g3337 (.Z(w3423), .A1(w3477), .B1(w3376), .C1(w3479), .D2(w3374), .A2(w3377), .B2(w3478), .C2(w3375), .D1(w3480), .E2(w3373), .F1(w3372), .E1(w3481), .F2(w3482), .G1(w3483), .H2(w3484), .G2(w3370), .H1(w3371) );
	vdp_aon2x8 g3338 (.Z(w3421), .A1(w3345), .B1(w3344), .C1(w3352), .D2(w3348), .A2(w3372), .B2(w3371), .C2(w3376), .D1(w3374), .E2(w3373), .F1(w3370), .E1(w3342), .F2(w3398), .G1(w3395), .H2(w3343), .G2(w3377), .H1(w3375) );
	vdp_aon2x8 g3339 (.Z(w3416), .A1(w3379), .B1(w3371), .C1(w3492), .D2(w3374), .A2(w3372), .B2(w3488), .C2(w3376), .D1(w3383), .E2(w3373), .F1(w3370), .E1(w3480), .F2(w3484), .G1(w3473), .H2(w3470), .G2(w3377), .H1(w3375) );
	vdp_aon2x8 g3340 (.Z(w3419), .A1(w3380), .B1(w3371), .C1(w3485), .D2(w3374), .A2(w3372), .B2(w3489), .C2(w3376), .D1(w3382), .E2(w3373), .F1(w3370), .E1(w3479), .F2(w3483), .G1(w3474), .H2(w3469), .G2(w3377), .H1(w3375) );
	vdp_aon2x8 g3341 (.Z(w3418), .A1(w3381), .B1(w3376), .C1(w3485), .D2(w3374), .A2(w3377), .B2(w3491), .C2(w3375), .D1(w3492), .E2(w3373), .F1(w3372), .E1(w3493), .F2(w3494), .G1(w3382), .H2(w3383), .G2(w3370), .H1(w3371) );
	vdp_aon2x8 g3342 (.A1(w3378), .B1(w3376), .C1(w3380), .D2(w3374), .A2(w3377), .B2(w3487), .C2(w3375), .D1(w3379), .E2(w3373), .F1(w3372), .E1(w3486), .F2(w3490), .G1(w3489), .H2(w3488), .G2(w3370), .H1(w3371), .Z(w3424) );
	vdp_sr_bit g3343 (.Q(w3367), .D(w3522), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3344 (.Q(w3522), .D(w3426), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3345 (.Q(w3427), .D(w3523), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3346 (.Q(w3523), .D(w3429), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3347 (.Q(w3428), .D(w3403), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3348 (.Q(w4044), .D(w3428), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3349 (.Q(w3507), .D(w3425), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3350 (.Q(w3402), .D(w3507), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3351 (.Q(w4046), .D(w3412), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3352 (.Q(w3401), .D(w4046), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3353 (.Q(w3400), .D(w3368), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3354 (.Q(w3368), .D(w3411), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3355 (.Q(w2816), .D(w3413), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3356 (.Q(w3508), .D(w2816), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3357 (.Q(w3192), .D(w3210), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3358 (.Q(w3194), .D(w3192), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3359 (.Q(w3197), .D(w3193), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3360 (.Q(w3193), .D(w3209), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3361 (.Q(w3208), .D(w3190), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3362 (.Q(w3190), .D(w3211), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3363 (.Q(w3191), .D(w3207), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3364 (.Q(w3199), .D(w3191), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3365 (.Q(w3277), .D(w2815), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3366 (.Q(w2815), .D(w3262), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3367 (.Q(w4025), .D(w3212), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3368 (.Q(w3198), .D(w4025), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3369 (.Q(w4024), .D(w3263), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3370 (.Q(w3196), .D(w4024), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3371 (.Q(w3124), .D(VRAMA[1]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3372 (.Q(w3156), .D(VRAMA[2]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3373 (.Q(w3158), .D(VRAMA[3]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3374 (.Q(w3159), .D(VRAMA[4]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3375 (.Q(w3160), .D(VRAMA[5]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3376 (.Q(w3161), .D(VRAMA[6]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3377 (.Q(w4022), .D(w3147), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3378 (.Q(w3509), .D(w4022), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3379 (.Q(w3146), .D(w3510), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3380 (.Q(w3510), .D(w3509), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_dlatch_inv g3381 (.nQ(w3147), .D(w3112), .C(DCLK1), .nC(nDCLK1) );
	vdp_slatch g3382 (.Q(w3271), .D(w4380), .C(w3264), .nC(w3025) );
	vdp_slatch g3383 (.Q(w3270), .D(w4381), .C(w3264), .nC(w3025) );
	vdp_slatch g3384 (.Q(w3269), .D(w4382), .C(w3264), .nC(w3025) );
	vdp_slatch g3385 (.Q(w3268), .D(w4383), .C(w3264), .nC(w3025) );
	vdp_slatch g3386 (.Q(w3267), .D(w4384), .C(w3264), .nC(w3025) );
	vdp_slatch g3387 (.Q(w3266), .D(w4385), .C(w3264), .nC(w3025) );
	vdp_slatch g3388 (.Q(w3265), .D(w4387), .C(w3264), .nC(w3025) );
	vdp_slatch g3389 (.Q(w3026), .D(w4386), .C(w3264), .nC(w3025) );
	vdp_slatch g3390 (.Q(w4380), .D(w3093), .C(w3284), .nC(w3316) );
	vdp_slatch g3391 (.Q(w4381), .D(w3067), .C(w3284), .nC(w3316) );
	vdp_slatch g3392 (.Q(w4382), .D(w3069), .C(w3284), .nC(w3316) );
	vdp_slatch g3393 (.Q(w4383), .D(w3070), .C(w3284), .nC(w3316) );
	vdp_slatch g3394 (.Q(w4384), .D(w3071), .C(w3284), .nC(w3316) );
	vdp_slatch g3395 (.Q(w4385), .D(w3094), .C(w3284), .nC(w3316) );
	vdp_slatch g3396 (.Q(w4387), .D(w3098), .C(w3284), .nC(w3316) );
	vdp_slatch g3397 (.Q(w4386), .D(w3097), .C(w3284), .nC(w3316) );
	vdp_slatch g3398 (.Q(w4388), .D(w3033), .C(w3035), .nC(w3034) );
	vdp_slatch g3399 (.Q(w4389), .D(w3066), .C(w3035), .nC(w3034) );
	vdp_slatch g3400 (.Q(w4390), .D(w3032), .C(w3035), .nC(w3034) );
	vdp_slatch g3401 (.Q(w4391), .D(w4077), .C(w3035), .nC(w3034) );
	vdp_slatch g3402 (.Q(w4392), .D(w3518), .C(w3035), .nC(w3034) );
	vdp_slatch g3403 (.Q(w4393), .D(w3073), .C(w3035), .nC(w3034) );
	vdp_slatch g3404 (.Q(w4394), .D(w3029), .C(w3035), .nC(w3034) );
	vdp_slatch g3405 (.Q(w4395), .D(w3074), .C(w3035), .nC(w3034) );
	vdp_slatch g3406 (.Q(w3325), .D(w4388), .C(w3036), .nC(w3318) );
	vdp_slatch g3407 (.Q(w3324), .D(w4389), .C(w3036), .nC(w3318) );
	vdp_slatch g3408 (.Q(w3323), .D(w4390), .C(w3036), .nC(w3318) );
	vdp_slatch g3409 (.Q(w3322), .D(w4391), .C(w3036), .nC(w3318) );
	vdp_slatch g3410 (.Q(w3321), .D(w4392), .C(w3036), .nC(w3318) );
	vdp_slatch g3411 (.Q(w3320), .D(w4393), .C(w3036), .nC(w3318) );
	vdp_slatch g3412 (.Q(w3319), .D(w4394), .C(w3036), .nC(w3318) );
	vdp_slatch g3413 (.Q(w4421), .D(w4395), .C(w3036), .nC(w3318) );
	vdp_slatch g3414 (.Q(w3461), .D(w3455), .C(w3144), .nC(w3452) );
	vdp_slatch g3415 (.Q(w3454), .D(w3151), .C(w3144), .nC(w3452) );
	vdp_slatch g3416 (.Q(w3855), .D(w3453), .C(w3144), .nC(w3452) );
	vdp_slatch g3417 (.Q(w3448), .D(w3451), .C(w3144), .nC(w3452) );
	vdp_slatch g3418 (.Q(w3033), .D(w3093), .C(w3096), .nC(w3095) );
	vdp_slatch g3419 (.Q(w3066), .D(w3067), .C(w3096), .nC(w3095) );
	vdp_slatch g3420 (.Q(w3032), .D(w3069), .C(w3096), .nC(w3095) );
	vdp_slatch g3421 (.Q(w4077), .D(w3070), .C(w3096), .nC(w3095) );
	vdp_slatch g3422 (.Q(w3518), .D(w3071), .C(w3096), .nC(w3095) );
	vdp_slatch g3423 (.Q(w3073), .D(w3094), .C(w3096), .nC(w3095) );
	vdp_slatch g3424 (.Q(w3029), .D(w3098), .C(w3096), .nC(w3095) );
	vdp_slatch g3425 (.Q(w3074), .D(w3097), .C(w3096), .nC(w3095) );
	vdp_cnt_bit_load g3426 (.D(w3453), .nL(w3116), .L(w3113), .R(1'b0), .Q(w3115), .CI(w3514), .CO(w3515), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3427 (.D(w3151), .nL(w3116), .L(w3113), .R(1'b0), .Q(w4011), .CI(w3515), .CO(w3516), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3428 (.D(w3117), .nL(w3116), .L(w3113), .R(1'b0), .Q(w3101), .CI(w3516), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3429 (.CO(w3514), .CI(1'b1), .D(w3451), .nL(w3116), .L(w3113), .R(1'b0), .Q(w3111), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3430 (.CO(w3513), .CI(1'b1), .D(w3448), .nL(w3450), .L(w3143), .R(1'b0), .Q(w3468), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3431 (.CO(w3512), .CI(w3513), .D(w3855), .nL(w3450), .L(w3143), .R(1'b0), .Q(w3414), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3432 (.CO(w3511), .CI(w3512), .D(w3454), .nL(w3450), .L(w3143), .R(1'b0), .Q(w3456), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3433 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .CI(w3511), .D(w3461), .nL(w3450), .L(w3143), .R(1'b0), .Q(w3366) );
	vdp_xor g3434 (.Z(w3254), .B(w4011), .A(w3110) );
	vdp_xor g3435 (.B(w3115), .A(w3110), .Z(w3102) );
	vdp_xor g3436 (.Z(w3257), .B(w3111), .A(w3110) );
	vdp_sr_bit g3437 (.Q(w3109), .D(w4020), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3438 (.Q(w4019), .D(w3109), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3439 (.Q(w3276), .D(w4019), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3440 (.Q(w4028), .D(w3517), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3441 (.Q(w3517), .D(w4029), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3442 (.Q(w4029), .D(w4030), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3443 (.Q(w3031), .D(w3030), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3444 (.Q(w3030), .D(w3028), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3445 (.Q(w3028), .D(w3027), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3446 (.Q(w4032), .D(w4033), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3447 (.Q(w3999), .D(w4032), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3448 (.Q(w4031), .D(w3999), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3449 (.Q(w4036), .D(w4035), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3450 (.Q(w4037), .D(w4036), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3451 (.Q(w4034), .D(w4037), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3452 (.Q(w3123), .D(w4034), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3453 (.Q(w4120), .D(w4121), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3454 (.Q(w4121), .D(w4039), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_xor g3455 (.Z(w3328), .A(w3410), .B(w3456) );
	vdp_xor g3456 (.Z(w3333), .A(w3410), .B(w3467) );
	vdp_xor g3457 (.Z(w3327), .A(w3410), .B(w3468) );
	vdp_dlatch_inv g3458 (.nQ(w4018), .D(w4017), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g3459 (.nQ(w3027), .D(w3072), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g3460 (.nQ(w4033), .D(w3023), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g3461 (.nQ(w3466), .D(w4040), .nC(nHCLK1), .C(HCLK1) );
	vdp_xor g3462 (.Z(w3467), .A(w3414), .B(M5) );
	vdp_sr_bit g3463 (.Q(w3520), .D(w3415), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_dlatch_inv g3464 (.nQ(w4035), .D(w3121), .nC(nDCLK1), .C(DCLK1) );
	vdp_comp_strong g3465 (.Z(w3040), .nZ(w3041), .A(w3317) );
	vdp_comp_strong g3466 (.Z(w3048), .nZ(w3043), .A(w3317) );
	vdp_comp_strong g3467 (.Z(w3045), .nZ(w3046), .A(w3317) );
	vdp_comp_strong g3468 (.Z(w3038), .nZ(w3037), .A(w3317) );
	vdp_comp_strong g3469 (.Z(w3039), .nZ(w3079), .A(w3075) );
	vdp_comp_strong g3470 (.Z(w3042), .nZ(w3080), .A(w3075) );
	vdp_comp_strong g3471 (.Z(w3047), .nZ(w3081), .A(w3075) );
	vdp_comp_strong g3472 (.Z(w3044), .nZ(w3049), .A(w3075) );
	vdp_comp_strong g3473 (.Z(w3052), .nZ(w3077), .A(w3076) );
	vdp_comp_strong g3474 (.Z(w3056), .nZ(w3082), .A(w3385) );
	vdp_comp_strong g3475 (.Z(w3057), .nZ(w3083), .A(w3384) );
	vdp_comp_strong g3476 (.Z(w3059), .nZ(w3078), .A(w3068) );
	vdp_comp_strong g3477 (.Z(w3051), .nZ(w3085), .A(w4027) );
	vdp_comp_strong g3478 (.Z(w3055), .nZ(w3089), .A(w3090) );
	vdp_comp_strong g3479 (.Z(w3058), .nZ(w3086), .A(w3092) );
	vdp_comp_strong g3480 (.Z(w3060), .nZ(w3084), .A(w3091) );
	vdp_comp_strong g3481 (.Z(w3291), .nZ(w3278), .A(w3024) );
	vdp_comp_strong g3482 (.Z(w3099), .nZ(w3279), .A(w3024) );
	vdp_comp_strong g3483 (.Z(w3285), .nZ(w3087), .A(w3024) );
	vdp_comp_strong g3484 (.Z(w3286), .nZ(w3088), .A(w3024) );
	vdp_comp_strong g3485 (.Z(w3290), .nZ(w3292), .A(w3100) );
	vdp_comp_strong g3486 (.Z(w3289), .nZ(w3300), .A(w3100) );
	vdp_comp_strong g3487 (.Z(w3288), .nZ(w3301), .A(w3100) );
	vdp_comp_strong g3488 (.Z(w3287), .nZ(w3293), .A(w3100) );
	vdp_comp_strong g3489 (.Z(w3141), .nZ(w3167), .A(w3100) );
	vdp_comp_strong g3490 (.Z(w3120), .nZ(w3177), .A(w3100) );
	vdp_comp_strong g3491 (.Z(w3132), .nZ(w3178), .A(w3100) );
	vdp_comp_strong g3492 (.Z(w3133), .nZ(w3107), .A(w3100) );
	vdp_comp_strong g3493 (.Z(w3119), .nZ(w3136), .A(w3024) );
	vdp_comp_strong g3494 (.Z(w3137), .nZ(w3128), .A(w3024) );
	vdp_comp_strong g3495 (.Z(w3138), .nZ(w3126), .A(w3024) );
	vdp_comp_strong g3496 (.Z(w3134), .nZ(w3135), .A(w3024) );
	vdp_comp_strong g3497 (.Z(w3149), .nZ(w3139), .A(w3150) );
	vdp_comp_strong g3498 (.Z(w3130), .nZ(w3129), .A(w3152) );
	vdp_comp_strong g3499 (.Z(w3131), .nZ(w3127), .A(w3153) );
	vdp_comp_strong g3500 (.Z(w3148), .nZ(w3140), .A(w3154) );
	vdp_comp_strong g3501 (.Z(w3459), .nZ(w3431), .A(w3274) );
	vdp_comp_strong g3502 (.Z(w3460), .nZ(w3447), .A(w3462) );
	vdp_comp_strong g3503 (.Z(w3458), .nZ(w3434), .A(w3463) );
	vdp_comp_strong g3504 (.Z(w3457), .nZ(w3435), .A(w3464) );
	vdp_comp_strong g3505 (.Z(w3404), .nZ(w3438), .A(w3075) );
	vdp_comp_strong g3506 (.Z(w3430), .nZ(w3432), .A(w3075) );
	vdp_comp_strong g3507 (.Z(w3405), .nZ(w3433), .A(w3075) );
	vdp_comp_strong g3508 (.Z(w3437), .nZ(w3436), .A(w3075) );
	vdp_comp_strong g3509 (.Z(w3439), .nZ(w3440), .A(w3317) );
	vdp_comp_strong g3510 (.Z(w3444), .nZ(w3443), .A(w3317) );
	vdp_comp_strong g3511 (.Z(w3441), .nZ(w3442), .A(w3317) );
	vdp_comp_strong g3512 (.Z(w3445), .nZ(w3446), .A(w3317) );
	vdp_not g3513 (.nZ(w3117), .A(w3455) );
	vdp_not g3514 (.nZ(w4020), .A(w3235) );
	vdp_not g3515 (.nZ(w3237), .A(w98) );
	vdp_not g3516 (.nZ(w3236), .A(w436) );
	vdp_not g3517 (.nZ(w3103), .A(w3236) );
	vdp_comp_strong g3518 (.Z(w3264), .nZ(w3025), .A(w3100) );
	vdp_comp_strong g3519 (.Z(w3284), .nZ(w3316), .A(w3024) );
	vdp_comp_strong g3520 (.Z(w3096), .nZ(w3095), .A(w3274) );
	vdp_comp_strong g3521 (.Z(w3036), .nZ(w3318), .A(w3317) );
	vdp_comp_strong g3522 (.Z(w3035), .nZ(w3034), .A(w3075) );
	vdp_comp_strong g3523 (.Z(w3144), .nZ(w3452), .A(w3520) );
	vdp_not g3524 (.nZ(w3334), .A(w3327) );
	vdp_not g3525 (.nZ(w3326), .A(w3333) );
	vdp_not g3526 (.nZ(w3337), .A(w3328) );
	vdp_nand3 g3527 (.Z(w3331), .A(w3337), .B(w3333), .C(w3327) );
	vdp_not g3528 (.nZ(w3376), .A(w3330) );
	vdp_nand3 g3529 (.Z(w3330), .A(w3328), .B(w3326), .C(w3327) );
	vdp_nand3 g3530 (.Z(w3329), .A(w3328), .B(w3333), .C(w3327) );
	vdp_nand3 g3531 (.Z(w3335), .A(w3328), .B(w3333), .C(w3334) );
	vdp_nand3 g3532 (.Z(w3332), .A(w3337), .B(w3326), .C(w3327) );
	vdp_nand3 g3533 (.Z(w3338), .A(w3337), .B(w3333), .C(w3334) );
	vdp_nand3 g3534 (.Z(w3336), .A(w3328), .B(w3326), .C(w3334) );
	vdp_nand3 g3535 (.Z(w3339), .A(w3334), .B(w3337), .C(w3326) );
	vdp_not g3536 (.nZ(w3377), .A(w3329) );
	vdp_not g3537 (.nZ(w3375), .A(w3331) );
	vdp_not g3538 (.nZ(w3374), .A(w3332) );
	vdp_not g3539 (.nZ(w3372), .A(w3336) );
	vdp_not g3540 (.nZ(w3373), .A(w3335) );
	vdp_not g3541 (.nZ(w3371), .A(w3339) );
	vdp_not g3542 (.nZ(w3370), .A(w3338) );
	vdp_not g3543 (.nZ(w3247), .A(w3257) );
	vdp_not g3544 (.nZ(w3255), .A(w3108) );
	vdp_not g3545 (.nZ(w3246), .A(w3254) );
	vdp_nand3 g3546 (.Z(w3259), .A(w3246), .B(w3108), .C(w3257) );
	vdp_not g3547 (.nZ(w3221), .A(w3261) );
	vdp_nand3 g3548 (.Z(w3261), .A(w3254), .B(w3255), .C(w3257) );
	vdp_nand3 g3549 (.Z(w3260), .A(w3254), .B(w3108), .C(w3257) );
	vdp_nand3 g3550 (.Z(w4026), .A(w3254), .B(w3108), .C(w3247) );
	vdp_nand3 g3551 (.Z(w3258), .A(w3246), .B(w3255), .C(w3257) );
	vdp_nand3 g3552 (.Z(w3256), .A(w3254), .B(w3255), .C(w3247) );
	vdp_not g3553 (.nZ(w3220), .A(w3260) );
	vdp_not g3554 (.nZ(w3226), .A(w3259) );
	vdp_not g3555 (.nZ(w3225), .A(w3258) );
	vdp_not g3556 (.nZ(w3224), .A(w3256) );
	vdp_not g3557 (.nZ(w3223), .A(w4026) );
	vdp_aon22 g3558 (.Z(w3262), .A1(w3265), .B1(w3272), .A2(w3273), .B2(w3026) );
	vdp_aon22 g3559 (.Z(w3263), .A1(w3267), .B1(w3272), .A2(w3273), .B2(w3266) );
	vdp_aon22 g3560 (.Z(w3212), .A1(w3269), .B1(w3272), .A2(w3273), .B2(w3268) );
	vdp_aon22 g3561 (.Z(w3110), .A1(w3271), .B1(w3272), .A2(w3273), .B2(w3270) );
	vdp_sr_bit g3562 (.Q(w3106), .D(w4021), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3563 (.Q(w4021), .D(w3105), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_xor g3564 (.Z(w3108), .A(w3102), .B(1'b1) );
	vdp_xor g3565 (.A(HPOS[3]), .B(w3125), .Z(w4076) );
	vdp_aon22 g3566 (.Z(w3163), .A1(w3156), .B1(w3157), .A2(w3155), .B2(w4075) );
	vdp_aon22 g3567 (.Z(w3164), .A1(w3158), .B1(w3157), .A2(w3155), .B2(w4074) );
	vdp_aon22 g3568 (.Z(w3166), .A1(w3159), .B1(w3157), .A2(w3155), .B2(w4073) );
	vdp_aon22 g3569 (.Z(w3165), .A1(w3160), .B1(w3157), .A2(w3155), .B2(w4072) );
	vdp_aon22 g3570 (.Z(w3601), .A1(w3161), .B1(w3157), .A2(w3155), .B2(w4071) );
	vdp_aon22 g3571 (.Z(w3207), .A1(w3303), .B1(w4013), .A2(w3200), .B2(w3302) );
	vdp_aon22 g3572 (.Z(w3211), .A1(w3303), .B1(w3201), .A2(w3202), .B2(w3302) );
	vdp_aon22 g3573 (.Z(w3209), .A1(w3303), .B1(w3206), .A2(w3205), .B2(w3302) );
	vdp_aon22 g3574 (.Z(w3210), .A1(w3303), .B1(w3203), .A2(w3204), .B2(w3302) );
	vdp_aon222 g3575 (.Z(w3426), .A1(w3418), .B1(w3417), .C1(w3416), .A2(w3364), .B2(w3365), .C2(w3363) );
	vdp_aon222 g3576 (.Z(w3429), .A1(w3422), .B1(w3387), .C1(w3421), .A2(w3364), .B2(w3365), .C2(w3363) );
	vdp_aon222 g3577 (.Z(w3403), .A1(w3423), .B1(w3420), .C1(w3388), .A2(w3364), .B2(w3365), .C2(w3363) );
	vdp_aon222 g3578 (.A1(w3424), .B1(w3389), .C1(w3419), .A2(w3364), .B2(w3365), .C2(w3363), .Z(w3425) );
	vdp_and5 g3579 (.Z(w3465), .A(w3415), .B(w3461), .C(w3454), .D(w3855), .E(w3448) );
	vdp_aon22 g3580 (.Z(w3412), .A1(w3321), .B1(w3521), .A2(w3142), .B2(w3320) );
	vdp_aon22 g3581 (.Z(w3411), .A1(w3323), .B1(w3521), .A2(w3142), .B2(w3322) );
	vdp_aon22 g3582 (.Z(w3410), .A1(w3325), .B1(w3521), .A2(w3142), .B2(w3324) );
	vdp_aon22 g3583 (.Z(w3413), .A1(w3319), .B1(w3521), .A2(w3142), .B2(w4421) );
	vdp_aon22 g3584 (.Z(w3122), .A1(w3407), .B1(w3146), .A2(w3123), .B2(M5) );
	vdp_and4 g3585 (.Z(w3408), .A(w3468), .B(w3414), .C(w3456), .D(w3409) );
	vdp_comp_we g3586 (.Z(w3142), .nZ(w3521), .A(w3406) );
	vdp_comp_we g3587 (.Z(w3302), .nZ(w3303), .A(w3101) );
	vdp_comp_we g3588 (.Z(w3273), .nZ(w3272), .A(w3101) );
	vdp_comp_we g3589 (.Z(w3113), .nZ(w3116), .A(w3195) );
	vdp_comp_we g3590 (.Z(w3155), .nZ(w3157), .A(w3689) );
	vdp_comp_we g3591 (.Z(w3143), .nZ(w3450), .A(w3415) );
	vdp_not g3592 (.nZ(w4041), .A(M5) );
	vdp_dlatch_inv g3593 (.nQ(w4030), .D(w3118), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g3594 (.Z(w3282), .A(DCLK2), .B(w3028) );
	vdp_and g3595 (.Z(w3283), .A(DCLK2), .B(w3027) );
	vdp_and g3596 (.Z(w3281), .A(DCLK2), .B(w3030) );
	vdp_and g3597 (.Z(w3280), .A(DCLK2), .B(w3031) );
	vdp_and g3598 (.Z(w3091), .A(w4030), .B(DCLK2) );
	vdp_and g3599 (.Z(w3092), .A(w4029), .B(DCLK2) );
	vdp_and g3600 (.Z(w3090), .A(w3517), .B(DCLK2) );
	vdp_and g3601 (.Z(w4027), .A(w4028), .B(DCLK2) );
	vdp_and g3602 (.Z(w3076), .A(DCLK2), .B(w4031) );
	vdp_and g3603 (.Z(w3385), .A(DCLK2), .B(w3999) );
	vdp_and g3604 (.Z(w3384), .A(DCLK2), .B(w4032) );
	vdp_and g3605 (.Z(w3068), .A(DCLK2), .B(w4033) );
	vdp_and g3606 (.Z(w3100), .A(w4018), .B(HCLK2) );
	vdp_and g3607 (.Z(w3275), .A(w3237), .B(w3109) );
	vdp_and g3608 (.Z(w3317), .A(w3466), .B(HCLK2) );
	vdp_or g3609 (.Z(w3409), .A(w4041), .B(w3366) );
	vdp_and g3610 (.Z(w3075), .A(w3122), .B(DCLK2) );
	vdp_and g3611 (.Z(w3464), .A(DCLK2), .B(w4035) );
	vdp_and g3612 (.Z(w3463), .A(DCLK2), .B(w4036) );
	vdp_and g3613 (.Z(w3462), .A(DCLK2), .B(w4037) );
	vdp_and g3614 (.Z(w3274), .A(DCLK2), .B(w4034) );
	vdp_and g3615 (.Z(w3406), .A(M5), .B(w3366) );
	vdp_and g3616 (.Z(w4072), .A(w44), .B(HPOS[7]) );
	vdp_and g3617 (.Z(w4071), .A(w44), .B(HPOS[8]) );
	vdp_and g3618 (.Z(w3154), .A(DCLK2), .B(w3147) );
	vdp_and g3619 (.Z(w4073), .A(w44), .B(HPOS[6]) );
	vdp_and g3620 (.Z(w3153), .A(DCLK2), .B(w4022) );
	vdp_and g3621 (.Z(w3152), .A(DCLK2), .B(w3509) );
	vdp_and g3622 (.Z(w3150), .A(DCLK2), .B(w3510) );
	vdp_and g3623 (.Z(w4074), .A(w44), .B(HPOS[5]) );
	vdp_and g3624 (.Z(w3024), .A(DCLK2), .B(w3146) );
	vdp_and g3625 (.Z(w4075), .A(w44), .B(HPOS[4]) );
	vdp_aon22 g3626 (.Z(w3162), .A1(w3124), .B1(w3157), .A2(w3155), .B2(w4076) );
	vdp_and g3627 (.nZ(w3125), .A(w44), .B(M5) );
	vdp_or4 g3628 (.Z(w2846), .D(w3190), .C(w3191), .B(w3192), .A(w3193) );
	vdp_or g3629 (.Z(w3195), .A(w87), .B(w15) );
	vdp_or g3630 (.Z(w3415), .A(w10), .B(w85) );
	vdp_or4 g3631 (.Z(w2847), .A(w3523), .B(w3522), .C(w3507), .D(w3428) );
	vdp_not g3632 (.nZ(w4039), .A(w3369) );
	vdp_not g3633 (.nZ(w3105), .A(w3213) );
	vdp_not g3634 (.nZ(w3407), .A(M5) );
	vdp_aoi21 g3635 (.Z(w3369), .A1(w100), .A2(w3103), .B(w17) );
	vdp_aoi21 g3636 (.Z(w3213), .A1(w101), .A2(w3103), .B(w11) );
	vdp_aoi21 g3637 (.Z(w3235), .A1(w98), .A2(w3103), .B(w4047) );
	vdp_nand4 g3638 (.D(w3101), .C(w3111), .Z(w4017), .A(w4011), .B(w3115) );
	vdp_nand3 g3639 (.Z(w3248), .A(w3246), .B(w3108), .C(w3247) );
	vdp_not g3640 (.nZ(w3228), .A(w3248) );
	vdp_nand3 g3641 (.Z(w3315), .A(w3247), .B(w3246), .C(w3255) );
	vdp_not g3642 (.nZ(w3218), .A(w3315) );
	vdp_not g3643 (.nZ(w3365), .A(w3361) );
	vdp_not g3644 (.nZ(w3364), .A(w3362) );
	vdp_not g3645 (.nZ(w4016), .A(w3366) );
	vdp_not g3646 (.nZ(w3363), .A(M5) );
	vdp_not g3647 (.nZ(w4045), .A(PLANE_A_PRIO) );
	vdp_not g3648 (.nZ(w4023), .A(PLANE_B_PRIO) );
	vdp_bufif0 g3649 (.Z(COL[5]), .A(w3196), .nE(w4023) );
	vdp_bufif0 g3650 (.Z(COL[6]), .A(w3277), .nE(w4023) );
	vdp_bufif0 g3651 (.Z(COL[4]), .A(w3198), .nE(w4023) );
	vdp_bufif0 g3652 (.Z(COL[3]), .A(w3199), .nE(w4023) );
	vdp_bufif0 g3653 (.Z(COL[2]), .A(w3194), .nE(w4023) );
	vdp_bufif0 g3654 (.Z(COL[1]), .A(w3208), .nE(w4023) );
	vdp_bufif0 g3655 (.Z(COL[0]), .A(w3197), .nE(w4023) );
	vdp_bufif0 g3656 (.Z(COL[5]), .A(w3401), .nE(w4045) );
	vdp_bufif0 g3657 (.Z(COL[6]), .A(w3508), .nE(w4045) );
	vdp_bufif0 g3658 (.Z(COL[4]), .A(w3400), .nE(w4045) );
	vdp_bufif0 g3659 (.Z(COL[3]), .A(w3402), .nE(w4045) );
	vdp_bufif0 g3660 (.Z(COL[2]), .A(w3367), .nE(w4045) );
	vdp_bufif0 g3661 (.Z(COL[1]), .A(w4044), .nE(w4045) );
	vdp_bufif0 g3662 (.Z(COL[0]), .A(w3427), .nE(w4045) );
	vdp_nand g3663 (.Z(w3112), .B(HCLK1), .A(w3106) );
	vdp_nand g3664 (.Z(w3118), .B(HCLK1), .A(w3105) );
	vdp_nand g3665 (.Z(w3072), .A(w3618), .B(HCLK1) );
	vdp_nand g3666 (.Z(w3023), .A(w4039), .B(HCLK1) );
	vdp_nor g3667 (.Z(w4040), .A(w3408), .B(w3465) );
	vdp_nand g3668 (.Z(w3121), .A(w4120), .B(HCLK1) );
	vdp_nand g3669 (.Z(w3362), .A(M5), .B(w3366) );
	vdp_nand g3670 (.Z(w3361), .A(M5), .B(w4016) );
	vdp_xor g3671 (.Z(w3538), .A(w3537), .B(w3536) );
	vdp_aon22 g3672 (.Z(w3536), .A1(w3534), .B1(w3613), .A2(VPOS[3]), .B2(w3535) );
	vdp_xnor g3673 (.Z(w3540), .A(w3537), .B(w3614) );
	vdp_aon22 g3674 (.Z(w3614), .A1(w3534), .B1(w3613), .A2(VPOS[2]), .B2(w3539) );
	vdp_xnor g3675 (.Z(w3542), .A(w3537), .B(w3612) );
	vdp_aon22 g3676 (.Z(w3612), .A1(w3534), .B1(w3613), .A2(VPOS[1]), .B2(w3541) );
	vdp_notif0 g3677 (.nZ(VRAMA[4]), .A(w3540), .nE(w3591) );
	vdp_notif0 g3678 (.nZ(VRAMA[3]), .A(w3542), .nE(w3591) );
	vdp_xnor g3679 (.Z(w3610), .A(w3537), .B(w3611) );
	vdp_aon22 g3680 (.Z(w3611), .A1(w3534), .B1(w3613), .A2(VPOS[0]), .B2(w3543) );
	vdp_notif0 g3681 (.nZ(VRAMA[2]), .A(w3610), .nE(w3591) );
	vdp_notif0 g3682 (.nZ(VRAMA[1]), .A(w3609), .nE(w3591) );
	vdp_notif0 g3683 (.nZ(VRAMA[0]), .A(1'b1), .nE(w3591) );
	vdp_not g3684 (.nZ(w3606), .A(w3617) );
	vdp_not g3685 (.nZ(w3591), .A(w3616) );
	vdp_comp_we g3686 (.Z(w3534), .nZ(w3613), .A(w4114) );
	vdp_comp_we g3687 (.Z(w3544), .nZ(w3608), .A(w1) );
	vdp_notif0 g3688 (.nZ(VRAMA[5]), .A(w3546), .nE(w3606) );
	vdp_aoi22 g3689 (.Z(w3546), .A1(w3538), .B1(w3545), .A2(w3544), .B2(w3608) );
	vdp_notif0 g3690 (.nZ(VRAMA[6]), .A(w3547), .nE(w3606) );
	vdp_aoi22 g3691 (.Z(w3547), .A1(w3545), .B1(w3548), .A2(w3544), .B2(w3608) );
	vdp_notif0 g3692 (.nZ(VRAMA[7]), .A(w3549), .nE(w3606) );
	vdp_aoi22 g3693 (.Z(w3549), .A1(w3548), .B1(w3550), .A2(w3544), .B2(w3608) );
	vdp_notif0 g3694 (.nZ(VRAMA[8]), .A(w3551), .nE(w3606) );
	vdp_aoi22 g3695 (.Z(w3551), .A1(w3550), .B1(w3552), .A2(w3544), .B2(w3608) );
	vdp_notif0 g3696 (.nZ(VRAMA[9]), .A(w4049), .nE(w3606) );
	vdp_aoi22 g3697 (.Z(w4049), .A1(w3552), .B1(w3554), .A2(w3544), .B2(w3608) );
	vdp_notif0 g3698 (.nZ(VRAMA[10]), .A(w3553), .nE(w3606) );
	vdp_aoi22 g3699 (.Z(w3553), .A1(w3554), .B1(w3555), .A2(w3544), .B2(w3608) );
	vdp_notif0 g3700 (.nZ(VRAMA[11]), .A(w4048), .nE(w3606) );
	vdp_aoi22 g3701 (.Z(w4048), .A1(w3555), .B1(w3557), .A2(w3544), .B2(w3608) );
	vdp_notif0 g3702 (.nZ(VRAMA[12]), .A(w3558), .nE(w3606) );
	vdp_aoi22 g3703 (.Z(w3558), .A1(w3557), .B1(w3556), .A2(w3544), .B2(w3608) );
	vdp_notif0 g3704 (.nZ(VRAMA[13]), .A(w3560), .nE(w3606) );
	vdp_aoi22 g3705 (.Z(w3560), .A1(w3556), .B1(w3559), .A2(w3544), .B2(w3608) );
	vdp_not g3706 (.nZ(w3607), .A(w4069) );
	vdp_notif0 g3707 (.nZ(VRAMA[14]), .A(w3562), .nE(w3607) );
	vdp_aoi22 g3708 (.Z(w3562), .A1(w3559), .B1(w3561), .A2(w3544), .B2(w3608) );
	vdp_notif0 g3709 (.nZ(VRAMA[15]), .A(w3564), .nE(w3607) );
	vdp_aoi22 g3710 (.Z(w3564), .A1(w3561), .B1(w3563), .A2(w3544), .B2(w3608) );
	vdp_notif0 g3711 (.nZ(VRAMA[16]), .A(w3566), .nE(w3607) );
	vdp_aoi22 g3712 (.Z(w3566), .A1(w3563), .B1(w3565), .A2(w3544), .B2(w3608) );
	vdp_notif0 g3713 (.nZ(VRAMA[5]), .A(w3569), .nE(w3605) );
	vdp_aoi22 g3714 (.Z(w3569), .A1(w3567), .B1(w3538), .A2(w3568), .B2(w3604) );
	vdp_notif0 g3715 (.nZ(VRAMA[6]), .A(w3571), .nE(w3605) );
	vdp_aoi22 g3716 (.Z(w3571), .A1(w3567), .B1(w3568), .A2(w3570), .B2(w3604) );
	vdp_notif0 g3717 (.nZ(VRAMA[7]), .A(w3572), .nE(w3605) );
	vdp_aoi22 g3718 (.Z(w3572), .A1(w3567), .B1(w3570), .A2(w3590), .B2(w3604) );
	vdp_notif0 g3719 (.nZ(VRAMA[8]), .A(w3573), .nE(w3605) );
	vdp_aoi22 g3720 (.Z(w3573), .A1(w3567), .B1(w3590), .A2(w3574), .B2(w3604) );
	vdp_notif0 g3721 (.nZ(VRAMA[9]), .A(w3575), .nE(w3605) );
	vdp_aoi22 g3722 (.Z(w3575), .A1(w3567), .B1(w3574), .A2(w3576), .B2(w3604) );
	vdp_notif0 g3723 (.nZ(VRAMA[10]), .A(w3578), .nE(w3605) );
	vdp_aoi22 g3724 (.Z(w3578), .A1(w3567), .B1(w3576), .A2(w3577), .B2(w3604) );
	vdp_notif0 g3725 (.nZ(VRAMA[11]), .A(w3580), .nE(w3603) );
	vdp_aoi22 g3726 (.Z(w3580), .A1(w3567), .B1(w3577), .A2(w3579), .B2(w3604) );
	vdp_notif0 g3727 (.nZ(VRAMA[12]), .A(w3582), .nE(w3603) );
	vdp_aoi22 g3728 (.Z(w3582), .A1(w3567), .B1(w3579), .A2(w3581), .B2(w3604) );
	vdp_notif0 g3729 (.nZ(VRAMA[14]), .A(w3585), .nE(w3603) );
	vdp_aoi22 g3730 (.Z(w3585), .A1(w3567), .B1(w3583), .A2(w3586), .B2(w3604) );
	vdp_notif0 g3731 (.nZ(VRAMA[15]), .A(w3588), .nE(w3603) );
	vdp_aoi22 g3732 (.Z(w3588), .A1(w3567), .B1(w3586), .A2(w3587), .B2(w3604) );
	vdp_notif0 g3733 (.nZ(VRAMA[16]), .A(w3589), .nE(w3603) );
	vdp_aoi22 g3734 (.Z(w3589), .A1(w3567), .B1(w3587), .A2(w3565), .B2(w3604) );
	vdp_notif0 g3735 (.nZ(VRAMA[13]), .A(w3584), .nE(w3603) );
	vdp_aoi22 g3736 (.Z(w3584), .A1(w3567), .B1(w3581), .A2(w3583), .B2(w3604) );
	vdp_not g3737 (.nZ(w3605), .A(w3533) );
	vdp_comp_we g3738 (.Z(w3604), .nZ(w3567), .A(w1) );
	vdp_aon22 g3739 (.Z(w3565), .A1(w3528), .B1(w3527), .A2(w3529), .B2(w3600) );
	vdp_not g3740 (.nZ(w3603), .A(w3533) );
	vdp_not g3741 (.nZ(w3529), .A(w3600) );
	vdp_sr_bit g3742 (.Q(w3616), .D(w3631), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3743 (.Q(w3600), .D(HPOS[3]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3744 (.Q(w3609), .D(w3668), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3745 (.Q(w3617), .D(w4122), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3746 (.Q(w3615), .D(w4113), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3747 (.Q(w3635), .D(w4112), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3748 (.Q(w3602), .D(w4111), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3749 (.Q(w4087), .D(w4088), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3750 (.Q(w4089), .D(w4087), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3751 (.Q(w3618), .D(w4089), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3752 (.Q(w3650), .D(w104), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3753 (.Q(w3628), .D(w37), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3754 (.Q(w4090), .D(w38), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3755 (.Q(w3690), .D(w4090), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3756 (.Q(w3691), .D(w3628), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3757 (.Q(w3688), .D(w3650), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3758 (.Q(w3692), .D(w3601), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3759 (.Q(w3693), .D(w3165), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3760 (.Q(w3694), .D(w3166), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3761 (.Q(w3695), .D(w3164), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3762 (.Q(w3723), .D(w3163), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3763 (.Q(w3724), .D(w3162), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3764 (.Q(w3626), .D(w3624), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3765 (.Q(w3627), .D(w3626), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3766 (.Q(w4091), .D(w3627), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_aon22 g3767 (.Z(w3640), .A1(H40), .B1(HPOS[8]), .A2(w3638), .B2(w3637) );
	vdp_aon22 g3768 (.Z(w3720), .A1(w3620), .B1(HPOS[8]), .A2(w3640), .B2(w3630) );
	vdp_aon22 g3769 (.Z(w3683), .A1(w3625), .B1(w3638), .A2(w3640), .B2(w3630) );
	vdp_or3 g3770 (.Z(w3689), .A(w3650), .B(w3628), .C(w4090) );
	vdp_or g3771 (.Z(w3641), .A(M5), .B(w3455) );
	vdp_bufif0 g3772 (.Z(VRAMA[1]), .A(w4086), .nE(w3629) );
	vdp_or g3773 (.Z(w3716), .A(w3640), .B(HPOS[4]) );
	vdp_bufif0 g3774 (.Z(VRAMA[2]), .A(w3643), .nE(w3629) );
	vdp_or g3775 (.Z(w3717), .A(w3640), .B(HPOS[5]) );
	vdp_bufif0 g3776 (.Z(VRAMA[3]), .A(w3644), .nE(w3629) );
	vdp_or g3777 (.Z(w3721), .A(w3640), .B(HPOS[6]) );
	vdp_bufif0 g3778 (.Z(VRAMA[4]), .A(w3645), .nE(w3629) );
	vdp_or g3779 (.Z(w3719), .A(w3640), .B(HPOS[7]) );
	vdp_bufif0 g3780 (.Z(VRAMA[5]), .A(w3646), .nE(w3629) );
	vdp_bufif0 g3781 (.Z(VRAMA[5]), .A(w3619), .nE(w3629) );
	vdp_not g3782 (.nZ(w3634), .A(w3526) );
	vdp_not g3783 (.nZ(w4092), .A(HPOS[3]) );
	vdp_dlatch_inv g3784 (.nQ(w3624), .D(w3623), .C(DCLK1), .nC(nDCLK1) );
	vdp_not g3785 (.nZ(w3638), .A(w4068) );
	vdp_not g3786 (.nZ(w3630), .A(w3640) );
	vdp_not g3787 (.nZ(w3637), .A(H40) );
	vdp_not g3788 (.nZ(w3629), .A(w3636) );
	vdp_bufif0 g3789 (.Z(VRAMA[0]), .A(1'b0), .nE(w3629) );
	vdp_or g3790 (.Z(w3636), .A(w3615), .B(w3635) );
	vdp_or g3791 (.Z(w4088), .A(w3633), .B(w6) );
	vdp_nand3 g3792 (.Z(w3687), .A(M5), .B(w3634), .C(HPOS[3]) );
	vdp_nand3 g3793 (.Z(w3648), .A(M5), .B(w3634), .C(w4092) );
	vdp_and g3794 (.Z(w3649), .A(DCLK2), .B(w4091) );
	vdp_and g3795 (.Z(w3622), .A(w3627), .B(DCLK2) );
	vdp_and g3796 (.Z(w3686), .A(w3626), .B(DCLK2) );
	vdp_and g3797 (.Z(w3621), .A(w3624), .B(DCLK2) );
	vdp_and g3798 (.Z(w4069), .A(M5), .B(w3617) );
	vdp_and g3799 (.Z(w3676), .A(HPOS[3]), .B(w3639) );
	vdp_and g3800 (.Z(w4111), .A(w3526), .B(w6) );
	vdp_and g3801 (.Z(w4112), .A(w3634), .B(w6) );
	vdp_and3 g3802 (.Z(w4113), .A(w3633), .B(M5), .C(w3632) );
	vdp_nor g3803 (.Z(w3639), .A(M5), .B(w3640) );
	vdp_nand g3804 (.Z(w3623), .A(w3276), .B(HCLK1) );
	vdp_oai21 g3805 (.A1(HPOS[6]), .A2(HPOS[7]), .B(HPOS[8]), .Z(w4068) );
	vdp_slatch g3806 (.Q(w3665), .D(REG_BUS[0]), .C(w3711), .nC(w3710) );
	vdp_slatch g3807 (.Q(w3661), .D(S[0]), .C(w3706), .nC(w3705) );
	vdp_slatch g3808 (.Q(w3662), .D(S[0]), .C(w3707), .nC(w3704) );
	vdp_slatch g3809 (.Q(w3663), .D(REG_BUS[1]), .C(w3711), .nC(w3710) );
	vdp_slatch g3810 (.Q(w3659), .D(S[1]), .C(w3706), .nC(w3705) );
	vdp_slatch g3811 (.Q(w3732), .D(S[1]), .C(w3707), .nC(w3704) );
	vdp_slatch g3812 (.Q(w3733), .D(REG_BUS[2]), .C(w3711), .nC(w3710) );
	vdp_slatch g3813 (.Q(w3653), .D(S[2]), .C(w3706), .nC(w3705) );
	vdp_slatch g3814 (.Q(w3734), .D(S[2]), .C(w3707), .nC(w3704) );
	vdp_slatch g3815 (.Q(w3730), .D(REG_BUS[3]), .C(w3711), .nC(w3710) );
	vdp_slatch g3816 (.Q(w3729), .D(S[3]), .C(w3706), .nC(w3705) );
	vdp_slatch g3817 (.Q(w4410), .D(S[3]), .C(w3707), .nC(w3704) );
	vdp_slatch g3818 (.Q(w3675), .D(REG_BUS[4]), .C(w3711), .nC(w3710) );
	vdp_slatch g3819 (.Q(w3728), .D(S[4]), .C(w3706), .nC(w3705) );
	vdp_slatch g3820 (.Q(w3727), .D(S[4]), .C(w3707), .nC(w3704) );
	vdp_slatch g3821 (.Q(w3726), .D(REG_BUS[5]), .C(w3711), .nC(w3710) );
	vdp_slatch g3822 (.Q(w3714), .D(S[5]), .C(w3706), .nC(w3705) );
	vdp_slatch g3823 (.Q(w3713), .D(S[5]), .C(w3707), .nC(w3704) );
	vdp_slatch g3824 (.Q(w3712), .D(REG_BUS[6]), .C(w3711), .nC(w3710) );
	vdp_slatch g3825 (.Q(w3708), .D(S[6]), .C(w3706), .nC(w3705) );
	vdp_slatch g3826 (.Q(w3709), .D(S[6]), .C(w3707), .nC(w3704) );
	vdp_slatch g3827 (.Q(w3703), .D(REG_BUS[7]), .C(w3711), .nC(w3710) );
	vdp_slatch g3828 (.Q(w3702), .D(S[7]), .C(w3706), .nC(w3705) );
	vdp_slatch g3829 (.Q(w3701), .D(S[7]), .C(w3707), .nC(w3704) );
	vdp_slatch g3830 (.Q(w3699), .D(S[0]), .C(w3679), .nC(w3696) );
	vdp_slatch g3831 (.Q(w3681), .D(S[0]), .C(w3680), .nC(w3700) );
	vdp_slatch g3832 (.Q(w3685), .D(S[1]), .C(w3680), .nC(w3700) );
	vdp_slatch g3833 (.Q(w3684), .D(S[1]), .C(w3679), .nC(w3696) );
	vdp_slatch g3834 (.Q(w3677), .D(w3703), .C(w3658), .nC(w3657) );
	vdp_slatch g3835 (.Q(w3671), .D(w3712), .C(w3658), .nC(w3657) );
	vdp_slatch g3836 (.Q(w3674), .D(w3726), .C(w3658), .nC(w3657) );
	vdp_slatch g3837 (.Q(w3736), .D(w3675), .C(w3658), .nC(w3657) );
	vdp_slatch g3838 (.Q(w3651), .D(w3730), .C(w3658), .nC(w3657) );
	vdp_slatch g3839 (.Q(w3652), .D(w3733), .C(w3658), .nC(w3657) );
	vdp_slatch g3840 (.Q(w3660), .D(w3663), .C(w3658), .nC(w3657) );
	vdp_slatch g3841 (.Q(w3664), .D(w3665), .C(w3658), .nC(w3657) );
	vdp_fa g3842 (.CI(w4066), .SUM(w4010), .B(w3683), .A(w3698) );
	vdp_fa g3843 (.CO(w4066), .CI(w3682), .SUM(w3882), .B(w3720), .A(w3725) );
	vdp_fa g3844 (.CO(w3725), .CI(w3678), .SUM(w3646), .B(w3719), .A(w4065) );
	vdp_fa g3845 (.CO(w4065), .CI(w3672), .SUM(w3645), .B(w3721), .A(w3722) );
	vdp_fa g3846 (.CO(w3722), .CI(w3673), .SUM(w3644), .B(w3717), .A(w3718) );
	vdp_fa g3847 (.CO(w3718), .CI(w3778), .SUM(w3643), .B(w3716), .A(w3715) );
	vdp_fa g3848 (.CO(w3715), .CI(w3641), .SUM(w4086), .B(w3676), .A(1'b1) );
	vdp_aon222 g3849 (.A1(w3655), .B1(w3642), .C1(w3654), .A2(w3684), .B2(w3685), .C2(1'b0), .Z(w3698) );
	vdp_aon222 g3850 (.A1(w3655), .B1(w3642), .C1(w3654), .A2(w3699), .B2(w3681), .C2(1'b0), .Z(w3682) );
	vdp_aon222 g3851 (.A1(w3655), .B1(w3642), .C1(w3654), .A2(w3701), .B2(w3702), .C2(w3677), .Z(w3678) );
	vdp_aon222 g3852 (.A1(w3655), .B1(w3642), .C1(w3654), .A2(w3709), .B2(w3708), .C2(w3671), .Z(w3672) );
	vdp_aon222 g3853 (.A1(w3655), .B1(w3642), .C1(w3654), .A2(w3713), .B2(w3714), .C2(w3674), .Z(w3673) );
	vdp_aon222 g3854 (.A1(w3655), .B1(w3642), .C1(w3654), .A2(w3727), .B2(w3728), .C2(w3736), .Z(w3778) );
	vdp_aon222 g3855 (.A1(w3655), .B1(w3642), .C1(w3654), .A2(w4410), .B2(w3729), .C2(w3651), .Z(w3455) );
	vdp_aon222 g3856 (.A1(w3655), .B1(w3642), .C1(w3654), .A2(w3734), .B2(w3653), .C2(w3652), .Z(w3151) );
	vdp_aon222 g3857 (.A1(w3655), .B1(w3642), .A2(w3732), .B2(w3659), .C2(w3660), .Z(w3453), .C1(w3654) );
	vdp_aon222 g3858 (.A1(w3655), .B1(w3642), .C1(w3654), .A2(w3662), .B2(w3661), .C2(w3664), .Z(w3451) );
	vdp_comp_strong g3859 (.Z(w3679), .nZ(w3696), .A(w3649) );
	vdp_comp_strong g3860 (.Z(w3680), .nZ(w3700), .A(w3686) );
	vdp_not g3861 (.nZ(w3642), .A(w3648) );
	vdp_not g3862 (.nZ(w3655), .A(w3687) );
	vdp_not g3863 (.nZ(w3654), .A(w3731) );
	vdp_not g3864 (.nZ(w3666), .A(w91) );
	vdp_not g3865 (.nZ(w3632), .A(w99) );
	vdp_not g3866 (.nZ(w3667), .A(w3668) );
	vdp_not g3867 (.nZ(w3633), .A(w3669) );
	vdp_not g3868 (.nZ(w3670), .A(M5) );
	vdp_comp_strong g3869 (.Z(w3706), .nZ(w3705), .A(w3621) );
	vdp_comp_strong g3870 (.Z(w3707), .nZ(w3704), .A(w3622) );
	vdp_comp_strong g3871 (.Z(w3711), .nZ(w3710), .A(w170) );
	vdp_comp_strong g3872 (.Z(w3658), .nZ(w3657), .A(w3735) );
	vdp_or g3873 (.Z(w3731), .A(w4070), .B(M5) );
	vdp_or g3874 (.Z(w4122), .A(w13), .B(w3667) );
	vdp_or g3875 (.Z(w3631), .A(w13), .B(w14) );
	vdp_or g3876 (.Z(w3735), .A(w4), .B(w98) );
	vdp_or5 g3877 (.E(w3666), .C(VPOS[6]), .D(VPOS[5]), .Z(w4070), .A(VPOS[7]), .B(VPOS[4]) );
	vdp_aoi21 g3878 (.Z(w3669), .A1(w99), .A2(w3103), .B(w8) );
	vdp_nand g3879 (.Z(w3668), .A(w14), .B(w3670) );
	vdp_slatch g3880 (.Q(w3772), .D(w4400), .C(w3741), .nC(w3742) );
	vdp_slatch g3881 (.Q(w3747), .D(w4401), .C(w3741), .nC(w3742) );
	vdp_slatch g3882 (.Q(w3748), .D(w4402), .C(w3741), .nC(w3742) );
	vdp_slatch g3883 (.Q(w3749), .D(w4399), .C(w3741), .nC(w3742) );
	vdp_slatch g3884 (.Q(w3751), .D(w4398), .C(w3741), .nC(w3742) );
	vdp_slatch g3885 (.Q(w3750), .D(w4397), .C(w3741), .nC(w3742) );
	vdp_slatch g3886 (.nQ(w3756), .D(w4405), .C(w3743), .nC(w3744) );
	vdp_slatch g3887 (.Q(w3767), .D(w4406), .C(w3743), .nC(w3744) );
	vdp_slatch g3888 (.Q(w3755), .D(w4407), .C(w3743), .nC(w3744) );
	vdp_slatch g3889 (.Q(w3754), .D(w4408), .C(w3743), .nC(w3744) );
	vdp_slatch g3890 (.Q(w3753), .D(w4404), .C(w3743), .nC(w3744) );
	vdp_slatch g3891 (.Q(w3752), .D(w4403), .C(w3743), .nC(w3744) );
	vdp_comp_strong g3892 (.Z(w3741), .nZ(w3742), .A(w3761) );
	vdp_comp_strong g3893 (.Z(w3743), .nZ(w3744), .A(w4093) );
	vdp_cgi2a g3894 (.Z(w4009), .A(w3752), .B(HPOS[4]), .C(1'b1) );
	vdp_cgi2a g3895 (.Z(w4004), .A(w3753), .B(HPOS[5]), .C(w4009) );
	vdp_cgi2a g3896 (.Z(w4003), .A(w3754), .B(HPOS[6]), .C(w4004) );
	vdp_cgi2a g3897 (.Z(w4005), .A(w3755), .B(HPOS[7]), .C(w4003) );
	vdp_cgi2a g3898 (.X(w3757), .A(w3767), .B(HPOS[8]), .C(w4005) );
	vdp_cgi2a g3899 (.Z(w3762), .A(w3759), .B(w3747), .C(w4095) );
	vdp_cgi2a g3900 (.Z(w4095), .A(w3760), .B(w3748), .C(w4006) );
	vdp_cgi2a g3901 (.Z(w4006), .A(w3763), .B(w3749), .C(w4007) );
	vdp_cgi2a g3902 (.Z(w4007), .A(w3766), .B(w3751), .C(w4008) );
	vdp_cgi2a g3903 (.Z(w4008), .A(w3765), .B(w3750), .C(1'b0) );
	vdp_slatch g3904 (.Q(w4400), .D(REG_BUS[7]), .C(w3769), .nC(w3746) );
	vdp_slatch g3905 (.Q(w4401), .D(REG_BUS[4]), .C(w3769), .nC(w3746) );
	vdp_slatch g3906 (.Q(w4402), .D(REG_BUS[3]), .C(w3769), .nC(w3746) );
	vdp_slatch g3907 (.Q(w4399), .D(REG_BUS[2]), .C(w3769), .nC(w3746) );
	vdp_slatch g3908 (.Q(w4398), .D(REG_BUS[1]), .C(w3769), .nC(w3746) );
	vdp_slatch g3909 (.Q(w4397), .D(REG_BUS[0]), .C(w3769), .nC(w3746) );
	vdp_comp_strong g3910 (.Z(w3769), .nZ(w3746), .A(w74) );
	vdp_slatch g3911 (.Q(w4405), .D(REG_BUS[7]), .C(w3770), .nC(w3768) );
	vdp_slatch g3912 (.Q(w4406), .D(REG_BUS[4]), .C(w3770), .nC(w3768) );
	vdp_slatch g3913 (.Q(w4407), .D(REG_BUS[3]), .C(w3770), .nC(w3768) );
	vdp_slatch g3914 (.Q(w4408), .D(REG_BUS[2]), .C(w3770), .nC(w3768) );
	vdp_slatch g3915 (.Q(w4404), .D(REG_BUS[1]), .C(w3770), .nC(w3768) );
	vdp_slatch g3916 (.Q(w4403), .D(REG_BUS[0]), .C(w3770), .nC(w3768) );
	vdp_comp_strong g3917 (.Z(w3770), .nZ(w3768), .A(w168) );
	vdp_xor g3918 (.Z(w3771), .A(w3772), .B(w3762) );
	vdp_xor g3919 (.Z(w3758), .A(w3756), .B(w3757) );
	vdp_aon22 g3920 (.Z(w3759), .A1(w3764), .B1(w3775), .A2(VPOS[8]), .B2(VPOS[7]) );
	vdp_aon22 g3921 (.Z(w3760), .A1(w3764), .B1(w3775), .A2(VPOS[7]), .B2(VPOS[6]) );
	vdp_aon22 g3922 (.Z(w3763), .A1(w3764), .B1(w3775), .A2(VPOS[6]), .B2(VPOS[5]) );
	vdp_aon22 g3923 (.Z(w3766), .A1(w3764), .B1(w3775), .A2(VPOS[5]), .B2(VPOS[4]) );
	vdp_aon22 g3924 (.Z(w3765), .A1(w3764), .B1(w3775), .A2(VPOS[4]), .B2(VPOS[3]) );
	vdp_aon22 g3925 (.Z(w3783), .A1(w3764), .B1(w3775), .A2(VPOS[3]), .B2(VPOS[2]) );
	vdp_aon22 g3926 (.Z(w3782), .A1(w3764), .B1(w3775), .A2(VPOS[2]), .B2(VPOS[1]) );
	vdp_aon22 g3927 (.Z(w3781), .A1(w3764), .B1(w3775), .A2(VPOS[1]), .B2(VPOS[0]) );
	vdp_comp_we g3928 (.Z(w3764), .nZ(w3775), .A(w1) );
	vdp_not g3929 (.nZ(w3526), .A(w4094) );
	vdp_not g3930 (.nZ(w3774), .A(HPOS[3]) );
	vdp_not g3931 (.nZ(w4097), .A(w4096) );
	vdp_or g3932 (.Z(w4093), .A(w98), .B(w4) );
	vdp_or g3933 (.Z(w3761), .A(w98), .B(w4097) );
	vdp_oai21 g3934 (.Z(w4096), .A1(w5), .A2(M5), .B(w4) );
	vdp_and g3935 (.Z(w3773), .A(w3758), .B(w3776) );
	vdp_oai211 g3936 (.Z(w4094), .A1(w3774), .A2(M5), .B(w3773), .C(w3771) );
	vdp_slatch g3937 (.nQ(w3816), .D(REG_BUS[4]), .C(w3788), .nC(w3789) );
	vdp_slatch g3938 (.nQ(w3818), .D(REG_BUS[4]), .C(w3786), .nC(w3787) );
	vdp_slatch g3939 (.nQ(w3817), .D(REG_BUS[5]), .C(w3788), .nC(w3789) );
	vdp_slatch g3940 (.nQ(w3819), .D(REG_BUS[5]), .C(w3786), .nC(w3787) );
	vdp_slatch g3941 (.nQ(w3792), .D(REG_BUS[6]), .C(w3788), .nC(w3789) );
	vdp_slatch g3942 (.nQ(w3793), .D(REG_BUS[6]), .C(w3786), .nC(w3787) );
	vdp_slatch g3943 (.nQ(w4396), .D(REG_BUS[1]), .C(w3786), .nC(w3787) );
	vdp_slatch g3944 (.nQ(w3812), .D(REG_BUS[2]), .C(w3788), .nC(w3789) );
	vdp_slatch g3945 (.nQ(w3813), .D(REG_BUS[2]), .C(w3786), .nC(w3787) );
	vdp_slatch g3946 (.nQ(w3814), .D(REG_BUS[3]), .C(w3788), .nC(w3789) );
	vdp_slatch g3947 (.nQ(w3815), .D(REG_BUS[3]), .C(w3786), .nC(w3787) );
	vdp_slatch g3948 (.nQ(w3820), .D(REG_BUS[0]), .C(w3786), .nC(w3787) );
	vdp_slatch g3949 (.nQ(w3790), .D(REG_BUS[1]), .C(w3788), .nC(w3789) );
	vdp_slatch g3950 (.Q(w3528), .D(REG_BUS[0]), .C(w3779), .nC(w3780) );
	vdp_slatch g3951 (.Q(w3527), .D(REG_BUS[4]), .C(w3779), .nC(w3780) );
	vdp_not g3952 (.nZ(w4099), .A(w3790) );
	vdp_aoi22 g3953 (.Z(w3809), .A1(HPOS[8]), .B1(w3765), .A2(w3785), .B2(w3784) );
	vdp_aoi22 g3954 (.Z(w3810), .A1(w3765), .B1(w3766), .A2(w3785), .B2(w3784) );
	vdp_aoi22 g3955 (.Z(w3797), .A1(w3766), .B1(w3763), .A2(w3785), .B2(w3784) );
	vdp_aoi22 g3956 (.Z(w3822), .A1(w3760), .B1(w3759), .A2(w3785), .B2(w3784) );
	vdp_aoi22 g3957 (.Z(w3811), .A1(w3763), .B1(w3760), .A2(w3785), .B2(w3784) );
	vdp_comp_strong g3958 (.Z(w3779), .nZ(w3780), .A(w169) );
	vdp_comp_strong g3959 (.Z(w3788), .nZ(w3789), .A(w71) );
	vdp_comp_strong g3960 (.Z(w3786), .nZ(w3787), .A(w68) );
	vdp_aoi22 g3961 (.Z(w3821), .A1(w3759), .B1(w3784), .A2(w3785), .B2(w4099) );
	vdp_nand g3962 (.Z(w3823), .A(w3759), .B(w88) );
	vdp_nand g3963 (.Z(w3796), .A(w3760), .B(w88) );
	vdp_nand g3964 (.Z(w3824), .A(w3766), .B(w88) );
	vdp_nand g3965 (.Z(w3798), .A(w3763), .B(w88) );
	vdp_nand g3966 (.Z(w3808), .A(w3765), .B(w88) );
	vdp_nand g3967 (.Z(w4098), .A(w3783), .B(w86) );
	vdp_nand g3968 (.Z(w4123), .A(w3782), .B(w86) );
	vdp_nand g3969 (.Z(w3804), .A(w3781), .B(w86) );
	vdp_nand g3970 (.Z(w3776), .A(HPOS[7]), .B(HPOS[8]) );
	vdp_comp_we g3971 (.Z(w3785), .nZ(w3784), .A(H40) );
	vdp_notif0 g3972 (.nZ(VRAMA[16]), .A(w3793), .nE(w3791) );
	vdp_notif0 g3973 (.nZ(VRAMA[16]), .A(w3792), .nE(w3795) );
	vdp_notif0 g3974 (.nZ(VRAMA[15]), .A(w3819), .nE(w3791) );
	vdp_notif0 g3975 (.nZ(VRAMA[15]), .A(w3817), .nE(w3795) );
	vdp_notif0 g3976 (.nZ(VRAMA[14]), .A(w3818), .nE(w3791) );
	vdp_notif0 g3977 (.nZ(VRAMA[14]), .A(w3816), .nE(w3795) );
	vdp_notif0 g3978 (.nZ(VRAMA[13]), .A(w3815), .nE(w3791) );
	vdp_notif0 g3979 (.nZ(VRAMA[13]), .A(w3814), .nE(w3795) );
	vdp_notif0 g3980 (.nZ(VRAMA[12]), .A(w3813), .nE(w3791) );
	vdp_notif0 g3981 (.nZ(VRAMA[12]), .A(w3812), .nE(w3795) );
	vdp_notif0 g3982 (.nZ(VRAMA[11]), .A(w4396), .nE(w3791) );
	vdp_notif0 g3983 (.nZ(VRAMA[11]), .A(w3821), .nE(w3795) );
	vdp_notif0 g3984 (.nZ(VRAMA[10]), .A(w3820), .nE(w3791) );
	vdp_notif0 g3985 (.nZ(VRAMA[10]), .A(w3822), .nE(w3795) );
	vdp_notif0 g3986 (.nZ(VRAMA[9]), .A(w3823), .nE(w3794) );
	vdp_notif0 g3987 (.nZ(VRAMA[9]), .A(w3811), .nE(w3795) );
	vdp_notif0 g3988 (.nZ(VRAMA[6]), .A(w3824), .nE(w3794) );
	vdp_notif0 g3989 (.nZ(VRAMA[6]), .A(w3809), .nE(w3799) );
	vdp_notif0 g3990 (.nZ(VRAMA[5]), .A(w3808), .nE(w3794) );
	vdp_notif0 g3991 (.nZ(VRAMA[5]), .A(w3807), .nE(w3799) );
	vdp_notif0 g3992 (.nZ(VRAMA[4]), .A(w4098), .nE(w3794) );
	vdp_notif0 g3993 (.nZ(VRAMA[4]), .A(w3806), .nE(w3799) );
	vdp_notif0 g3994 (.nZ(VRAMA[3]), .A(w4123), .nE(w3794) );
	vdp_notif0 g3995 (.nZ(VRAMA[3]), .A(w3805), .nE(w3799) );
	vdp_notif0 g3996 (.nZ(VRAMA[2]), .A(w3804), .nE(w3794) );
	vdp_notif0 g3997 (.nZ(VRAMA[2]), .A(w3803), .nE(w3799) );
	vdp_notif0 g3998 (.nZ(VRAMA[1]), .A(1'b1), .nE(w3794) );
	vdp_notif0 g3999 (.nZ(VRAMA[1]), .A(1'b1), .nE(w3799) );
	vdp_notif0 g4000 (.nZ(VRAMA[0]), .A(w3801), .nE(w3794) );
	vdp_notif0 g4001 (.nZ(VRAMA[0]), .A(w3801), .nE(w3799) );
	vdp_notif0 g4002 (.nZ(VRAMA[8]), .A(w3796), .nE(w3794) );
	vdp_notif0 g4003 (.nZ(VRAMA[8]), .A(w3797), .nE(w3799) );
	vdp_notif0 g4004 (.nZ(VRAMA[7]), .A(w3798), .nE(w3794) );
	vdp_notif0 g4005 (.nZ(VRAMA[7]), .A(w3810), .nE(w3799) );
	vdp_not g4006 (.nZ(w3801), .A(1'b0) );
	vdp_not g4007 (.nZ(w3803), .A(HPOS[4]) );
	vdp_not g4008 (.nZ(w3805), .A(HPOS[5]) );
	vdp_not g4009 (.nZ(w3806), .A(HPOS[6]) );
	vdp_not g4010 (.nZ(w3807), .A(HPOS[7]) );
	vdp_not g4011 (.nZ(w3794), .A(w3275) );
	vdp_not g4012 (.nZ(w3791), .A(w3275) );
	vdp_not g4013 (.nZ(w3799), .A(w3602) );
	vdp_not g4014 (.nZ(w3795), .A(w3602) );
	vdp_not g4015 (.nZ(w3833), .A(w4002) );
	vdp_comp_strong g4016 (.Z(w3827), .nZ(w3828), .A(w70) );
	vdp_comp_we g4017 (.Z(w3832), .nZ(w3831), .A(w3615) );
	vdp_comp_strong g4018 (.Z(w3830), .nZ(w3829), .A(w72) );
	vdp_slatch g4019 (.Q(w3853), .D(REG_BUS[6]), .C(w3827), .nC(w3828) );
	vdp_slatch g4020 (.Q(w4108), .D(REG_BUS[3]), .C(w3830), .nC(w3829) );
	vdp_slatch g4021 (.Q(w3852), .D(REG_BUS[5]), .C(w3827), .nC(w3828) );
	vdp_slatch g4022 (.Q(w3850), .D(REG_BUS[2]), .C(w3830), .nC(w3829) );
	vdp_slatch g4023 (.Q(w3836), .D(REG_BUS[4]), .C(w3827), .nC(w3828) );
	vdp_slatch g4024 (.Q(w4411), .D(REG_BUS[1]), .C(w3830), .nC(w3829) );
	vdp_slatch g4025 (.Q(w3839), .D(REG_BUS[3]), .C(w3827), .nC(w3828) );
	vdp_slatch g4026 (.Q(w4109), .D(REG_BUS[0]), .C(w3830), .nC(w3829) );
	vdp_slatch g4027 (.Q(w3847), .D(REG_BUS[1]), .C(w3827), .nC(w3828) );
	vdp_slatch g4028 (.Q(w3844), .D(REG_BUS[2]), .C(w3827), .nC(w3828) );
	vdp_bufif0 g4029 (.Z(VRAMA[11]), .A(w3846), .nE(w3835) );
	vdp_bufif0 g4030 (.Z(VRAMA[10]), .A(w3840), .nE(w3835) );
	vdp_bufif0 g4031 (.Z(VRAMA[13]), .A(w3848), .nE(w3835) );
	vdp_bufif0 g4032 (.Z(VRAMA[9]), .A(w3838), .nE(w3835) );
	vdp_bufif0 g4033 (.Z(VRAMA[8]), .A(w3837), .nE(w3835) );
	vdp_bufif0 g4034 (.Z(VRAMA[14]), .A(w3849), .nE(w3833) );
	vdp_bufif0 g4035 (.Z(VRAMA[7]), .A(w3834), .nE(w3835) );
	vdp_bufif0 g4036 (.Z(VRAMA[15]), .A(w4067), .nE(w3833) );
	vdp_bufif0 g4037 (.Z(VRAMA[16]), .A(w3851), .nE(w3833) );
	vdp_aon22 g4038 (.Z(w3851), .A1(w3831), .B1(w3832), .A2(w3853), .B2(w4108) );
	vdp_aon22 g4039 (.Z(w4067), .A1(w3831), .B1(w3832), .A2(w3852), .B2(w3850) );
	vdp_aon22 g4040 (.Z(w3849), .A1(w3831), .B1(w3832), .A2(w3836), .B2(w4411) );
	vdp_aon22 g4041 (.Z(w3848), .A1(w3831), .B1(w3832), .A2(w3839), .B2(w4109) );
	vdp_aon22 g4042 (.Z(w3846), .A1(w3842), .B1(w3845), .A2(w3847), .B2(w3843) );
	vdp_aon22 g4043 (.Z(w3841), .A1(w3842), .B1(w3856), .A2(w3844), .B2(w3843) );
	vdp_bufif0 g4044 (.Z(VRAMA[12]), .A(w3841), .nE(w3835) );
	vdp_not g4045 (.nZ(w3835), .A(w3636) );
	vdp_and g4046 (.Z(w4002), .A(w3636), .B(M5) );
	vdp_comp_we g4047 (.Z(w3843), .nZ(w3842), .A(M5) );
	vdp_fa g4048 (.CO(w3871), .CI(w4056), .SUM(w3891), .B(VPOS[6]), .A(w4055) );
	vdp_fa g4049 (.CO(w4055), .CI(w4058), .SUM(w3872), .B(VPOS[5]), .A(w4057) );
	vdp_fa g4050 (.CO(w4057), .CI(w4060), .SUM(w3873), .B(VPOS[4]), .A(w4059) );
	vdp_fa g4051 (.CO(w4059), .CI(w3939), .SUM(w3535), .B(VPOS[3]), .A(w4061) );
	vdp_fa g4052 (.CO(w4061), .CI(w4063), .SUM(w3539), .B(VPOS[2]), .A(w4062) );
	vdp_fa g4053 (.CO(w4062), .CI(w3997), .SUM(w3541), .B(VPOS[1]), .A(w4064) );
	vdp_fa g4054 (.CO(w4064), .CI(w3952), .SUM(w3543), .B(VPOS[0]), .A(1'b0) );
	vdp_fa g4055 (.CO(w3890), .CI(w4054), .SUM(w3888), .B(VPOS[7]), .A(w3871) );
	vdp_fa g4056 (.CO(w3870), .CI(w3925), .SUM(w3899), .B(VPOS[8]), .A(w3890) );
	vdp_fa g4057 (.CO(w3898), .CI(w3926), .SUM(w3865), .B(1'b0), .A(w3870) );
	vdp_fa g4058 (.CI(w3910), .SUM(w3866), .B(1'b0), .A(w3898) );
	vdp_aon22 g4059 (.Z(w3910), .A1(w3908), .B1(w3909), .A2(w3869), .B2(w3868) );
	vdp_aon22 g4060 (.Z(w3926), .A1(w4000), .B1(w3913), .A2(w3869), .B2(w3868) );
	vdp_aon22 g4061 (.Z(w3925), .A1(w3914), .B1(w3915), .A2(w3869), .B2(w3868) );
	vdp_aon22 g4062 (.Z(w4054), .A1(w3917), .B1(w3918), .A2(w3869), .B2(w3868) );
	vdp_aon22 g4063 (.Z(w4056), .A1(w3924), .B1(w3921), .A2(w3869), .B2(w3868) );
	vdp_aon22 g4064 (.Z(w4058), .A1(w3929), .B1(w3928), .A2(w3869), .B2(w3868) );
	vdp_aon22 g4065 (.Z(w4060), .A1(w3933), .B1(w3934), .A2(w3869), .B2(w3868) );
	vdp_aon22 g4066 (.Z(w3939), .A1(w3938), .B1(w3937), .A2(w3869), .B2(w3868) );
	vdp_aon22 g4067 (.Z(w4063), .A1(w3940), .B1(w3941), .A2(w3869), .B2(w3868) );
	vdp_aon22 g4068 (.Z(w3997), .A1(w3944), .B1(w4001), .A2(w3869), .B2(w3868) );
	vdp_aon22 g4069 (.Z(w3952), .A1(w3946), .B1(w3945), .A2(w3869), .B2(w3868) );
	vdp_comp_we g4070 (.Z(w3869), .nZ(w3868), .A(w3877) );
	vdp_comp_strong g4071 (.Z(w3879), .nZ(w3874), .A(w69) );
	vdp_sr_bit g4072 (.Q(w3900), .D(RD_DATA[1]), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4073 (.Q(w3875), .D(RD_DATA[2]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4074 (.Q(w3949), .D(w3900), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4075 (.Q(w3967), .D(w3875), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4076 (.Q(w3948), .D(HPOS[3]), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4077 (.Q(w3620), .D(REG_BUS[0]), .C(w3879), .nC(w3874) );
	vdp_slatch g4078 (.Q(w3625), .D(REG_BUS[1]), .C(w3879), .nC(w3874) );
	vdp_slatch g4079 (.Q(w3895), .D(REG_BUS[5]), .C(w3879), .nC(w3874) );
	vdp_slatch g4080 (.Q(w3894), .D(REG_BUS[4]), .C(w3879), .nC(w3874) );
	vdp_slatch g4081 (.Q(w3946), .D(w3950), .C(w3901), .nC(w3905) );
	vdp_slatch g4082 (.Q(w4119), .D(w3951), .C(w3907), .nC(w3902) );
	vdp_slatch g4083 (.Q(w3944), .D(w3943), .C(w3901), .nC(w3905) );
	vdp_slatch g4084 (.Q(w4118), .D(w3942), .C(w3907), .nC(w3902) );
	vdp_slatch g4085 (.Q(w3940), .D(w3969), .C(w3901), .nC(w3905) );
	vdp_slatch g4086 (.Q(w4117), .D(w3936), .C(w3907), .nC(w3902) );
	vdp_slatch g4087 (.Q(w3938), .D(w3935), .C(w3901), .nC(w3905) );
	vdp_slatch g4088 (.Q(w4116), .D(w3932), .C(w3907), .nC(w3902) );
	vdp_slatch g4089 (.Q(w3933), .D(w3931), .C(w3901), .nC(w3905) );
	vdp_slatch g4090 (.Q(w4115), .D(w3930), .C(w3907), .nC(w3902) );
	vdp_slatch g4091 (.Q(w3929), .D(w3923), .C(w3901), .nC(w3905) );
	vdp_slatch g4092 (.Q(w4126), .D(w3922), .C(w3907), .nC(w3902) );
	vdp_slatch g4093 (.Q(w3924), .D(w3919), .C(w3901), .nC(w3905) );
	vdp_slatch g4094 (.Q(w4127), .D(w3920), .C(w3907), .nC(w3902) );
	vdp_slatch g4095 (.Q(w3917), .D(w3916), .C(w3901), .nC(w3905) );
	vdp_slatch g4096 (.Q(w3915), .D(w3927), .C(w3907), .nC(w3902) );
	vdp_slatch g4097 (.Q(w3914), .D(w3974), .C(w3901), .nC(w3905) );
	vdp_slatch g4098 (.Q(w3913), .D(w3912), .C(w3907), .nC(w3902) );
	vdp_slatch g4099 (.Q(w4000), .D(w3911), .C(w3901), .nC(w3905) );
	vdp_slatch g4100 (.Q(w3909), .D(w3989), .C(w3907), .nC(w3902) );
	vdp_slatch g4101 (.Q(w3908), .D(w3906), .C(w3901), .nC(w3905) );
	vdp_slatch g4102 (.Q(w4102), .D(REG_BUS[0]), .C(w3958), .nC(w3957) );
	vdp_aon22 g4103 (.Z(w3947), .A1(w3950), .B1(w3966), .A2(w3968), .B2(w4102) );
	vdp_slatch g4104 (.Q(w3970), .D(REG_BUS[1]), .C(w3958), .nC(w3957) );
	vdp_aon22 g4105 (.Z(w3951), .A1(w3943), .B1(w3966), .A2(w3968), .B2(w3970) );
	vdp_slatch g4106 (.Q(w4101), .D(REG_BUS[2]), .C(w3958), .nC(w3957) );
	vdp_aon22 g4107 (.Z(w3942), .A1(w3969), .B1(w3966), .A2(w3968), .B2(w4101) );
	vdp_slatch g4108 (.Q(w3971), .D(REG_BUS[3]), .C(w3958), .nC(w3957) );
	vdp_aon22 g4109 (.Z(w3936), .A1(w3935), .B1(w3966), .A2(w3968), .B2(w3971) );
	vdp_slatch g4110 (.Q(w3972), .D(REG_BUS[4]), .C(w3958), .nC(w3957) );
	vdp_aon22 g4111 (.Z(w3932), .A1(w3931), .B1(w3966), .A2(w3968), .B2(w3972) );
	vdp_slatch g4112 (.Q(w3998), .D(REG_BUS[5]), .C(w3958), .nC(w3957) );
	vdp_aon22 g4113 (.Z(w3930), .A1(w3923), .B1(w3966), .A2(w3968), .B2(w3998) );
	vdp_slatch g4114 (.Q(w4100), .D(REG_BUS[6]), .C(w3958), .nC(w3957) );
	vdp_aon22 g4115 (.Z(w3922), .A1(w3919), .B1(w3966), .A2(w3968), .B2(w4100) );
	vdp_slatch g4116 (.Q(w3973), .D(REG_BUS[7]), .C(w3958), .nC(w3957) );
	vdp_aon22 g4117 (.Z(w3920), .A1(w3916), .B1(w3966), .A2(w3968), .B2(w3973) );
	vdp_aon22 g4118 (.Z(w3927), .A1(w3974), .B1(w3966), .A2(w3968), .B2(1'b0) );
	vdp_aon22 g4119 (.Z(w3912), .A1(w3911), .B1(w3966), .A2(w3968), .B2(1'b0) );
	vdp_aon22 g4120 (.Z(w3989), .A1(w3906), .B1(w3966), .A2(w3968), .B2(1'b0) );
	vdp_notif0 g4121 (.nZ(RD_DATA[2]), .A(w3990), .nE(w3962) );
	vdp_slatch g4122 (.nQ(w3990), .D(w3906), .C(w3961), .nC(w3960) );
	vdp_notif0 g4123 (.nZ(RD_DATA[1]), .A(w3975), .nE(w3962) );
	vdp_slatch g4124 (.nQ(w3975), .D(w3911), .C(w3961), .nC(w3960) );
	vdp_notif0 g4125 (.nZ(RD_DATA[0]), .A(w4125), .nE(w3962) );
	vdp_slatch g4126 (.nQ(w4125), .D(w3974), .C(w3961), .nC(w3960) );
	vdp_notif0 g4127 (.nZ(AD_DATA[7]), .A(w4420), .nE(w3962) );
	vdp_slatch g4128 (.nQ(w4420), .D(w3916), .C(w3961), .nC(w3960) );
	vdp_notif0 g4129 (.nZ(AD_DATA[6]), .A(w3976), .nE(w3962) );
	vdp_slatch g4130 (.nQ(w3976), .D(w3919), .C(w3961), .nC(w3960) );
	vdp_notif0 g4131 (.nZ(AD_DATA[5]), .A(w3977), .nE(w3962) );
	vdp_slatch g4132 (.nQ(w3977), .D(w3923), .C(w3961), .nC(w3960) );
	vdp_notif0 g4133 (.nZ(AD_DATA[4]), .A(w3978), .nE(w3962) );
	vdp_slatch g4134 (.nQ(w3978), .D(w3931), .C(w3961), .nC(w3960) );
	vdp_notif0 g4135 (.nZ(AD_DATA[3]), .A(w3987), .nE(w3962) );
	vdp_slatch g4136 (.nQ(w3987), .D(w3935), .C(w3961), .nC(w3960) );
	vdp_notif0 g4137 (.nZ(AD_DATA[2]), .A(w3985), .nE(w3962) );
	vdp_slatch g4138 (.nQ(w3985), .D(w3969), .C(w3961), .nC(w3960) );
	vdp_notif0 g4139 (.nZ(AD_DATA[1]), .A(w3980), .nE(w3962) );
	vdp_slatch g4140 (.nQ(w3980), .D(w3943), .C(w3961), .nC(w3960) );
	vdp_notif0 g4141 (.nZ(AD_DATA[0]), .A(w3984), .nE(w3962) );
	vdp_slatch g4142 (.nQ(w3984), .D(w3950), .C(w3961), .nC(w3960) );
	vdp_sr_bit g4143 (.Q(w3983), .D(w3688), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4144 (.Q(w3991), .D(w3995), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4145 (.Q(w3995), .D(RD_DATA[0]), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4146 (.Q(w4124), .D(w3947), .C(w3907), .nC(w3902) );
	vdp_comp_strong g4147 (.Z(w3907), .nZ(w3902), .A(w3965) );
	vdp_comp_strong g4148 (.Z(w3901), .nZ(w3905), .A(w3963) );
	vdp_comp_strong g4149 (.Z(w3958), .nZ(w3957), .A(w171) );
	vdp_sr_bit g4150 (.Q(w3903), .D(w4105), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_comp_strong g4151 (.Z(w3961), .nZ(w3960), .A(w3982) );
	vdp_not g4152 (.nZ(w3962), .A(w3983) );
	vdp_and g4153 (.Z(w3982), .A(w3688), .B(HCLK1) );
	vdp_and g4154 (.Z(w3918), .A(w4127), .B(w3903) );
	vdp_and g4155 (.Z(w3921), .A(w4126), .B(w3903) );
	vdp_and g4156 (.Z(w3928), .A(w4115), .B(w3903) );
	vdp_and g4157 (.Z(w3934), .A(w4116), .B(w3903) );
	vdp_and g4158 (.Z(w3937), .A(w4117), .B(w3903) );
	vdp_and g4159 (.Z(w3941), .A(w4118), .B(w3903) );
	vdp_and g4160 (.Z(w4001), .A(w4119), .B(w3903) );
	vdp_and g4161 (.Z(w3945), .A(w4124), .B(w3903) );
	vdp_not g4162 (.nZ(w4104), .A(w4103) );
	vdp_not g4163 (.nZ(w3963), .A(w3964) );
	vdp_not g4164 (.nZ(w3877), .A(w3876) );
	vdp_not g4165 (.nZ(w3881), .A(w3620) );
	vdp_not g4166 (.nZ(w3880), .A(w3625) );
	vdp_not g4167 (.nZ(w3858), .A(w4106) );
	vdp_not g4168 (.nZ(w3857), .A(w4107) );
	vdp_not g4169 (.nZ(w3859), .A(w4110) );
	vdp_not g4170 (.nZ(w4053), .A(M5) );
	vdp_not g4171 (.nZ(w3897), .A(w4052) );
	vdp_aon22 g4172 (.Z(w3885), .A1(w3864), .B1(w3872), .A2(w3891), .B2(w3867) );
	vdp_aon22 g4173 (.Z(w3889), .A1(w3864), .B1(w3891), .A2(w3888), .B2(w3867) );
	vdp_ha g4174 (.CO(w3893), .SUM(w3863), .B(w3892), .A(w3889) );
	vdp_aon222 g4175 (.A1(w3859), .B1(w3857), .C1(w3858), .A2(w3887), .B2(w3886), .C2(w3863), .Z(w3838) );
	vdp_aon22 g4176 (.Z(w4051), .A1(w3864), .B1(w3888), .A2(w3899), .B2(w3867) );
	vdp_ha g4177 (.SUM(w3862), .B(w3893), .A(w4051) );
	vdp_aon222 g4178 (.A1(w3859), .B1(w3857), .C1(w3858), .A2(w3886), .B2(w3863), .C2(w3862), .Z(w3840) );
	vdp_ha g4179 (.CO(w3892), .SUM(w3886), .B(w3885), .A(w3896) );
	vdp_aon222 g4180 (.A1(w3859), .B1(w3857), .C1(w3858), .A2(w3883), .B2(w3887), .C2(w3886), .Z(w3837) );
	vdp_aon22 g4181 (.Z(w3887), .A1(w3864), .B1(w3873), .A2(w3872), .B2(w3867) );
	vdp_aon222 g4182 (.A1(w3859), .B1(w3857), .C1(w3858), .A2(w4010), .B2(w3883), .C2(w3887), .Z(w3834) );
	vdp_aon222 g4183 (.A1(w3859), .B1(w3857), .C1(w3858), .A2(w3882), .B2(w3882), .C2(w3883), .Z(w3619) );
	vdp_aon22 g4184 (.Z(w3883), .A1(w3864), .B1(w3535), .A2(w3873), .B2(w3867) );
	vdp_comp_we g4185 (.Z(w3968), .nZ(w3966), .A(M5) );
	vdp_comp_we g4186 (.Z(w3864), .nZ(w3867), .A(w1) );
	vdp_and g4187 (.Z(w3896), .A(w3897), .B(w4053) );
	vdp_aon222 g4188 (.A1(w3859), .B1(w3857), .C1(w3858), .A2(w3863), .B2(w3862), .C2(w3860), .Z(w3845) );
	vdp_aon222 g4189 (.A1(w3859), .B1(w3857), .C1(w3858), .A2(w3862), .B2(w3860), .C2(w4050), .Z(w3856) );
	vdp_aon22 g4190 (.Z(w3861), .A1(w3864), .B1(w3865), .A2(w3866), .B2(w3867) );
	vdp_aon22 g4191 (.Z(w3884), .A1(w3864), .B1(w3899), .A2(w3865), .B2(w3867) );
	vdp_and g4192 (.Z(w3860), .B(w3884), .A(w3894) );
	vdp_and g4193 (.Z(w4050), .B(w3861), .A(w3895) );
	vdp_oai21 g4194 (.Z(w3876), .A1(w44), .A2(w3948), .B(M5) );
	vdp_aoi21 g4195 (.Z(w3964), .A1(HCLK1), .A2(w16), .B(w98) );
	vdp_oai211 g4196 (.Z(w4103), .A1(HCLK1), .A2(w4), .B(w5), .C(M5) );
	vdp_or g4197 (.Z(w3965), .A(w98), .B(w4104) );
	vdp_nand3 g4198 (.Z(w4105), .A(w90), .B(HPOS[6]), .C(HPOS[7]) );
	vdp_nand g4199 (.Z(w4110), .A(w3625), .B(w3620) );
	vdp_nand g4200 (.Z(w4107), .A(w3620), .B(w3880) );
	vdp_nand g4201 (.Z(w4106), .A(w3880), .B(w3881) );
	vdp_aoi31 g4202 (.Z(w4052), .B3(w4051), .B2(w3889), .B1(w3885), .A(w3884) );
	vdp_slatch g4203 (.Q(w3568), .D(S[0]), .C(w3530), .nC(w3145) );
	vdp_slatch g4204 (.Q(w3570), .D(S[1]), .C(w3530), .nC(w3145) );
	vdp_slatch g4205 (.Q(w3590), .D(S[2]), .C(w3530), .nC(w3145) );
	vdp_slatch g4206 (.Q(w3574), .D(S[3]), .C(w3530), .nC(w3145) );
	vdp_slatch g4207 (.Q(w3576), .D(S[4]), .C(w3530), .nC(w3145) );
	vdp_slatch g4208 (.Q(w3577), .D(S[5]), .C(w3530), .nC(w3145) );
	vdp_slatch g4209 (.Q(w3579), .D(S[6]), .C(w3530), .nC(w3145) );
	vdp_slatch g4210 (.Q(w3581), .D(S[7]), .C(w3530), .nC(w3145) );
	vdp_slatch g4211 (.Q(w3583), .D(S[0]), .C(w3525), .nC(w3524) );
	vdp_slatch g4212 (.Q(w3586), .D(S[1]), .C(w3525), .nC(w3524) );
	vdp_slatch g4213 (.Q(w3587), .D(S[2]), .C(w3525), .nC(w3524) );
	vdp_slatch g4214 (.Q(w3093), .D(S[3]), .C(w3525), .nC(w3524) );
	vdp_slatch g4215 (.Q(w3594), .D(S[4]), .C(w3525), .nC(w3524) );
	vdp_slatch g4216 (.Q(w3069), .D(S[5]), .C(w3525), .nC(w3524) );
	vdp_slatch g4217 (.Q(w3071), .D(S[6]), .C(w3525), .nC(w3524) );
	vdp_slatch g4218 (.Q(w3098), .D(S[7]), .C(w3525), .nC(w3524) );
	vdp_comp_strong g4219 (.Z(w3525), .nZ(w3524), .A(w3280) );
	vdp_comp_strong g4220 (.Z(w3530), .nZ(w3145), .A(w3281) );
	vdp_comp_strong g4221 (.Z(w3531), .nZ(w3592), .A(w3282) );
	vdp_slatch g4222 (.Q(w4085), .D(S[7]), .C(w3531), .nC(w3592) );
	vdp_slatch g4223 (.Q(w4084), .D(S[6]), .C(w3531), .nC(w3592) );
	vdp_slatch g4224 (.Q(w4083), .D(S[5]), .C(w3531), .nC(w3592) );
	vdp_slatch g4225 (.Q(w3597), .D(S[4]), .C(w3531), .nC(w3592) );
	vdp_slatch g4226 (.Q(w3598), .D(S[3]), .C(w3531), .nC(w3592) );
	vdp_slatch g4227 (.Q(w3563), .D(S[2]), .C(w3531), .nC(w3592) );
	vdp_slatch g4228 (.Q(w3561), .D(S[1]), .C(w3531), .nC(w3592) );
	vdp_slatch g4229 (.Q(w3559), .D(S[0]), .C(w3531), .nC(w3592) );
	vdp_slatch g4230 (.Q(w3556), .D(S[7]), .C(w3532), .nC(w3593) );
	vdp_slatch g4231 (.Q(w3557), .D(S[6]), .C(w3532), .nC(w3593) );
	vdp_slatch g4232 (.Q(w3555), .D(S[5]), .C(w3532), .nC(w3593) );
	vdp_slatch g4233 (.Q(w3554), .D(S[4]), .C(w3532), .nC(w3593) );
	vdp_slatch g4234 (.Q(w3552), .D(S[3]), .C(w3532), .nC(w3593) );
	vdp_slatch g4235 (.Q(w3550), .D(S[2]), .C(w3532), .nC(w3593) );
	vdp_slatch g4236 (.Q(w3548), .D(S[1]), .C(w3532), .nC(w3593) );
	vdp_slatch g4237 (.Q(w3545), .D(S[0]), .C(w3532), .nC(w3593) );
	vdp_sr_bit g4238 (.Q(w4114), .D(w3526), .C1(HCLK2), .C2(HCLK1), .nC2(nHCLK1), .nC1(nHCLK2) );
	vdp_sr_bit g4239 (.Q(w3533), .D(w4082), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and g4240 (.Z(w4082), .A(w14), .B(M5) );
	vdp_not g4241 (.nZ(w4080), .A(w3533) );
	vdp_aon22 g4242 (.Z(w3097), .A1(w4085), .B1(w3597), .A2(w3596), .B2(w4042) );
	vdp_aon22 g4243 (.Z(w3094), .A1(w4084), .B1(1'b0), .A2(w3596), .B2(w4042) );
	vdp_aon22 g4244 (.Z(w3595), .A1(w3597), .B1(w3563), .A2(w3596), .B2(w4042) );
	vdp_aon22 g4245 (.Z(w3067), .A1(w3598), .B1(w3561), .A2(w3596), .B2(w4042) );
	vdp_aon22 g4246 (.Z(w3070), .A1(w4083), .B1(w3598), .A2(w3596), .B2(w4042) );
	vdp_comp_strong g4247 (.Z(w3532), .nZ(w3593), .A(w3283) );
	vdp_comp_we g4248 (.Z(w3596), .nZ(w4042), .A(M5) );
	vdp_aon22 g4249 (.Z(w3537), .A1(w3594), .B1(w3595), .A2(w3533), .B2(w4080) );
	vdp_sr_bit g4250 (.Q(w3992), .D(FIFOo[0]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4251 (.Q(w3996), .D(FIFOo[1]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4252 (.Q(w3994), .D(FIFOo[2]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4253 (.Q(w3993), .D(FIFOo[3]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4254 (.Q(w3981), .D(FIFOo[4]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4255 (.Q(w3979), .D(FIFOo[5]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4256 (.Q(w3986), .D(FIFOo[6]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4257 (.Q(w3988), .D(FIFOo[7]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_aon22 g4258 (.Z(w1401), .B1(w4463), .A1(w1429), .B2(w4481), .A2(w43) );
	vdp_not g4259 (.nZ(w4481), .A(w43) );
	vdp_not g4260 (.nZ(w4453), .A(w4440) );
	vdp_not g4261 (.nZ(w4452), .A(w4453) );
	vdp_not g4262 (.nZ(w4451), .A(w4452) );
	vdp_not g4263 (.nZ(w4450), .A(w4451) );
	vdp_and g4264 (.Z(w4463), .B(w4454), .A(w4458) );
	vdp_not g4265 (.nZ(w4454), .A(w4457) );
	vdp_not g4266 (.nZ(w4457), .A(w4456) );
	vdp_not g4267 (.nZ(w4456), .A(w4455) );
	vdp_not g4268 (.nZ(w4455), .A(w4458) );
	vdp_or g4269 (.Z(w4458), .B(w4438), .A(w4437) );
	vdp_dff g4270 (.Q(w4438), .R(w4427), .D(w4437), .C(w4436) );
	vdp_not g4271 (.nZ(w4436), .A(w4459) );
	vdp_nor g4272 (.Z(w4435), .B(w4460), .A(w4437) );
	vdp_dff g4273 (.Q(w4437), .R(w4427), .D(w4460), .C(w4459) );
	vdp_dff g4274 (.Q(w4460), .R(w4427), .D(w4435), .C(w4459) );
	vdp_not g4275 (.nZ(w4459), .A(w4446) );
	vdp_not g4276 (.nZ(w4433), .A(w4446) );
	vdp_dff g4277 (.Q(w4430), .R(w4427), .D(w4461), .C(w4429) );
	vdp_dff g4278 (.Q(w4461), .R(w4427), .D(w4428), .C(w4426) );
	vdp_not g4279 (.nZ(w4426), .A(w4469) );
	vdp_dff g4280 (.Q(w4428), .R(w4427), .D(w4447), .C(w4426) );
	vdp_not g4281 (.nZ(w4429), .A(w4426) );
	vdp_nor g4282 (.Z(w4488), .B(w4464), .A(w4465) );
	vdp_nor g4283 (.Z(w4466), .B(w4464), .A(H40) );
	vdp_not g4284 (.nZ(w4465), .A(H40) );
	vdp_not g4285 (.nZ(w4441), .A(PAL) );
	vdp_AOI222 g4286 (.Z(w4434), .B1(w4468), .A1(w4467), .B2(w4488), .A2(w4464), .C1(w4433), .C2(w4466) );
	vdp_not g4287 (.nZ(EDCLK_O), .A(w4434) );
	vdp_or g4288 (.Z(w4462), .B(w4430), .A(w4461) );
	vdp_nor g4289 (.Z(w4447), .B(w4428), .A(w4461) );
	vdp_not g4290 (.nZ(w4423), .A(w4487) );
	vdp_nand g4291 (.Z(w4442), .B(w4423), .A(w4422) );
	vdp_sr_bit g4292 (.Q(w4487), .D(w4422), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_not g4293 (.nZ(w4486), .A(w4472) );
	vdp_not g4294 (.nZ(w1161), .A(w4485) );
	vdp_not g4295 (.nZ(SYSRES), .A(w4486) );
	vdp_comp_dff g4296 (.Q(w4422), .D(w4472), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_not g4297 (.nZ(w4482), .A(w4483) );
	vdp_not g4298 (.nZ(w4427), .A(w4484) );
	vdp_not g4299 (.nZ(w4471), .A(w4470) );
	vdp_nand g4300 (.Z(w4484), .B(w4471), .A(w4425) );
	vdp_not g4301 (.nZ(w4469), .A(w4473) );
	vdp_nand g4302 (.Z(w4476), .B(w4475), .A(w4474) );
	vdp_not g4303 (.nZ(w4446), .A(w4431) );
	vdp_nand g4304 (.Z(w4479), .B(w4478), .A(w4477) );
	vdp_not g4305 (.nZ(w4440), .A(w4445) );
	vdp_not g4306 (.nZ(RES), .A(w4442) );
	vdp_dff g4307 (.Q(w4425), .R(1'b0), .D(w4472), .C(w4443) );
	vdp_dff g4308 (.Q(w4470), .R(1'b0), .D(w4425), .C(w4443) );
	vdp_dff g4309 (.Q(w4483), .R(w4427), .D(w4473), .C(w4443) );
	vdp_dff g4310 (.Q(w4473), .R(w4427), .D(w4482), .C(w4443) );
	vdp_dff g4311 (.Q(w4474), .R(w4427), .D(w4431), .C(w4443) );
	vdp_dff g4312 (.Q(w4475), .R(w4427), .D(w4474), .C(w4443) );
	vdp_dff g4313 (.Q(w4431), .R(w4427), .D(w4476), .C(w4443) );
	vdp_dff g4314 (.Q(w4477), .R(w4427), .D(w4445), .C(w4443) );
	vdp_dff g4315 (.Q(w4478), .R(w4427), .D(w4477), .C(w4443) );
	vdp_dff g4316 (.Q(w4480), .R(w4427), .D(w4479), .C(w4443) );
	vdp_dff g4317 (.Q(w4445), .R(w4427), .D(w4480), .C(w4443) );
	vdp_not g4318 (.nZ(w4468), .A(w4469) );
	vdp_nand g4319 (.Z(w4472), .B(w1430), .A(w4485) );
	vdp_not g4320 (.nZ(68K CPU CLOCK), .A(w4439) );
	vdp_or g4321 (.Z(w4464), .B(w43), .A(w1142) );
	vdp_aon22 g4322 (.Z(w4432), .B1(w4462), .A1(w4463), .B2(PAL), .A2(w4441) );
	vdp_or g4323 (.Z(w4439), .B(w4450), .A(w4440) );
	vdp_comp_we g4324 (.A(w2627), .nZ(nHCLK2), .Z(HCLK2) );
	vdp_comp_we g4325 (.A(w2626), .nZ(nHCLK1), .Z(HCLK1) );
	vdp_comp_we g4326 (.A(w4496), .nZ(nDCLK2), .Z(DCLK2) );
	vdp_comp_we g4327 (.A(EDCLK_O), .nZ(nDCLK1), .Z(DCLK1) );
	vdp_not g4328 (.nZ(w4496), .A(EDCLK_O) );
	vdp_sr_bit g4329 (.Q(w4591), .D(w4590), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4330 (.Q(w4609), .D(w4586), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4331 (.Q(w4586), .D(w4571), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4332 (.Q(w4571), .D(w4563), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4333 (.Q(w4566), .D(w6526), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4334 (.Q(w6526), .D(w6527), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4335 (.Q(w6527), .D(w6529), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4336 (.Q(w6529), .D(w6528), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4337 (.Q(w6528), .D(w6530), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4338 (.Q(w6530), .D(w6531), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4339 (.Q(w6531), .D(w6533), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4340 (.Q(w6533), .D(w6532), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4341 (.Q(w6532), .D(w6358), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4342 (.Q(w6358), .D(w4511), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4343 (.Q(w4547), .D(w4548), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4344 (.Q(w4548), .D(w24), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4345 (.Q(w4812), .D(w6534), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4346 (.Q(w4516), .D(w4846), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4347 (.Q(w4515), .D(w6522), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4348 (.Q(w6220), .D(w4593), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4349 (.Q(w4592), .D(w6535), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4350 (.Q(w4594), .D(w4584), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4351 (.Q(w6524), .D(w4), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4352 (.Q(w4535), .D(w4556), .nC(w4559), .C(w4560) );
	vdp_slatch g4353 (.Q(w4540), .D(w4557), .nC(w4559), .C(w4560) );
	vdp_slatch g4354 (.Q(w4527), .D(w4558), .nC(w4559), .C(w4560) );
	vdp_slatch g4355 (.Q(w4519), .D(w4564), .nC(w4559), .C(w4560) );
	vdp_slatch g4356 (.Q(w4518), .D(w4555), .nC(w4559), .C(w4560) );
	vdp_slatch g4357 (.Q(w4517), .D(w4554), .nC(w4559), .C(w4560) );
	vdp_slatch g4358 (.Q(w4568), .D(w4553), .nC(w4559), .C(w4560) );
	vdp_slatch g4359 (.Q(w4520), .D(w4551), .nC(w4559), .C(w4560) );
	vdp_slatch g4360 (.Q(w4523), .D(w4552), .nC(w4559), .C(w4560) );
	vdp_slatch g4361 (.Q(w4524), .D(w4550), .nC(w4559), .C(w4560) );
	vdp_comp_str g4362 (.nZ(w4559), .A(w4565), .Z(w4560) );
	vdp_sr_bit g4363 (.Q(w4587), .D(w4610), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4364 (.Q(w6206), .D(w7), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_xor g4365 (.Z(w4533), .B(w4525), .A(w4536) );
	vdp_xor g4366 (.Z(w4528), .B(w4526), .A(w4534) );
	vdp_xor g4367 (.Z(w4530), .B(w4513), .A(w4527) );
	vdp_xor g4368 (.Z(w6309), .B(w4513), .A(w4519) );
	vdp_xor g4369 (.Z(w6310), .B(w4513), .A(w4518) );
	vdp_xor g4370 (.Z(w6305), .B(w4513), .A(w4517) );
	vdp_aon22 g4371 (.Z(w6306), .B2(w4541), .B1(w4535), .A1(w4533), .A2(w4529) );
	vdp_aon22 g4372 (.Z(w6307), .B2(w4541), .B1(w4533), .A1(w4528), .A2(w4529) );
	vdp_aon22 g4373 (.Z(w6308), .B2(w4541), .B1(w4528), .A1(w4530), .A2(w4529) );
	vdp_aon22 g4374 (.Z(w4531), .B2(w4522), .B1(w4527), .A1(w4540), .A2(w4532) );
	vdp_aon22 g4375 (.Z(w4537), .B2(w4522), .B1(w4540), .A1(w4535), .A2(w4532) );
	vdp_aon22 g4376 (.Z(w4602), .B2(w4595), .B1(w4598), .A1(w4599), .A2(w79) );
	vdp_aon22 g4377 (.Z(w4603), .B2(w4597), .B1(w4598), .A1(w4599), .A2(w78) );
	vdp_aon22 g4378 (.Z(w4604), .B2(w4596), .B1(w4598), .A1(w4599), .A2(w77) );
	vdp_aon22 g4379 (.Z(w4605), .B2(w4600), .B1(w4598), .A1(w4599), .A2(w76) );
	vdp_aon22 g4380 (.Z(w4606), .B2(w4601), .B1(w4598), .A1(w4599), .A2(w75) );
	vdp_not g4381 (.nZ(w4572), .A(w4511) );
	vdp_not g4382 (.nZ(w4544), .A(w4576) );
	vdp_not g4383 (.nZ(w4575), .A(w120) );
	vdp_not g4384 (.nZ(w4580), .A(w4578) );
	vdp_not g4385 (.nZ(w4567), .A(M5) );
	vdp_not g4386 (.nZ(w4608), .A(w80) );
	vdp_not g4387 (.nZ(w4607), .A(w81) );
	vdp_not g4388 (.nZ(w4582), .A(1'b0) );
	vdp_not g4389 (.nZ(w4583), .A(M5) );
	vdp_not g4390 (.nZ(w4510), .A(w4511) );
	vdp_not g4391 (.nZ(w4514), .A(w4545) );
	vdp_not g4392 (.nZ(w4521), .A(w4524) );
	vdp_not g4393 (.nZ(w4526), .A(w4562) );
	vdp_and g4394 (.Z(w4563), .B(w4572), .A(w4573) );
	vdp_and g4395 (.Z(w4577), .B(w4575), .A(w4586) );
	vdp_or g4396 (.Z(w4574), .B(w4577), .A(w4589) );
	vdp_or g4397 (.Z(w4570), .B(w4612), .A(w4577) );
	vdp_and g4398 (.Z(w4588), .B(w4581), .A(1'b0) );
	vdp_and g4399 (.Z(w4611), .B(w4581), .A(w4582) );
	vdp_or g4400 (.Z(w4610), .B(w7), .A(w27) );
	vdp_and g4401 (.Z(w122), .B(w6668), .A(w4) );
	vdp_and g4402 (.Z(w6522), .B(w4510), .A(w4512) );
	vdp_or g4403 (.Z(w4561), .B(w4516), .A(w4515) );
	vdp_and g4404 (.Z(w4525), .B(w4520), .A(w4513) );
	vdp_comp_we g4405 (.nZ(w4522), .A(w1), .Z(w4532) );
	vdp_comp_we g4406 (.nZ(w4541), .A(w1), .Z(w4529) );
	vdp_comp_we g4407 (.nZ(w4598), .A(w120), .Z(w4599) );
	vdp_not g4408 (.nZ(w4620), .A(w4590) );
	vdp_rs_ff g4409 (.Q(w6523), .R(w6524), .S(w4561) );
	vdp_rs_ff g4410 (.Q(w6668), .R(w6524), .S(w4515) );
	vdp_ha g4411 (.SUM(w4536), .B(w4537), .A(w4538) );
	vdp_ha g4412 (.SUM(w4534), .B(w4531), .A(w4539), .CO(w4538) );
	vdp_not g4413 (.nZ(w4546), .A(w4509) );
	vdp_and g4414 (.Z(w4549), .B(w4511), .A(w4512) );
	vdp_and3 g4415 (.Z(w4539), .B(w4520), .A(w4513), .C(w4521) );
	vdp_and3 g4416 (.Z(w4593), .B(w4591), .A(M5), .C(w4620) );
	vdp_and3 g4417 (.Z(w6535), .B(w4596), .A(w4595), .C(w4594) );
	vdp_and3 g4418 (.Z(w4612), .B(w81), .A(w4608), .C(w113) );
	vdp_and3 g4419 (.Z(w6525), .B(w80), .A(w4607), .C(w113) );
	vdp_and3 g4420 (.Z(w4589), .B(w4608), .A(w4607), .C(w113) );
	vdp_or3 g4421 (.Z(w4569), .B(w6525), .A(w4577), .C(w4580) );
	vdp_and3 g4422 (.Z(w4565), .B(HCLK1), .A(w4547), .C(DCLK1) );
	vdp_or3 g4423 (.Z(w4581), .B(w4584), .A(w4609), .C(w4583) );
	vdp_oai21 g4424 (.Z(w4562), .B(w4513), .A1(w4520), .A2(w4524) );
	vdp_nor g4425 (.Z(w4509), .B(w4549), .A(w4548) );
	vdp_nor g4426 (.Z(w6534), .B(w4514), .A(w6523) );
	vdp_nand g4427 (.Z(w4585), .B(w4567), .A(w4566) );
	vdp_nand g4428 (.Z(w4543), .B(w4608), .A(w4607) );
	vdp_nand g4429 (.Z(w4576), .B(w80), .A(w4607) );
	vdp_nand g4430 (.Z(w4542), .B(w81), .A(w4608) );
	vdp_nor g4431 (.Z(w4590), .B(w4592), .A(w4507) );
	vdp_cnt_bit_rev g4432 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4595), .CI(w4624), .B(w4587), .A(w4588) );
	vdp_cnt_bit_rev g4433 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4597), .CI(w4623), .B(w4587), .A(w4588), .CO(w4624) );
	vdp_cnt_bit_rev g4434 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4596), .CI(w4622), .B(w4587), .A(w4588), .CO(w4623) );
	vdp_cnt_bit_rev g4435 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4600), .CI(w4621), .B(w4587), .A(w4588), .CO(w4622) );
	vdp_cnt_bit_rev g4436 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4601), .CI(w4611), .B(w4587), .A(w4588), .CO(w4621) );
	vdp_cnt_bit_load g4437 (.Q(w4631), .D(w4671), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4633), .CI(w6571), .L(w4672), .nL(w4637) );
	vdp_cnt_bit_load g4438 (.Q(w4634), .D(w4676), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4633), .CI(w6570), .L(w4672), .nL(w4637), .CO(w6571) );
	vdp_cnt_bit_load g4439 (.Q(w4636), .D(w4677), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4633), .CI(w6569), .L(w4672), .nL(w4637), .CO(w6570) );
	vdp_cnt_bit_load g4440 (.Q(w4638), .D(w4701), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4633), .CI(w6568), .L(w4672), .nL(w4637), .CO(w6569) );
	vdp_cnt_bit_load g4441 (.Q(w4642), .D(w4702), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4633), .CI(w6567), .L(w4672), .nL(w4637), .CO(w6568) );
	vdp_cnt_bit_load g4442 (.Q(w4639), .D(w4703), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4633), .CI(w6566), .L(w4672), .nL(w4637), .CO(w6567) );
	vdp_cnt_bit_load g4443 (.Q(w4635), .D(w4704), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4633), .CI(w4632), .L(w4672), .nL(w4637), .CO(w6566) );
	vdp_fa g4444 (.SUM(w4779), .CO(w6581), .CI(1'b1), .A(w4834), .B(w4782) );
	vdp_fa g4445 (.SUM(w4781), .CO(w6582), .CI(w6581), .A(w4833), .B(w4786) );
	vdp_fa g4446 (.SUM(w4787), .CO(w6583), .CI(w6582), .A(w4832), .B(w4790) );
	vdp_fa g4447 (.SUM(w4789), .CO(w6584), .CI(w6583), .A(w4831), .B(w4792) );
	vdp_fa g4448 (.SUM(w4794), .CO(w6585), .CI(w6584), .A(w4830), .B(w4796) );
	vdp_fa g4449 (.SUM(w4800), .CO(w6586), .CI(w6585), .A(w4829), .B(w4825) );
	vdp_fa g4450 (.SUM(w4803), .CO(w6587), .CI(w6586), .A(w4827), .B(w4802) );
	vdp_fa g4451 (.SUM(w4807), .CO(w6588), .CI(w6587), .A(w4839), .B(w4806) );
	vdp_fa g4452 (.SUM(w4809), .CO(w6589), .CI(w6588), .A(w4840), .B(w4808) );
	vdp_fa g4453 (.SUM(w4823), .CI(w6589), .A(w4844), .B(w4822) );
	vdp_fa g4454 (.SUM(w4834), .CO(w6572), .CI(1'b0), .A(VPOS[0]), .B(w4835) );
	vdp_fa g4455 (.SUM(w4833), .CO(w6573), .CI(w6572), .A(VPOS[1]), .B(w1) );
	vdp_fa g4456 (.SUM(w4832), .CO(w6574), .CI(w6573), .A(VPOS[2]), .B(1'b0) );
	vdp_fa g4457 (.SUM(w4831), .CO(w6575), .CI(w6574), .A(VPOS[3]), .B(1'b0) );
	vdp_fa g4458 (.SUM(w4830), .CO(w6576), .CI(w6575), .A(VPOS[4]), .B(1'b0) );
	vdp_fa g4459 (.SUM(w4829), .CO(w6577), .CI(w6576), .A(VPOS[5]), .B(1'b0) );
	vdp_fa g4460 (.SUM(w4827), .CO(w6578), .CI(w6577), .A(VPOS[6]), .B(1'b0) );
	vdp_fa g4461 (.SUM(w4839), .CO(w6579), .CI(w6578), .A(VPOS[7]), .B(w4835) );
	vdp_fa g4462 (.SUM(w4840), .CO(w6580), .CI(w6579), .A(VPOS[8]), .B(w1) );
	vdp_fa g4463 (.SUM(w4844), .CI(w6580), .A(VPOS[9]), .B(1'b0) );
	vdp_slatch g4464 (.nC(w4727), .C(w4726), .Q(w4773), .D(S[0]) );
	vdp_dlatch_inv g4465 (.nQ(w4772), .D(w4740), .nC(nHCLK2), .C(HCLK2) );
	vdp_slatch g4466 (.nC(w4712), .C(w4711), .Q(w4740), .D(w4729) );
	vdp_slatch g4467 (.nC(w4727), .C(w4726), .Q(w4770), .D(S[1]) );
	vdp_slatch g4468 (.nC(w4712), .C(w4711), .Q(w6611), .D(w4731) );
	vdp_slatch g4469 (.nC(w4727), .C(w4726), .Q(w4768), .D(S[2]) );
	vdp_slatch g4470 (.nC(w4712), .C(w4711), .Q(w6612), .D(w4722) );
	vdp_slatch g4471 (.nC(w4727), .C(w4726), .Q(w4766), .D(S[3]) );
	vdp_slatch g4472 (.nC(w4712), .C(w4711), .Q(w6613), .D(w4718) );
	vdp_slatch g4473 (.nC(w4727), .C(w4726), .Q(w4762), .D(S[4]) );
	vdp_slatch g4474 (.nC(w4712), .C(w4711), .Q(w6614), .D(w4714) );
	vdp_slatch g4475 (.nC(w4727), .C(w4726), .Q(w4761), .D(S[5]) );
	vdp_slatch g4476 (.nC(w4712), .C(w4711), .Q(w6615), .D(w4710) );
	vdp_slatch g4477 (.nC(w4727), .C(w4726), .Q(w4758), .D(S[6]) );
	vdp_slatch g4478 (.nC(w4712), .C(w4711), .Q(w6616), .D(w6558) );
	vdp_slatch g4479 (.nC(w4727), .C(w4726), .Q(w6617), .D(S[7]) );
	vdp_slatch g4480 (.nC(w4712), .C(w4711), .Q(w6618), .D(w4742) );
	vdp_slatch g4481 (.nC(w4712), .C(w4711), .Q(w4743), .D(w4744) );
	vdp_slatch g4482 (.nC(w4712), .C(w4711), .Q(w6619), .D(w4746) );
	vdp_dlatch_inv g4483 (.nQ(w4769), .D(w6611), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4484 (.nQ(w4767), .D(w6612), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4485 (.nQ(w4764), .D(w6613), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4486 (.nQ(w4763), .D(w6614), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4487 (.nQ(w4760), .D(w6615), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4488 (.nQ(w4757), .D(w6616), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4489 (.nQ(w4756), .D(w6618), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4490 (.nQ(w4755), .D(w4743), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4491 (.nQ(w4745), .D(w6619), .nC(nHCLK2), .C(HCLK2) );
	vdp_sr_bit g4492 (.Q(w4697), .D(w4628), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4493 (.Z(w4545), .B2(w4693), .B1(w4699), .A1(M5), .A2(w4698) );
	vdp_sr_bit g4494 (.Q(w4628), .D(w4694), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4495 (.Q(w4694), .D(w4695), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4496 (.Q(w4695), .D(w4673), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4497 (.Q(w4734), .D(w4736), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4498 (.Q(w4725), .D(w4739), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4499 (.Q(w4721), .D(w4732), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4500 (.Q(w4717), .D(w4733), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4501 (.Q(w4713), .D(w4715), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4502 (.Q(w4709), .D(w4707), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4503 (.Q(w4741), .D(w4708), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4504 (.Q(w6620), .D(w4706), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4505 (.Q(w4655), .D(w4705), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4506 (.Q(w4662), .D(w4700), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4507 (.Q(w4696), .D(w4629), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4508 (.Q(w4629), .D(w4651), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4509 (.Q(w4881), .D(w126), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4510 (.Q(w4883), .D(VRAMA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4511 (.Q(w4651), .D(w9), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4512 (.Q(w4884), .D(w6565), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4513 (.Q(w6565), .D(w4881), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4514 (.Q(w6609), .D(w4867), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4515 (.Q(w6607), .D(w4870), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4516 (.Q(w6605), .D(w4885), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4517 (.Q(w6603), .D(w4847), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4518 (.Q(w6601), .D(w4671), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4519 (.Q(w6599), .D(w4676), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4520 (.Q(w6597), .D(w4677), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4521 (.Q(w6595), .D(w4701), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4522 (.Q(w6593), .D(w4702), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4523 (.Q(w6591), .D(w4703), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4524 (.Q(w4865), .D(w4704), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4525 (.Q(w4857), .D(w6590), .nC(w4856), .C(w4848) );
	vdp_dlatch_inv g4526 (.nQ(w6590), .D(w4865), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4527 (.Q(w4858), .D(w6592), .nC(w4856), .C(w4848) );
	vdp_dlatch_inv g4528 (.nQ(w6592), .D(w6591), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4529 (.Q(w4859), .D(w6594), .nC(w4856), .C(w4848) );
	vdp_dlatch_inv g4530 (.nQ(w6594), .D(w6593), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4531 (.Q(w4860), .D(w6596), .nC(w4856), .C(w4848) );
	vdp_dlatch_inv g4532 (.nQ(w6596), .D(w6595), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4533 (.Q(w4861), .D(w6598), .nC(w4856), .C(w4848) );
	vdp_dlatch_inv g4534 (.nQ(w6598), .D(w6597), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4535 (.Q(w6564), .D(w6600), .nC(w4856), .C(w4848) );
	vdp_dlatch_inv g4536 (.nQ(w6600), .D(w6599), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4537 (.Q(w4862), .D(w6602), .nC(w4856), .C(w4848) );
	vdp_dlatch_inv g4538 (.nQ(w6602), .D(w6601), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4539 (.Q(w4852), .D(w6604), .nC(w4856), .C(w4848) );
	vdp_dlatch_inv g4540 (.nQ(w6604), .D(w6603), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4541 (.Q(w4855), .D(w6606), .nC(w4856), .C(w4848) );
	vdp_dlatch_inv g4542 (.nQ(w6606), .D(w6605), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4543 (.Q(w4853), .D(w6608), .nC(w4856), .C(w4848) );
	vdp_dlatch_inv g4544 (.nQ(w6608), .D(w6607), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4545 (.Q(w4854), .D(w6610), .nC(w4856), .C(w4848) );
	vdp_dlatch_inv g4546 (.nQ(w6610), .D(w6609), .nC(nHCLK1), .C(HCLK1) );
	vdp_aon22 g4547 (.Z(w6377), .B2(w4681), .B1(w4631), .A1(w4630), .A2(w6356) );
	vdp_aon22 g4548 (.Z(w6378), .B2(w4681), .B1(w4634), .A1(w4630), .A2(w4686) );
	vdp_aon22 g4549 (.Z(w6379), .B2(w4681), .B1(w4636), .A1(w4630), .A2(w4685) );
	vdp_aon22 g4550 (.Z(w6380), .B2(w4681), .B1(w4638), .A1(w4630), .A2(w4684) );
	vdp_aon22 g4551 (.Z(w6381), .B2(w4681), .B1(w4642), .A1(w4630), .A2(w4683) );
	vdp_aon22 g4552 (.Z(w6383), .B2(w4681), .B1(w4639), .A1(w4630), .A2(w4682) );
	vdp_aon22 g4553 (.Z(w6382), .B2(w4681), .B1(w4635), .A1(w4630), .A2(w4680) );
	vdp_aon22 g4554 (.Z(w4906), .B2(w4644), .B1(w3), .A1(w4640), .A2(w4635) );
	vdp_aon22 g4555 (.Z(w4793), .B2(w4753), .B1(w4762), .A1(w4763), .A2(w4777) );
	vdp_2x_sr_bit g4556 (.Q(w4692), .D(w4635), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4557 (.Z(w6357), .B2(w4644), .B1(w4692), .A1(w4640), .A2(w4639) );
	vdp_2x_sr_bit g4558 (.Q(w4641), .D(w4639), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4559 (.Z(w4961), .B2(w4644), .B1(w4641), .A1(w4640), .A2(w4642) );
	vdp_2x_sr_bit g4560 (.Q(w4679), .D(w4642), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4561 (.Z(w4967), .B2(w4644), .B1(w4679), .A1(w4640), .A2(w4638) );
	vdp_2x_sr_bit g4562 (.Q(w4643), .D(w4638), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4563 (.Z(w5017), .B2(w4644), .B1(w4643), .A1(w4640), .A2(w4636) );
	vdp_2x_sr_bit g4564 (.Q(w4646), .D(w4636), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4565 (.Z(w5069), .B2(w4644), .B1(w4646), .A1(w4640), .A2(w4634) );
	vdp_aon22 g4566 (.Z(w5084), .B2(w4644), .B1(1'b1), .A1(w4640), .A2(w4631) );
	vdp_aon22 g4567 (.Z(w4729), .B2(w4654), .B1(w4730), .A1(w4657), .A2(w4728) );
	vdp_dlatch_inv g4568 (.nQ(w4728), .D(w4734), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4569 (.nZ(w4730), .A(S[0]) );
	vdp_aon22 g4570 (.Z(w4731), .B2(w4654), .B1(w4724), .A1(w4657), .A2(w4723) );
	vdp_dlatch_inv g4571 (.nQ(w4723), .D(w4725), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4572 (.nZ(w4724), .A(S[1]) );
	vdp_aon22 g4573 (.Z(w4722), .B2(w4654), .B1(w4720), .A1(w4657), .A2(w4719) );
	vdp_dlatch_inv g4574 (.nQ(w4719), .D(w4721), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4575 (.nZ(w4720), .A(S[2]) );
	vdp_aon22 g4576 (.Z(w4718), .B2(w4654), .B1(w4678), .A1(w4657), .A2(w4716) );
	vdp_dlatch_inv g4577 (.nQ(w4716), .D(w4717), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4578 (.nZ(w4678), .A(S[3]) );
	vdp_aon22 g4579 (.Z(w4714), .B2(w4654), .B1(w4674), .A1(w4657), .A2(w4675) );
	vdp_dlatch_inv g4580 (.nQ(w4675), .D(w4713), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4581 (.nZ(w4674), .A(S[4]) );
	vdp_aon22 g4582 (.Z(w4710), .B2(w4654), .B1(w4670), .A1(w4657), .A2(w4669) );
	vdp_dlatch_inv g4583 (.nQ(w4669), .D(w4709), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4584 (.nZ(w4670), .A(S[5]) );
	vdp_aon22 g4585 (.Z(w6558), .B2(w4654), .B1(w4665), .A1(w4657), .A2(w4664) );
	vdp_dlatch_inv g4586 (.nQ(w4664), .D(w4741), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4587 (.nZ(w4665), .A(S[6]) );
	vdp_aon22 g4588 (.Z(w4742), .B2(w4654), .B1(w4658), .A1(w4657), .A2(w4656) );
	vdp_dlatch_inv g4589 (.nQ(w4656), .D(w6620), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4590 (.nZ(w4658), .A(S[7]) );
	vdp_aon22 g4591 (.Z(w4744), .B2(w4654), .B1(w4901), .A1(w4657), .A2(1'b1) );
	vdp_dlatch_inv g4592 (.nQ(w4901), .D(w4655), .nC(nHCLK1), .C(HCLK1) );
	vdp_aon22 g4593 (.Z(w4746), .B2(w4654), .B1(1'b1), .A1(w4657), .A2(w4663) );
	vdp_dlatch_inv g4594 (.nQ(w4663), .D(w4662), .nC(nHCLK1), .C(HCLK1) );
	vdp_sr_bit g4595 (.Q(w4633), .D(w6552), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4596 (.Q(w4645), .D(w30), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4597 (.Q(w4666), .D(w4645), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4598 (.Q(w4650), .D(w5), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4599 (.Q(w4660), .D(w4650), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4600 (.Q(w4673), .D(w6551), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_not g4601 (.nZ(w4668), .A(w4667) );
	vdp_not g4602 (.nZ(w4661), .A(M5) );
	vdp_not g4603 (.nZ(w6552), .A(w4659) );
	vdp_not g4604 (.nZ(w4649), .A(w4660) );
	vdp_not g4605 (.nZ(w6551), .A(w4652) );
	vdp_not g4606 (.nZ(w4647), .A(w4632) );
	vdp_aon22 g4607 (.Z(w4752), .B2(w4748), .B1(w4558), .A1(w4747), .A2(w4557) );
	vdp_aon22 g4608 (.Z(w4751), .B2(w4748), .B1(w4557), .A1(w4747), .A2(w4556) );
	vdp_aon22 g4609 (.Z(w4750), .B2(w4748), .B1(w4556), .A1(w4747), .A2(1'b0) );
	vdp_slatch g4610 (.nQ(w6629), .D(w4880), .nC(w4864), .C(w4869) );
	vdp_aon22 g4611 (.Z(w4880), .B2(w4863), .B1(w4736), .A1(w4868), .A2(w4704) );
	vdp_notif0 g4612 (.A(w6629), .nZ(AD_DATA[0]), .nE(w4874) );
	vdp_slatch g4613 (.nQ(w6628), .D(w4879), .nC(w4864), .C(w4869) );
	vdp_aon22 g4614 (.Z(w4879), .B2(w4863), .B1(w4739), .A1(w4868), .A2(w4703) );
	vdp_notif0 g4615 (.A(w6628), .nZ(AD_DATA[1]), .nE(w4874) );
	vdp_slatch g4616 (.nQ(w6627), .D(w4878), .nC(w4864), .C(w4869) );
	vdp_aon22 g4617 (.Z(w4878), .B2(w4863), .B1(w4732), .A1(w4868), .A2(w4702) );
	vdp_notif0 g4618 (.A(w6627), .nZ(AD_DATA[2]), .nE(w4874) );
	vdp_slatch g4619 (.nQ(w6626), .D(w6562), .nC(w4864), .C(w4869) );
	vdp_aon22 g4620 (.Z(w6562), .B2(w4863), .B1(w4733), .A1(w4868), .A2(w4701) );
	vdp_notif0 g4621 (.A(w6626), .nZ(AD_DATA[3]), .nE(w4874) );
	vdp_slatch g4622 (.nQ(w6625), .D(w6561), .nC(w4864), .C(w4869) );
	vdp_aon22 g4623 (.Z(w6561), .B2(w4863), .B1(w4715), .A1(w4868), .A2(w4677) );
	vdp_notif0 g4624 (.A(w6625), .nZ(AD_DATA[4]), .nE(w4874) );
	vdp_slatch g4625 (.nQ(w6624), .D(w6560), .nC(w4864), .C(w4869) );
	vdp_aon22 g4626 (.Z(w6560), .B2(w4863), .B1(w4707), .A1(w4868), .A2(w4676) );
	vdp_notif0 g4627 (.A(w6624), .nZ(AD_DATA[5]), .nE(w4874) );
	vdp_slatch g4628 (.nQ(w6623), .D(w4877), .nC(w4864), .C(w4869) );
	vdp_aon22 g4629 (.Z(w4877), .B2(w4863), .B1(w4708), .A1(w4868), .A2(w4671) );
	vdp_notif0 g4630 (.A(w6623), .nZ(AD_DATA[6]), .nE(w4874) );
	vdp_slatch g4631 (.nQ(w6622), .D(w4886), .nC(w4864), .C(w4869) );
	vdp_aon22 g4632 (.Z(w4886), .B2(w4863), .B1(w4706), .A1(w4868), .A2(w4847) );
	vdp_notif0 g4633 (.A(w6622), .nZ(AD_DATA[7]), .nE(w4874) );
	vdp_slatch g4634 (.nQ(w4876), .D(w4875), .nC(w4864), .C(w4869) );
	vdp_aon22 g4635 (.Z(w4875), .B2(w4863), .B1(w4705), .A1(w4868), .A2(w4885) );
	vdp_notif0 g4636 (.A(w4876), .nZ(RD_DATA[0]), .nE(w4874) );
	vdp_slatch g4637 (.nQ(w4873), .D(w4872), .nC(w4864), .C(w4869) );
	vdp_aon22 g4638 (.Z(w4872), .B2(w4863), .B1(w4700), .A1(w4868), .A2(w4870) );
	vdp_notif0 g4639 (.A(w4873), .nZ(RD_DATA[1]), .nE(w4874) );
	vdp_slatch g4640 (.nQ(w4871), .D(w4866), .nC(w4864), .C(w4869) );
	vdp_aon22 g4641 (.Z(w4866), .B2(w4863), .B1(1'b0), .A1(w4868), .A2(w4867) );
	vdp_notif0 g4642 (.A(w4871), .nZ(RD_DATA[2]), .nE(w4874) );
	vdp_not g4643 (.nZ(w4874), .A(w4884) );
	vdp_sr_bit g4644 (.Q(w4551), .D(w6633), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4645 (.Q(w4552), .D(w4842), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4646 (.Q(w4838), .D(w4836), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_dlatch_inv g4647 (.nQ(w4837), .D(w4738), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4648 (.nQ(w4836), .D(w4776), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g4649 (.nQ(w4782), .D(w4778), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4650 (.nQ(w6559), .D(w4779), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4651 (.nQ(w4786), .D(w4780), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4652 (.nQ(w4784), .D(w4781), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4653 (.nQ(w4790), .D(w4785), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4654 (.nQ(w4788), .D(w4787), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4655 (.nQ(w4792), .D(w4791), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4656 (.nQ(w4801), .D(w4789), .nC(nHCLK2), .C(HCLK2) );
	vdp_aon22 g4657 (.Z(w4791), .B2(w4753), .B1(w4766), .A1(w4764), .A2(w4777) );
	vdp_aon22 g4658 (.Z(w4785), .B2(w4753), .B1(w4768), .A1(w4767), .A2(w4777) );
	vdp_aon22 g4659 (.Z(w4780), .B2(w4753), .B1(w4770), .A1(w4769), .A2(w4777) );
	vdp_aon22 g4660 (.Z(w4778), .B2(w4753), .B1(w4773), .A1(w4772), .A2(w4777) );
	vdp_not g4661 (.nZ(w4775), .A(w4738) );
	vdp_not g4662 (.nZ(w4554), .A(w6559) );
	vdp_not g4663 (.nZ(w4555), .A(w4784) );
	vdp_not g4664 (.nZ(w4564), .A(w4788) );
	vdp_not g4665 (.nZ(w4558), .A(w4801) );
	vdp_not g4666 (.nZ(w4797), .A(w4793) );
	vdp_not g4667 (.nZ(w4557), .A(w4795) );
	vdp_dlatch_inv g4668 (.nQ(w4796), .D(w4793), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4669 (.nQ(w4795), .D(w4794), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g4670 (.nZ(w4556), .A(w4804) );
	vdp_dlatch_inv g4671 (.nQ(w4825), .D(w4759), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4672 (.nQ(w4804), .D(w4800), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g4673 (.nZ(w4805), .A(w4826) );
	vdp_dlatch_inv g4674 (.nQ(w4802), .D(w4826), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4675 (.nQ(w4815), .D(w4803), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g4676 (.nZ(w4799), .A(w4810) );
	vdp_dlatch_inv g4677 (.nQ(w4806), .D(w4810), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4678 (.nQ(w4816), .D(w4807), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4679 (.nQ(w4808), .D(w4798), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4680 (.nQ(w4813), .D(w4809), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4681 (.nQ(w4822), .D(w4811), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4682 (.nQ(w4824), .D(w4823), .nC(nHCLK2), .C(HCLK2) );
	vdp_sr_bit g4683 (.Q(w4550), .D(w6621), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4684 (.Z(w4811), .B2(w4753), .B1(1'b0), .A1(w4745), .A2(w4777) );
	vdp_aon22 g4685 (.Z(w4798), .B2(w4753), .B1(1'b0), .A1(w4755), .A2(w4777) );
	vdp_aon22 g4686 (.Z(w6621), .B2(w4851), .B1(M5), .A1(w127), .A2(w4897) );
	vdp_not g4687 (.nZ(w4841), .A(w1) );
	vdp_not g4688 (.nZ(w4900), .A(w4854) );
	vdp_not g4689 (.nZ(w4842), .A(w4853) );
	vdp_not g4690 (.nZ(w4898), .A(w4855) );
	vdp_not g4691 (.nZ(w4851), .A(w4852) );
	vdp_not g4692 (.nZ(w4897), .A(M5) );
	vdp_not g4693 (.nZ(w4846), .A(w4849) );
	vdp_not g4694 (.nZ(w4843), .A(w4550) );
	vdp_not g4695 (.nZ(w6630), .A(w4551) );
	vdp_not g4696 (.nZ(w4899), .A(M5) );
	vdp_not g4697 (.nZ(w4814), .A(w1) );
	vdp_not g4698 (.nZ(w4818), .A(w4750) );
	vdp_bufif0 g4699 (.A(1'b0), .Z(VRAMA[0]), .nE(w4647) );
	vdp_bufif0 g4700 (.A(w4635), .Z(VRAMA[1]), .nE(w4647) );
	vdp_bufif0 g4701 (.A(w4639), .Z(VRAMA[2]), .nE(w4647) );
	vdp_bufif0 g4702 (.A(w4642), .Z(VRAMA[3]), .nE(w4647) );
	vdp_bufif0 g4703 (.A(w4638), .Z(VRAMA[4]), .nE(w4647) );
	vdp_bufif0 g4704 (.A(w4636), .Z(VRAMA[5]), .nE(w4647) );
	vdp_bufif0 g4705 (.A(1'b0), .Z(VRAMA[6]), .nE(w4647) );
	vdp_bufif0 g4706 (.A(1'b0), .Z(VRAMA[7]), .nE(w4647) );
	vdp_aon22 g4707 (.Z(w4810), .B2(w4753), .B1(w6617), .A1(w4756), .A2(w4777) );
	vdp_aon22 g4708 (.Z(w4826), .B2(w4753), .B1(w4758), .A1(w4757), .A2(w4777) );
	vdp_aon22 g4709 (.Z(w4759), .B2(w4753), .B1(w4761), .A1(w4760), .A2(w4777) );
	vdp_comp_str g4710 (.A(w4774), .nZ(w4712), .Z(w4711) );
	vdp_and g4711 (.Z(w4737), .B(w4697), .A(w4693) );
	vdp_comp_we g4712 (.A(w4737), .nZ(w4777), .Z(w4753) );
	vdp_comp_str g4713 (.A(w4771), .nZ(w4727), .Z(w4726) );
	vdp_not g4714 (.nZ(w4693), .A(M5) );
	vdp_comp_str g4715 (.A(w4845), .nZ(w4856), .Z(w4848) );
	vdp_comp_str g4716 (.A(w4882), .nZ(w4864), .Z(w4869) );
	vdp_comp_we g4717 (.A(M5), .nZ(w4654), .Z(w4657) );
	vdp_comp_we g4718 (.A(w4689), .nZ(w4681), .Z(w4630) );
	vdp_comp_we g4719 (.A(w4668), .nZ(w4637), .Z(w4672) );
	vdp_comp_we g4720 (.A(M5), .nZ(w4644), .Z(w4640) );
	vdp_comp_we g4721 (.A(w1), .nZ(w4748), .Z(w4747) );
	vdp_comp_we g4722 (.nZ(w4863), .A(w4883), .Z(w4868) );
	vdp_and g4723 (.Z(w4774), .B(w4836), .A(DCLK2) );
	vdp_and g4724 (.Z(w4771), .B(w4838), .A(DCLK2) );
	vdp_and g4725 (.Z(w4835), .B(M5), .A(w4841) );
	vdp_and g4726 (.Z(w6633), .B(w4898), .A(M5) );
	vdp_and g4727 (.Z(w6632), .B(w4843), .A(w4551) );
	vdp_and g4728 (.Z(w4882), .B(w4881), .A(HCLK1) );
	vdp_or g4729 (.Z(w4817), .B(w4814), .A(w4824) );
	vdp_or g4730 (.Z(w6634), .B(w4899), .A(w4813) );
	vdp_and g4731 (.Z(w4632), .B(w4661), .A(w4645) );
	vdp_and g4732 (.Z(w4690), .B(w4626), .A(w4688) );
	vdp_and g4733 (.Z(w6374), .B(w4688), .A(w4627) );
	vdp_and g4734 (.Z(w6375), .B(w4625), .A(w4627) );
	vdp_and g4735 (.Z(w6376), .B(w4626), .A(w4625) );
	vdp_and g4736 (.Z(w6349), .B(H40), .A(VRAMA[9]) );
	vdp_or g4737 (.Z(w4699), .B(w4628), .A(w4697) );
	vdp_or g4738 (.Z(w4698), .B(w4628), .A(w4694) );
	vdp_not g4739 (.nZ(w4625), .A(w4688) );
	vdp_oai21 g4740 (.Z(w4652), .B(w30), .A1(w31), .A2(w5) );
	vdp_oai21 g4741 (.Z(w4849), .B(w4545), .A1(w4765), .A2(w4850) );
	vdp_aoi22 g4742 (.Z(w4738), .B2(w4693), .B1(w4694), .A1(M5), .A2(w4735) );
	vdp_or3 g4743 (.Z(w4735), .B(w4694), .A(w4695), .C(w4696) );
	vdp_and3 g4744 (.Z(w4845), .B(DCLK1), .A(HCLK2), .C(w4837) );
	vdp_oai21 g4745 (.Z(w4667), .B(M5), .A1(w4645), .A2(w4666) );
	vdp_2a3oi g4746 (.Z(w4659), .B(w4650), .A1(w4649), .A2(w4), .C(SYSRES) );
	vdp_or8 g4747 (.Z(w4850), .B(w4862), .A(M5), .C(w6564), .D(w4861), .F(w4859), .E(w4860), .G(w4858), .H(w4857) );
	vdp_and9 g4748 (.Z(w4512), .B(w4819), .A(w4821), .C(w4820), .D(w4818), .F(w4816), .E(w4817), .G(w4815), .H(w4812), .I(w6634) );
	vdp_nor12 g4749 (.Z(w4765), .B(w4759), .A(1'b0), .C(w4799), .D(M5), .F(w4811), .E(w4798), .G(w4805), .H(w4797), .J(w4780), .I(w4785), .K(w4778), .L(w4791) );
	vdp_or4 g4750 (.Z(w4689), .B(w4627), .A(w4626), .C(w4687), .D(w4629) );
	vdp_nand g4751 (.Z(w4776), .B(w4775), .A(HCLK1) );
	vdp_nand g4752 (.Z(w4821), .B(w4752), .A(w6631) );
	vdp_nand g4753 (.Z(w4820), .B(w4751), .A(w6630) );
	vdp_nor g4754 (.Z(w6631), .B(w4550), .A(w4551) );
	vdp_nand3 g4755 (.Z(w4819), .B(w4751), .A(w6632), .C(w4752) );
	vdp_sr_bit g4756 (.Q(w4553), .D(w4900), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4757 (.Q(w4908), .D(w28), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4758 (.Q(w4573), .D(w6553), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4759 (.Q(w4907), .D(w6537), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4760 (.Q(w6537), .D(w6538), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4761 (.Q(w6538), .D(w4906), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4762 (.Z(w4911), .B2(w4907), .B1(w5269), .A1(DB[4]), .A2(w5270) );
	vdp_notif0 g4763 (.A(HPOS[1]), .nZ(VRAMA[1]), .nE(w5128) );
	vdp_aon22 g4764 (.Z(w6553), .B2(w4905), .B1(w4908), .A1(M5), .A2(w28) );
	vdp_not g4765 (.nZ(w4905), .A(M5) );
	vdp_lfsr_bit g4766 (.Q(w4912), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6805), .A1(w4911), .A2(w6806) );
	vdp_lfsr_bit g4767 (.Q(w4915), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6803), .A1(w4912), .A2(w6804) );
	vdp_lfsr_bit g4768 (.Q(w4917), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6801), .A1(w4915), .A2(w6802) );
	vdp_lfsr_bit g4769 (.Q(w4918), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6799), .A1(w4917), .A2(w6800) );
	vdp_lfsr_bit g4770 (.Q(w4922), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6797), .A1(w4918), .A2(w6798) );
	vdp_lfsr_bit g4771 (.Q(w4920), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6795), .A1(w4922), .A2(w6796) );
	vdp_lfsr_bit g4772 (.Q(w4924), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6793), .A1(w4920), .A2(w6794) );
	vdp_lfsr_bit g4773 (.Q(w4904), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6792), .A1(w4924), .A2(w6791) );
	vdp_lfsr_bit g4774 (.Q(w4928), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5108), .A1(w4904), .A2(w6790) );
	vdp_lfsr_bit g4775 (.Q(w4930), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5273), .A1(w4928), .A2(w5274) );
	vdp_lfsr_bit g4776 (.Q(w4934), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5155), .A1(w4930), .A2(w5156) );
	vdp_lfsr_bit g4777 (.Q(w4931), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5152), .A1(w4934), .A2(w5153) );
	vdp_lfsr_bit g4778 (.Q(w4933), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5150), .A1(w4931), .A2(w5151) );
	vdp_lfsr_bit g4779 (.Q(w4937), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6788), .A1(w4933), .A2(w6787) );
	vdp_lfsr_bit g4780 (.Q(w4938), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5147), .A1(w4937), .A2(w5148) );
	vdp_lfsr_bit g4781 (.Q(w4942), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6785), .A1(w4938), .A2(w6786) );
	vdp_lfsr_bit g4782 (.Q(w4941), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6789), .A1(w4942), .A2(w6556) );
	vdp_lfsr_bit g4783 (.Q(w4946), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5144), .A1(w4941), .A2(w5145) );
	vdp_lfsr_bit g4784 (.Q(w4948), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5143), .A1(w4946), .A2(w5142) );
	vdp_lfsr_bit g4785 (.Q(w4903), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5140), .A1(w4948), .A2(w5141) );
	vdp_bufif0 g4786 (.A(w4904), .Z(VRAMA[1]), .nE(w6555) );
	vdp_bufif0 g4787 (.A(1'b0), .Z(VRAMA[1]), .nE(w5163) );
	vdp_notif0 g4788 (.A(w4903), .nZ(DB[4]), .nE(w5275) );
	vdp_sr_bit g4789 (.Q(w4955), .D(w6540), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4790 (.Q(w6540), .D(w6539), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4791 (.Q(w6539), .D(w6357), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4792 (.Z(w4910), .B2(w4955), .B1(w5269), .A1(DB[5]), .A2(w5270) );
	vdp_notif0 g4793 (.A(w4963), .nZ(VRAMA[2]), .nE(w5128) );
	vdp_lfsr_bit g4794 (.Q(w4913), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6805), .A1(w4910), .A2(w6806) );
	vdp_lfsr_bit g4795 (.Q(w4914), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6803), .A1(w4913), .A2(w6804) );
	vdp_lfsr_bit g4796 (.Q(w4916), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6801), .A1(w4914), .A2(w6802) );
	vdp_lfsr_bit g4797 (.Q(w4919), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6799), .A1(w4916), .A2(w6800) );
	vdp_lfsr_bit g4798 (.Q(w4923), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6797), .A1(w4919), .A2(w6798) );
	vdp_lfsr_bit g4799 (.Q(w4921), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6795), .A1(w4923), .A2(w6796) );
	vdp_lfsr_bit g4800 (.Q(w4925), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6793), .A1(w4921), .A2(w6794) );
	vdp_lfsr_bit g4801 (.Q(w4926), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6792), .A1(w4925), .A2(w6791) );
	vdp_lfsr_bit g4802 (.Q(w4929), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5108), .A1(w4926), .A2(w6790) );
	vdp_lfsr_bit g4803 (.Q(w4927), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5273), .A1(w4929), .A2(w5274) );
	vdp_lfsr_bit g4804 (.Q(w4935), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5155), .A1(w4927), .A2(w5156) );
	vdp_lfsr_bit g4805 (.Q(w4932), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5152), .A1(w4935), .A2(w5153) );
	vdp_lfsr_bit g4806 (.Q(w4936), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5150), .A1(w4932), .A2(w5151) );
	vdp_lfsr_bit g4807 (.Q(w4940), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6788), .A1(w4936), .A2(w6787) );
	vdp_lfsr_bit g4808 (.Q(w4939), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5147), .A1(w4940), .A2(w5148) );
	vdp_lfsr_bit g4809 (.Q(w4943), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6785), .A1(w4939), .A2(w6786) );
	vdp_lfsr_bit g4810 (.Q(w4944), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6789), .A1(w4943), .A2(w6556) );
	vdp_lfsr_bit g4811 (.Q(w4945), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5144), .A1(w4944), .A2(w5145) );
	vdp_lfsr_bit g4812 (.Q(w4949), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5143), .A1(w4945), .A2(w5142) );
	vdp_lfsr_bit g4813 (.Q(w4953), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5140), .A1(w4949), .A2(w5141) );
	vdp_bufif0 g4814 (.A(w4926), .Z(VRAMA[2]), .nE(w6555) );
	vdp_bufif0 g4815 (.A(1'b1), .Z(VRAMA[2]), .nE(w5163) );
	vdp_notif0 g4816 (.A(w4953), .nZ(DB[5]), .nE(w5275) );
	vdp_aon22 g4817 (.Z(w4952), .B2(w4942), .B1(w5137), .A1(w5136), .A2(w4903) );
	vdp_dlatch_inv g4818 (.nQ(w4964), .D(w4957), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g4819 (.nQ(w4959), .D(w4909), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g4820 (.Z(w4958), .B(w4959), .A(DCLK2) );
	vdp_nand g4821 (.Z(w4957), .B(HCLK1), .A(w4573) );
	vdp_nand g4822 (.Z(w4909), .B(HCLK1), .A(w28) );
	vdp_sr_bit g4823 (.Q(w4956), .D(w6542), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4824 (.Q(w6542), .D(w6541), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4825 (.Q(w6541), .D(w4961), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4826 (.Z(w4972), .B2(w4956), .B1(w5269), .A1(DB[6]), .A2(w5270) );
	vdp_notif0 g4827 (.A(w4970), .nZ(VRAMA[3]), .nE(w5128) );
	vdp_lfsr_bit g4828 (.Q(w4974), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6805), .A1(w4972), .A2(w6806) );
	vdp_lfsr_bit g4829 (.Q(w4975), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6803), .A1(w4974), .A2(w6804) );
	vdp_lfsr_bit g4830 (.Q(w4978), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6801), .A1(w4975), .A2(w6802) );
	vdp_lfsr_bit g4831 (.Q(w4979), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6799), .A1(w4978), .A2(w6800) );
	vdp_lfsr_bit g4832 (.Q(w4984), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6797), .A1(w4979), .A2(w6798) );
	vdp_lfsr_bit g4833 (.Q(w4983), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6795), .A1(w4984), .A2(w6796) );
	vdp_lfsr_bit g4834 (.Q(w4986), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6793), .A1(w4983), .A2(w6794) );
	vdp_lfsr_bit g4835 (.Q(w4988), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6792), .A1(w4986), .A2(w6791) );
	vdp_lfsr_bit g4836 (.Q(w4990), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5108), .A1(w4988), .A2(w6790) );
	vdp_lfsr_bit g4837 (.Q(w4992), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5273), .A1(w4990), .A2(w5274) );
	vdp_lfsr_bit g4838 (.Q(w4994), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5155), .A1(w4992), .A2(w5156) );
	vdp_lfsr_bit g4839 (.Q(w4996), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5152), .A1(w4994), .A2(w5153) );
	vdp_lfsr_bit g4840 (.Q(w4998), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5150), .A1(w4996), .A2(w5151) );
	vdp_lfsr_bit g4841 (.Q(w5001), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6788), .A1(w4998), .A2(w6787) );
	vdp_lfsr_bit g4842 (.Q(w5002), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5147), .A1(w5001), .A2(w5148) );
	vdp_lfsr_bit g4843 (.Q(w5003), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6785), .A1(w5002), .A2(w6786) );
	vdp_lfsr_bit g4844 (.Q(w5008), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6789), .A1(w5003), .A2(w6556) );
	vdp_lfsr_bit g4845 (.Q(w5007), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5144), .A1(w5008), .A2(w5145) );
	vdp_lfsr_bit g4846 (.Q(w5010), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5143), .A1(w5007), .A2(w5142) );
	vdp_lfsr_bit g4847 (.Q(w4954), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5140), .A1(w5010), .A2(w5141) );
	vdp_bufif0 g4848 (.A(w4988), .Z(VRAMA[3]), .nE(w6555) );
	vdp_bufif0 g4849 (.A(w4952), .Z(VRAMA[3]), .nE(w5163) );
	vdp_notif0 g4850 (.A(w4954), .nZ(DB[6]), .nE(w5275) );
	vdp_aon22 g4851 (.Z(w5011), .B2(w4943), .B1(w5137), .A1(w5136), .A2(w4953) );
	vdp_sr_bit g4852 (.Q(w4966), .D(w4964), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g4853 (.Q(w4960), .D(w4959), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_and g4854 (.Z(w4962), .B(w4964), .A(DCLK2) );
	vdp_and g4855 (.Z(w4968), .B(DCLK2), .A(w4966) );
	vdp_and g4856 (.Z(w4965), .B(w4960), .A(DCLK2) );
	vdp_sr_bit g4857 (.Q(w5024), .D(w6543), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4858 (.Q(w6543), .D(w6544), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4859 (.Q(w6544), .D(w4967), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4860 (.Z(w4971), .B2(w5024), .B1(w5269), .A1(DB[7]), .A2(w5270) );
	vdp_notif0 g4861 (.A(w5022), .nZ(VRAMA[4]), .nE(w5128) );
	vdp_lfsr_bit g4862 (.Q(w4973), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6805), .A1(w4971), .A2(w6806) );
	vdp_lfsr_bit g4863 (.Q(w4976), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6803), .A1(w4973), .A2(w6804) );
	vdp_lfsr_bit g4864 (.Q(w4977), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6801), .A1(w4976), .A2(w6802) );
	vdp_lfsr_bit g4865 (.Q(w4980), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6799), .A1(w4977), .A2(w6800) );
	vdp_lfsr_bit g4866 (.Q(w4981), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6797), .A1(w4980), .A2(w6798) );
	vdp_lfsr_bit g4867 (.Q(w4982), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6795), .A1(w4981), .A2(w6796) );
	vdp_lfsr_bit g4868 (.Q(w4985), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6793), .A1(w4982), .A2(w6794) );
	vdp_lfsr_bit g4869 (.Q(w4987), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6792), .A1(w4985), .A2(w6791) );
	vdp_lfsr_bit g4870 (.Q(w4989), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5108), .A1(w4987), .A2(w6790) );
	vdp_lfsr_bit g4871 (.Q(w4991), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5273), .A1(w4989), .A2(w5274) );
	vdp_lfsr_bit g4872 (.Q(w4993), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5155), .A1(w4991), .A2(w5156) );
	vdp_lfsr_bit g4873 (.Q(w4995), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5152), .A1(w4993), .A2(w5153) );
	vdp_lfsr_bit g4874 (.Q(w4997), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5150), .A1(w4995), .A2(w5151) );
	vdp_lfsr_bit g4875 (.Q(w5000), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6788), .A1(w4997), .A2(w6787) );
	vdp_lfsr_bit g4876 (.Q(w4999), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5147), .A1(w5000), .A2(w5148) );
	vdp_lfsr_bit g4877 (.Q(w5004), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6785), .A1(w4999), .A2(w6786) );
	vdp_lfsr_bit g4878 (.Q(w5005), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6789), .A1(w5004), .A2(w6556) );
	vdp_lfsr_bit g4879 (.Q(w5006), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5144), .A1(w5005), .A2(w5145) );
	vdp_lfsr_bit g4880 (.Q(w5009), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5143), .A1(w5006), .A2(w5142) );
	vdp_lfsr_bit g4881 (.Q(w5026), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5140), .A1(w5009), .A2(w5141) );
	vdp_bufif0 g4882 (.A(w4987), .Z(VRAMA[4]), .nE(w6555) );
	vdp_bufif0 g4883 (.A(w5011), .Z(VRAMA[4]), .nE(w5163) );
	vdp_notif0 g4884 (.A(w5026), .nZ(DB[7]), .nE(w5275) );
	vdp_aon22 g4885 (.Z(w5027), .B2(w5003), .B1(w5137), .A1(w5136), .A2(w4954) );
	vdp_aon22 g4886 (.Z(w5021), .B2(w5014), .B1(w127), .A1(w4969), .A2(w5020) );
	vdp_not g4887 (.nZ(w4969), .A(w127) );
	vdp_comp_str g4888 (.nZ(w5015), .A(w4965), .Z(w5016) );
	vdp_comp_str g4889 (.nZ(w5019), .A(w4968), .Z(w5018) );
	vdp_sr_bit g4890 (.Q(w5023), .D(w6546), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4891 (.Q(w6546), .D(w6545), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4892 (.Q(w6545), .D(w5017), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4893 (.Z(w5068), .B2(w5023), .B1(w5269), .A1(DB[8]), .A2(w5270) );
	vdp_notif0 g4894 (.A(w5021), .nZ(VRAMA[5]), .nE(w5128) );
	vdp_lfsr_bit g4895 (.Q(w5066), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6805), .A1(w5068), .A2(w6806) );
	vdp_lfsr_bit g4896 (.Q(w5063), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6803), .A1(w5066), .A2(w6804) );
	vdp_lfsr_bit g4897 (.Q(w5062), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6801), .A1(w5063), .A2(w6802) );
	vdp_lfsr_bit g4898 (.Q(w5059), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6799), .A1(w5062), .A2(w6800) );
	vdp_lfsr_bit g4899 (.Q(w5058), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6797), .A1(w5059), .A2(w6798) );
	vdp_lfsr_bit g4900 (.Q(w5055), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6795), .A1(w5058), .A2(w6796) );
	vdp_lfsr_bit g4901 (.Q(w5054), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6793), .A1(w5055), .A2(w6794) );
	vdp_lfsr_bit g4902 (.Q(w5032), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6792), .A1(w5054), .A2(w6791) );
	vdp_lfsr_bit g4903 (.Q(w5051), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5108), .A1(w5032), .A2(w6790) );
	vdp_lfsr_bit g4904 (.Q(w5025), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5273), .A1(w5051), .A2(w5274) );
	vdp_lfsr_bit g4905 (.Q(w5048), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5155), .A1(w5025), .A2(w5156) );
	vdp_lfsr_bit g4906 (.Q(w5047), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5152), .A1(w5048), .A2(w5153) );
	vdp_lfsr_bit g4907 (.Q(w5044), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5150), .A1(w5047), .A2(w5151) );
	vdp_lfsr_bit g4908 (.Q(w5042), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6788), .A1(w5044), .A2(w6787) );
	vdp_lfsr_bit g4909 (.Q(w5041), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5147), .A1(w5042), .A2(w5148) );
	vdp_lfsr_bit g4910 (.Q(w5030), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6785), .A1(w5041), .A2(w6786) );
	vdp_lfsr_bit g4911 (.Q(w5037), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6789), .A1(w5030), .A2(w6556) );
	vdp_lfsr_bit g4912 (.Q(w5035), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5144), .A1(w5037), .A2(w5145) );
	vdp_lfsr_bit g4913 (.Q(w5033), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5143), .A1(w5035), .A2(w5142) );
	vdp_lfsr_bit g4914 (.Q(w5050), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5140), .A1(w5033), .A2(w5141) );
	vdp_bufif0 g4915 (.A(w5032), .Z(VRAMA[5]), .nE(w6555) );
	vdp_bufif0 g4916 (.A(w5027), .Z(VRAMA[5]), .nE(w5163) );
	vdp_notif0 g4917 (.A(w5050), .nZ(DB[8]), .nE(w5275) );
	vdp_aon22 g4918 (.Z(w5029), .B2(w5004), .B1(w5137), .A1(w5136), .A2(w5026) );
	vdp_slatch g4919 (.D(S[0]), .nC(w5019), .C(w5018), .Q(w5073) );
	vdp_slatch g4920 (.D(S[0]), .nC(w5015), .C(w5016), .Q(w5013) );
	vdp_aoi22 g4921 (.Z(w5020), .B2(w5072), .B1(w5073), .A1(w5071), .A2(w5013) );
	vdp_sr_bit g4922 (.Q(w5081), .D(w6548), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4923 (.Q(w6548), .D(w6547), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4924 (.Q(w6547), .D(w5069), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4925 (.Z(w5067), .B2(w5081), .B1(w5269), .A1(DB[9]), .A2(w5270) );
	vdp_notif0 g4926 (.A(w5070), .nZ(VRAMA[6]), .nE(w5128) );
	vdp_lfsr_bit g4927 (.Q(w5065), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6805), .A1(w5067), .A2(w6806) );
	vdp_lfsr_bit g4928 (.Q(w5064), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6803), .A1(w5065), .A2(w6804) );
	vdp_lfsr_bit g4929 (.Q(w5061), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6801), .A1(w5064), .A2(w6802) );
	vdp_lfsr_bit g4930 (.Q(w5060), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6799), .A1(w5061), .A2(w6800) );
	vdp_lfsr_bit g4931 (.Q(w5057), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6797), .A1(w5060), .A2(w6798) );
	vdp_lfsr_bit g4932 (.Q(w5056), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6795), .A1(w5057), .A2(w6796) );
	vdp_lfsr_bit g4933 (.Q(w5053), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6793), .A1(w5056), .A2(w6794) );
	vdp_lfsr_bit g4934 (.Q(w5031), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6792), .A1(w5053), .A2(w6791) );
	vdp_lfsr_bit g4935 (.Q(w5052), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5108), .A1(w5031), .A2(w6790) );
	vdp_lfsr_bit g4936 (.Q(w5079), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5273), .A1(w5052), .A2(w5274) );
	vdp_lfsr_bit g4937 (.Q(w5049), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5155), .A1(w5079), .A2(w5156) );
	vdp_lfsr_bit g4938 (.Q(w5046), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5152), .A1(w5049), .A2(w5153) );
	vdp_lfsr_bit g4939 (.Q(w5045), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5150), .A1(w5046), .A2(w5151) );
	vdp_lfsr_bit g4940 (.Q(w5043), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6788), .A1(w5045), .A2(w6787) );
	vdp_lfsr_bit g4941 (.Q(w5040), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5147), .A1(w5043), .A2(w5148) );
	vdp_lfsr_bit g4942 (.Q(w5039), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6785), .A1(w5040), .A2(w6786) );
	vdp_lfsr_bit g4943 (.Q(w5038), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6789), .A1(w5039), .A2(w6556) );
	vdp_lfsr_bit g4944 (.Q(w5036), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5144), .A1(w5038), .A2(w5145) );
	vdp_lfsr_bit g4945 (.Q(w5034), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5143), .A1(w5036), .A2(w5142) );
	vdp_lfsr_bit g4946 (.Q(w5076), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5140), .A1(w5034), .A2(w5141) );
	vdp_bufif0 g4947 (.A(w5031), .Z(VRAMA[6]), .nE(w6555) );
	vdp_bufif0 g4948 (.A(w5029), .Z(VRAMA[6]), .nE(w5163) );
	vdp_notif0 g4949 (.A(w5076), .nZ(DB[9]), .nE(w5275) );
	vdp_aon22 g4950 (.Z(w5078), .B2(w5030), .B1(w5137), .A1(w5136), .A2(w5050) );
	vdp_aoi22 g4951 (.Z(w5070), .B2(w5072), .B1(w5083), .A1(w5071), .A2(w5074) );
	vdp_slatch g4952 (.D(S[1]), .nC(w5019), .C(w5018), .Q(w5083) );
	vdp_slatch g4953 (.D(S[1]), .nC(w5015), .C(w5016), .Q(w5074) );
	vdp_sr_bit g4954 (.Q(w5080), .D(w6550), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4955 (.Q(w6550), .D(w6549), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4956 (.Q(w6549), .D(w5084), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4957 (.Z(w5127), .B2(w5080), .B1(w5269), .A1(DB[10]), .A2(w5270) );
	vdp_notif0 g4958 (.A(w5130), .nZ(VRAMA[7]), .nE(w5131) );
	vdp_lfsr_bit g4959 (.Q(w5126), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6805), .A1(w5127), .A2(w6806) );
	vdp_lfsr_bit g4960 (.Q(w5121), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6803), .A1(w5126), .A2(w6804) );
	vdp_lfsr_bit g4961 (.Q(w5122), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6801), .A1(w5121), .A2(w6802) );
	vdp_lfsr_bit g4962 (.Q(w5116), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6799), .A1(w5122), .A2(w6800) );
	vdp_lfsr_bit g4963 (.Q(w5117), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6797), .A1(w5116), .A2(w6798) );
	vdp_lfsr_bit g4964 (.Q(w5114), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6795), .A1(w5117), .A2(w6796) );
	vdp_lfsr_bit g4965 (.Q(w5112), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6793), .A1(w5114), .A2(w6794) );
	vdp_lfsr_bit g4966 (.Q(w5077), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6792), .A1(w5112), .A2(w6791) );
	vdp_lfsr_bit g4967 (.Q(w5109), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5108), .A1(w5077), .A2(w6790) );
	vdp_lfsr_bit g4968 (.Q(w5104), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5273), .A1(w5109), .A2(w5274) );
	vdp_lfsr_bit g4969 (.Q(w5106), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5155), .A1(w5104), .A2(w5156) );
	vdp_lfsr_bit g4970 (.Q(w5103), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5152), .A1(w5106), .A2(w5153) );
	vdp_lfsr_bit g4971 (.Q(w5102), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5150), .A1(w5103), .A2(w5151) );
	vdp_lfsr_bit g4972 (.Q(w5099), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6788), .A1(w5102), .A2(w6787) );
	vdp_lfsr_bit g4973 (.Q(w5097), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5147), .A1(w5099), .A2(w5148) );
	vdp_lfsr_bit g4974 (.Q(w5095), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6785), .A1(w5097), .A2(w6786) );
	vdp_lfsr_bit g4975 (.Q(w5093), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6789), .A1(w5095), .A2(w6556) );
	vdp_lfsr_bit g4976 (.Q(w5091), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5144), .A1(w5093), .A2(w5145) );
	vdp_lfsr_bit g4977 (.Q(w5089), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5143), .A1(w5091), .A2(w5142) );
	vdp_lfsr_bit g4978 (.Q(w5087), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5140), .A1(w5089), .A2(w5141) );
	vdp_bufif0 g4979 (.A(w5077), .Z(VRAMA[7]), .nE(w6555) );
	vdp_bufif0 g4980 (.A(w5078), .Z(VRAMA[7]), .nE(w5163) );
	vdp_notif0 g4981 (.A(w5087), .nZ(DB[10]), .nE(w5275) );
	vdp_aon22 g4982 (.Z(w5086), .B2(w5039), .B1(w5137), .A1(w5136), .A2(w5076) );
	vdp_aoi22 g4983 (.Z(w5130), .B2(w5072), .B1(w5132), .A1(w5071), .A2(w5082) );
	vdp_slatch g4984 (.D(S[2]), .nC(w5019), .C(w5018), .Q(w5132) );
	vdp_slatch g4985 (.D(S[2]), .nC(w5015), .C(w5016), .Q(w5082) );
	vdp_sr_bit g4986 (.Q(w5158), .D(w29), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4987 (.Q(w5157), .D(w22), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4988 (.Z(w5124), .B2(w4548), .B1(w5269), .A1(DB[11]), .A2(w5270) );
	vdp_notif0 g4989 (.A(w5129), .nZ(VRAMA[8]), .nE(w5131) );
	vdp_lfsr_bit g4990 (.Q(w5125), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6805), .A1(w5124), .A2(w6806) );
	vdp_lfsr_bit g4991 (.Q(w5120), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6803), .A1(w5125), .A2(w6804) );
	vdp_lfsr_bit g4992 (.Q(w5123), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6801), .A1(w5120), .A2(w6802) );
	vdp_lfsr_bit g4993 (.Q(w5119), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6799), .A1(w5123), .A2(w6800) );
	vdp_lfsr_bit g4994 (.Q(w5118), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6797), .A1(w5119), .A2(w6798) );
	vdp_lfsr_bit g4995 (.Q(w5115), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6795), .A1(w5118), .A2(w6796) );
	vdp_lfsr_bit g4996 (.Q(w5113), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6793), .A1(w5115), .A2(w6794) );
	vdp_lfsr_bit g4997 (.Q(w5111), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6792), .A1(w5113), .A2(w6791) );
	vdp_lfsr_bit g4998 (.Q(w5110), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5108), .A1(w5111), .A2(w6790) );
	vdp_lfsr_bit g4999 (.Q(w5107), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5273), .A1(w5110), .A2(w5274) );
	vdp_lfsr_bit g5000 (.Q(w5105), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5155), .A1(w5107), .A2(w5156) );
	vdp_lfsr_bit g5001 (.Q(w5101), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5152), .A1(w5105), .A2(w5153) );
	vdp_lfsr_bit g5002 (.Q(w5100), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5150), .A1(w5101), .A2(w5151) );
	vdp_lfsr_bit g5003 (.Q(w5098), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6788), .A1(w5100), .A2(w6787) );
	vdp_lfsr_bit g5004 (.Q(w5096), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5147), .A1(w5098), .A2(w5148) );
	vdp_lfsr_bit g5005 (.Q(w5094), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6785), .A1(w5096), .A2(w6786) );
	vdp_lfsr_bit g5006 (.Q(w5092), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6789), .A1(w5094), .A2(w6556) );
	vdp_lfsr_bit g5007 (.Q(w5090), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5144), .A1(w5092), .A2(w5145) );
	vdp_lfsr_bit g5008 (.Q(w5088), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5143), .A1(w5090), .A2(w5142) );
	vdp_lfsr_bit g5009 (.Q(w5154), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5140), .A1(w5088), .A2(w5141) );
	vdp_bufif0 g5010 (.A(1'b0), .Z(VRAMA[0]), .nE(w6555) );
	vdp_bufif0 g5011 (.A(w5086), .Z(VRAMA[8]), .nE(w5163) );
	vdp_notif0 g5012 (.A(w5154), .nZ(DB[11]), .nE(w5275) );
	vdp_aon22 g5013 (.Z(w5164), .B2(w5138), .B1(w5137), .A1(w5136), .A2(w5087) );
	vdp_aoi22 g5014 (.Z(w5129), .B2(w5072), .B1(w5133), .A1(w5071), .A2(w5134) );
	vdp_slatch g5015 (.D(S[3]), .nC(w5019), .C(w5018), .Q(w5133) );
	vdp_slatch g5016 (.D(S[3]), .nC(w5015), .C(w5016), .Q(w5134) );
	vdp_bufif0 g5017 (.A(1'b0), .Z(VRAMA[0]), .nE(w5163) );
	vdp_bufif0 g5018 (.A(w5167), .Z(VRAMA[8]), .nE(w5171) );
	vdp_aon22 g5019 (.Z(w5194), .B2(w4558), .B1(w5269), .A1(DB[3]), .A2(w5270) );
	vdp_lfsr_bit g5020 (.Q(w5192), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6805), .A1(w5194), .A2(w6806) );
	vdp_lfsr_bit g5021 (.Q(w5190), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6803), .A1(w5192), .A2(w6804) );
	vdp_lfsr_bit g5022 (.Q(w5188), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6801), .A1(w5190), .A2(w6802) );
	vdp_lfsr_bit g5023 (.Q(w5186), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6799), .A1(w5188), .A2(w6800) );
	vdp_lfsr_bit g5024 (.Q(w5183), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6797), .A1(w5186), .A2(w6798) );
	vdp_lfsr_bit g5025 (.Q(w5182), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6795), .A1(w5183), .A2(w6796) );
	vdp_lfsr_bit g5026 (.Q(w5180), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6793), .A1(w5182), .A2(w6794) );
	vdp_lfsr_bit g5027 (.Q(w5178), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6792), .A1(w5180), .A2(w6791) );
	vdp_lfsr_bit g5028 (.Q(w5162), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5108), .A1(w5178), .A2(w6790) );
	vdp_lfsr_bit g5029 (.Q(w5160), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5273), .A1(w5162), .A2(w5274) );
	vdp_notif0 g5030 (.A(w5160), .nZ(DB[3]), .nE(w5275) );
	vdp_not g5031 (.nZ(w5149), .A(M5) );
	vdp_not g5032 (.nZ(w5159), .A(H40) );
	vdp_notif0 g5033 (.A(1'b1), .nZ(VRAMA[0]), .nE(w5128) );
	vdp_aoi22 g5034 (.Z(w5014), .B2(w5198), .B1(w5162), .A1(w5071), .A2(w5160) );
	vdp_not g5035 (.nZ(w5196), .A(M5) );
	vdp_or g5036 (.Z(w5197), .B(w5158), .A(w5157) );
	vdp_sr_bit g5037 (.Q(w5168), .D(w9), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5038 (.Q(w5174), .D(w30), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_comp_we g5039 (.nZ(w5140), .A(w5166), .Z(w5141) );
	vdp_comp_we g5040 (.nZ(w5143), .A(w5166), .Z(w5142) );
	vdp_comp_we g5041 (.nZ(w5144), .A(w5166), .Z(w5145) );
	vdp_comp_we g5042 (.nZ(w6789), .A(w5166), .Z(w6556) );
	vdp_comp_we g5043 (.nZ(w6785), .A(w5166), .Z(w6786) );
	vdp_comp_we g5044 (.nZ(w5137), .A(H40), .Z(w5136) );
	vdp_comp_we g5045 (.nZ(w5147), .A(w5166), .Z(w5148) );
	vdp_comp_we g5046 (.nZ(w6788), .A(w5166), .Z(w6787) );
	vdp_comp_we g5047 (.nZ(w5150), .A(w5166), .Z(w5151) );
	vdp_comp_we g5048 (.nZ(w5152), .A(w5166), .Z(w5153) );
	vdp_comp_we g5049 (.nZ(w5155), .A(w5166), .Z(w5156) );
	vdp_comp_we g5050 (.nZ(w5072), .A(w5157), .Z(w5071) );
	vdp_not g5051 (.nZ(w5131), .A(w5161) );
	vdp_not g5052 (.nZ(w5128), .A(w5161) );
	vdp_not g5053 (.nZ(w5163), .A(w5170) );
	vdp_not g5054 (.nZ(w6555), .A(w5146) );
	vdp_and g5055 (.Z(w5146), .B(w5168), .A(w5149) );
	vdp_oai21 g5056 (.Z(w5173), .B(w5149), .A1(w5174), .A2(w5168) );
	vdp_aon333 g5057 (.Z(w4511), .B1(M5), .A1(1'b1), .C1(M5), .A2(w5149), .A3(w5111), .B2(w5094), .B3(w5159), .C2(H40), .C3(w5154) );
	vdp_aon22 g5058 (.Z(w5193), .B2(w4564), .B1(w5269), .A1(DB[2]), .A2(w5270) );
	vdp_lfsr_bit g5059 (.Q(w5191), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6805), .A1(w5193), .A2(w6806) );
	vdp_lfsr_bit g5060 (.Q(w5189), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6803), .A1(w5191), .A2(w6804) );
	vdp_lfsr_bit g5061 (.Q(w5187), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6801), .A1(w5189), .A2(w6802) );
	vdp_lfsr_bit g5062 (.Q(w5185), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6799), .A1(w5187), .A2(w6800) );
	vdp_lfsr_bit g5063 (.Q(w5184), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6797), .A1(w5185), .A2(w6798) );
	vdp_lfsr_bit g5064 (.Q(w5181), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6795), .A1(w5184), .A2(w6796) );
	vdp_lfsr_bit g5065 (.Q(w5179), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6793), .A1(w5181), .A2(w6794) );
	vdp_lfsr_bit g5066 (.Q(w5177), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6792), .A1(w5179), .A2(w6791) );
	vdp_lfsr_bit g5067 (.Q(w5176), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5108), .A1(w5177), .A2(w6790) );
	vdp_lfsr_bit g5068 (.Q(w5175), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5273), .A1(w5176), .A2(w5274) );
	vdp_notif0 g5069 (.A(w5175), .nZ(DB[2]), .nE(w5275) );
	vdp_aoi22 g5070 (.Z(w5022), .B2(w5198), .B1(w5176), .A1(w5071), .A2(w5175) );
	vdp_aoi22 g5071 (.Z(w5211), .B2(w5198), .B1(w5212), .A1(w5071), .A2(w4513) );
	vdp_notif0 g5072 (.A(w5211), .nZ(VRAMA[9]), .nE(w5131) );
	vdp_slatch g5074 (.D(S[4]), .nC(w5016), .C(w5015), .Q(w4513) );
	vdp_and g5075 (.Z(w5161), .B(w5196), .A(w5197) );
	vdp_slatch g5076 (.D(REG_BUS[0]), .nC(w5272), .C(w5271), .Q(w5138) );
	vdp_slatch g5077 (.D(REG_BUS[7]), .nC(w5272), .C(w5271), .Q(w5169) );
	vdp_bufif0 g5078 (.A(w5164), .Z(VRAMA[9]), .nE(w5201) );
	vdp_bufif0 g5079 (.A(w5169), .Z(VRAMA[16]), .nE(w5201) );
	vdp_and g5080 (.Z(w5170), .B(w5168), .A(M5) );
	vdp_not g5081 (.nZ(w5201), .A(w5170) );
	vdp_not g5082 (.nZ(w5171), .A(w5172) );
	vdp_not g5083 (.nZ(w5172), .A(w5173) );
	vdp_xor g5084 (.Z(w5200), .B(w5169), .A(VRAMA[16]) );
	vdp_xor g5085 (.Z(w5204), .B(w5206), .A(w5205) );
	vdp_and3 g5086 (.Z(w6355), .B(w5210), .A(w5207), .C(M5) );
	vdp_nor g5087 (.Z(w5206), .B(H40), .A(w5138) );
	vdp_nor g5088 (.Z(w5205), .B(H40), .A(VRAMA[9]) );
	vdp_aon22 g5089 (.Z(w5231), .B2(w4555), .B1(w5269), .A1(DB[1]), .A2(w5270) );
	vdp_lfsr_bit g5090 (.Q(w5230), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6805), .A1(w5231), .A2(w6806) );
	vdp_lfsr_bit g5091 (.Q(w5229), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6803), .A1(w5230), .A2(w6804) );
	vdp_lfsr_bit g5092 (.Q(w5228), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6801), .A1(w5229), .A2(w6802) );
	vdp_lfsr_bit g5093 (.Q(w5227), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6799), .A1(w5228), .A2(w6800) );
	vdp_lfsr_bit g5094 (.Q(w5226), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6797), .A1(w5227), .A2(w6798) );
	vdp_lfsr_bit g5095 (.Q(w5225), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6795), .A1(w5226), .A2(w6796) );
	vdp_lfsr_bit g5096 (.Q(w5224), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6793), .A1(w5225), .A2(w6794) );
	vdp_lfsr_bit g5097 (.Q(w5223), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6792), .A1(w5224), .A2(w6791) );
	vdp_lfsr_bit g5098 (.Q(w5209), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5108), .A1(w5223), .A2(w6790) );
	vdp_lfsr_bit g5099 (.Q(w5221), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5273), .A1(w5209), .A2(w5274) );
	vdp_notif0 g5100 (.A(w5221), .nZ(DB[1]), .nE(w5275) );
	vdp_slatch g5101 (.D(REG_BUS[1]), .nC(w5272), .C(w5271), .Q(w5167) );
	vdp_slatch g5102 (.D(REG_BUS[6]), .nC(w5272), .C(w5271), .Q(w5220) );
	vdp_xor g5103 (.Z(w5203), .B(w5220), .A(VRAMA[15]) );
	vdp_xor g5104 (.Z(w5202), .B(w5167), .A(VRAMA[10]) );
	vdp_aon22 g5105 (.Z(w5240), .B2(w4554), .B1(w5269), .A1(DB[0]), .A2(w5270) );
	vdp_lfsr_bit g5106 (.Q(w5241), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6805), .A1(w5240), .A2(w6806) );
	vdp_lfsr_bit g5107 (.Q(w5242), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6803), .A1(w5241), .A2(w6804) );
	vdp_lfsr_bit g5108 (.Q(w5243), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6801), .A1(w5242), .A2(w6802) );
	vdp_lfsr_bit g5109 (.Q(w5245), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6799), .A1(w5243), .A2(w6800) );
	vdp_lfsr_bit g5110 (.Q(w5244), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6797), .A1(w5245), .A2(w6798) );
	vdp_lfsr_bit g5111 (.Q(w5247), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6795), .A1(w5244), .A2(w6796) );
	vdp_lfsr_bit g5112 (.Q(w5246), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6793), .A1(w5247), .A2(w6794) );
	vdp_lfsr_bit g5113 (.Q(w5248), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6792), .A1(w5246), .A2(w6791) );
	vdp_lfsr_bit g5114 (.Q(w5222), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5108), .A1(w5248), .A2(w6790) );
	vdp_lfsr_bit g5115 (.Q(w6554), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5273), .A1(w5222), .A2(w5274) );
	vdp_notif0 g5116 (.A(w6554), .nZ(DB[0]), .nE(w5275) );
	vdp_slatch g5117 (.D(REG_BUS[2]), .nC(w5272), .C(w5271), .Q(w5219) );
	vdp_slatch g5118 (.D(REG_BUS[5]), .nC(w5272), .C(w5271), .Q(w5263) );
	vdp_xor g5119 (.Z(w5216), .B(w5263), .A(VRAMA[14]) );
	vdp_xor g5120 (.Z(w5215), .B(w5219), .A(VRAMA[11]) );
	vdp_slatch g5121 (.D(S[5]), .nC(w5018), .C(w5019), .Q(w5234) );
	vdp_slatch g5122 (.D(S[5]), .nC(w5016), .C(w5015), .Q(w5213) );
	vdp_slatch g5123 (.D(S[6]), .nC(w5018), .C(w5019), .Q(w5235) );
	vdp_slatch g5124 (.D(S[6]), .nC(w5016), .C(w5015), .Q(w5233) );
	vdp_slatch g5125 (.D(S[7]), .nC(w5018), .C(w5019), .Q(w5268) );
	vdp_slatch g5126 (.D(S[7]), .nC(w5016), .C(w5015), .Q(w5198) );
	vdp_slatch g5127 (.D(REG_BUS[2]), .nC(w5238), .C(w5239), .Q(w5236) );
	vdp_slatch g5128 (.D(REG_BUS[5]), .nC(w5238), .C(w5239), .Q(w5232) );
	vdp_bufif0 g5129 (.A(w5219), .Z(VRAMA[9]), .nE(w5171) );
	vdp_bufif0 g5130 (.A(w5167), .Z(VRAMA[10]), .nE(w5201) );
	vdp_bufif0 g5131 (.A(w5257), .Z(VRAMA[10]), .nE(w5171) );
	vdp_bufif0 g5132 (.A(w5220), .Z(VRAMA[13]), .nE(w5171) );
	vdp_bufif0 g5133 (.A(w5263), .Z(VRAMA[14]), .nE(w5201) );
	vdp_bufif0 g5134 (.A(w5219), .Z(VRAMA[11]), .nE(w5201) );
	vdp_bufif0 g5135 (.A(w5256), .Z(VRAMA[13]), .nE(w5201) );
	vdp_bufif0 g5136 (.A(w5257), .Z(VRAMA[12]), .nE(w5201) );
	vdp_bufif0 g5137 (.A(w5256), .Z(VRAMA[11]), .nE(w5171) );
	vdp_bufif0 g5138 (.A(w5263), .Z(VRAMA[12]), .nE(w5171) );
	vdp_bufif0 g5139 (.A(w5220), .Z(VRAMA[15]), .nE(w5201) );
	vdp_slatch g5140 (.D(REG_BUS[3]), .nC(w5272), .C(w5271), .Q(w5257) );
	vdp_slatch g5141 (.D(REG_BUS[4]), .nC(w5272), .C(w5271), .Q(w5256) );
	vdp_xor g5142 (.Z(w5218), .B(w5256), .A(VRAMA[13]) );
	vdp_xor g5143 (.Z(w5217), .B(w5257), .A(VRAMA[12]) );
	vdp_dlatch_inv g5144 (.nQ(w5255), .D(w5260), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5145 (.nQ(w5254), .D(w5261), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5146 (.nQ(w5253), .D(w6661), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5147 (.nQ(w5252), .D(w6663), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5148 (.nQ(w5251), .D(w5262), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5149 (.nQ(w5250), .D(w5259), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5150 (.nQ(w5249), .D(w6662), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5151 (.nQ(w6350), .D(w5258), .nC(nDCLK1), .C(DCLK1) );
	vdp_comp_we g5152 (.nZ(w5273), .A(w5166), .Z(w5274) );
	vdp_comp_we g5153 (.nZ(w5108), .A(w5166), .Z(w6790) );
	vdp_comp_we g5154 (.nZ(w6792), .A(w5166), .Z(w6791) );
	vdp_comp_we g5155 (.nZ(w6793), .A(w5166), .Z(w6794) );
	vdp_comp_we g5156 (.nZ(w6795), .A(w5166), .Z(w6796) );
	vdp_comp_we g5157 (.nZ(w6797), .A(w5166), .Z(w6798) );
	vdp_comp_we g5158 (.nZ(w6799), .A(w5166), .Z(w6800) );
	vdp_comp_we g5159 (.nZ(w6801), .A(w5166), .Z(w6802) );
	vdp_comp_we g5160 (.nZ(w6803), .A(w5166), .Z(w6804) );
	vdp_comp_we g5161 (.nZ(w6805), .A(w5166), .Z(w6806) );
	vdp_comp_we g5162 (.nZ(w5269), .A(w114), .Z(w5270) );
	vdp_notif0 g5163 (.A(w5208), .nZ(VRAMA[10]), .nE(w5131) );
	vdp_notif0 g5164 (.A(w5237), .nZ(VRAMA[13]), .nE(w5131) );
	vdp_notif0 g5165 (.A(w5267), .nZ(VRAMA[11]), .nE(w5131) );
	vdp_notif0 g5166 (.A(w5266), .nZ(VRAMA[12]), .nE(w5131) );
	vdp_not g5167 (.nZ(w5210), .A(VRAMA[2]) );
	vdp_not g5168 (.nZ(w5237), .A(w5236) );
	vdp_not g5169 (.nZ(w5265), .A(w119) );
	vdp_aoi22 g5170 (.Z(w4970), .B2(w5198), .B1(w5209), .A1(w5071), .A2(w5221) );
	vdp_aoi22 g5171 (.Z(w5208), .B2(w5198), .B1(w5234), .A1(w5071), .A2(w5213) );
	vdp_aoi22 g5172 (.Z(w4963), .B2(w5198), .B1(w5222), .A1(w5071), .A2(w6554) );
	vdp_aoi22 g5173 (.Z(w5267), .B2(w5198), .B1(w5235), .A1(w5071), .A2(w5233) );
	vdp_aoi22 g5174 (.Z(w5266), .B2(w5198), .B1(w5268), .A1(w5071), .A2(w5198) );
	vdp_and g5175 (.Z(w5264), .B(w5265), .A(w4546) );
	vdp_nor8 g5176 (.Z(w5207), .B(w5217), .A(w5218), .C(w5216), .D(w5215), .F(w5204), .E(w5200), .G(w5202), .H(w5203) );
	vdp_not g5177 (.nZ(w5275), .A(w118) );
	vdp_comp_str g5178 (.nZ(w5272), .A(w137), .Z(w5271) );
	vdp_comp_str g5179 (.nZ(w5239), .A(w138), .Z(w5238) );
	vdp_or3 g5180 (.Z(w5166), .B(w114), .A(w118), .C(w5264) );
	vdp_not g5181 (.nZ(S[7]), .A(w5255) );
	vdp_not g5182 (.nZ(S[6]), .A(w5254) );
	vdp_not g5183 (.nZ(S[5]), .A(w5253) );
	vdp_not g5184 (.nZ(S[4]), .A(w5252) );
	vdp_not g5185 (.nZ(S[3]), .A(w5251) );
	vdp_not g5186 (.nZ(S[2]), .A(w5250) );
	vdp_not g5187 (.nZ(S[1]), .A(w5249) );
	vdp_not g5188 (.nZ(S[0]), .A(w6350) );
	vdp_aon21_sr g5189 (.Q(w5351), .A1(w5350), .A2(w6455), .B(w6462), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5190 (.Q(w6462), .A1(w5318), .A2(w6455), .B(w6461), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5191 (.Q(w6461), .A1(w5317), .A2(w6455), .B(w6460), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5192 (.Q(w6460), .A1(w5316), .A2(w6455), .B(w6459), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5193 (.Q(w6459), .A1(w5315), .A2(w6455), .B(w6458), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5194 (.Q(w6458), .A1(w5314), .A2(w6455), .B(w6457), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5195 (.Q(w6457), .A1(w5313), .A2(w6455), .B(w6456), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5196 (.Q(w6456), .A1(w5312), .A2(w6455), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5197 (.Q(w6464), .A1(w5307), .A2(w6463), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5198 (.Q(w6465), .A1(w5306), .A2(w6463), .B(w6464), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5199 (.Q(w6466), .A1(w5305), .A2(w6463), .B(w6465), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5200 (.Q(w6467), .A1(w5304), .A2(w6463), .B(w6466), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5201 (.Q(w6468), .A1(w5303), .A2(w6463), .B(w6467), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5202 (.Q(w6469), .A1(w5302), .A2(w6463), .B(w6468), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5203 (.Q(w6470), .A1(w5301), .A2(w6463), .B(w6469), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5204 (.Q(w5332), .A1(w5321), .A2(w6463), .B(w6470), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5205 (.Q(w5457), .A1(w5296), .A2(w6447), .B(w6448), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5206 (.Q(w6448), .A1(w5295), .A2(w6447), .B(w6449), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5207 (.Q(w6449), .A1(w5294), .A2(w6447), .B(w6450), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5208 (.Q(w6450), .A1(w5293), .A2(w6447), .B(w6451), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5209 (.Q(w6451), .A1(w5292), .A2(w6447), .B(w6452), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5210 (.Q(w6452), .A1(w5291), .A2(w6447), .B(w6453), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5211 (.Q(w6453), .A1(w5290), .A2(w6447), .B(w6454), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5212 (.Q(w6454), .A1(w5289), .A2(w6447), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5213 (.Q(w6440), .A1(w5284), .A2(w6439), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5214 (.Q(w6441), .A1(w5283), .A2(w6439), .B(w6440), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5215 (.Q(w6442), .A1(w5282), .A2(w6439), .B(w6441), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5216 (.Q(w6443), .A1(w5281), .A2(w6439), .B(w6442), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5217 (.Q(w6445), .A1(w5359), .A2(w6439), .B(w6443), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5218 (.Q(w6444), .A1(w5364), .A2(w6439), .B(w6445), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5219 (.Q(w6446), .A1(w5358), .A2(w6439), .B(w6444), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5220 (.Q(w5280), .A1(w5279), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .A2(w6439), .B(w6446) );
	vdp_not g5221 (.nZ(w6447), .A(w5344) );
	vdp_not g5222 (.nZ(w6439), .A(w5344) );
	vdp_not g5223 (.nZ(w6463), .A(w5344) );
	vdp_not g5224 (.nZ(w6455), .A(w5344) );
	vdp_or4 g5225 (.Z(w5349), .B(w5310), .A(w5367), .D(w5345), .C(w5311) );
	vdp_or4 g5226 (.Z(w5336), .B(w5308), .A(w5339), .D(w5343), .C(w5309) );
	vdp_or4 g5227 (.Z(w5352), .B(w5320), .A(w5279), .D(w5693), .C(w5319) );
	vdp_or4 g5228 (.Z(w5335), .B(w5300), .A(w5689), .D(w5358), .C(w5299) );
	vdp_or4 g5229 (.Z(w5331), .B(w5298), .A(w5688), .D(w5364), .C(w5297) );
	vdp_or4 g5230 (.Z(w5355), .B(w5286), .A(w5285), .D(w6351), .C(w5287) );
	vdp_or4 g5231 (.Z(w5326), .B(w5324), .A(w5325), .D(w5288), .C(w5323) );
	vdp_slatch g5232 (.Q(w5345), .D(w5403), .nC(w5340), .C(w5341) );
	vdp_comp_str g5233 (.nZ(w5340), .A(w5375), .Z(w5341) );
	vdp_slatch g5234 (.Q(w5311), .D(w5401), .nC(w5340), .C(w5341) );
	vdp_slatch g5235 (.Q(w5310), .D(w5400), .nC(w5340), .C(w5341) );
	vdp_slatch g5236 (.Q(w5367), .D(w5399), .nC(w5340), .C(w5341) );
	vdp_slatch g5237 (.Q(w5343), .D(w5398), .nC(w5340), .C(w5341) );
	vdp_slatch g5238 (.Q(w5309), .D(w5397), .nC(w5340), .C(w5341) );
	vdp_slatch g5239 (.Q(w5308), .D(w5395), .nC(w5340), .C(w5341) );
	vdp_slatch g5240 (.Q(w5339), .D(w5391), .nC(w5340), .C(w5341) );
	vdp_slatch g5241 (.Q(w5288), .D(w6436), .nC(w5322), .C(w5357) );
	vdp_slatch g5242 (.Q(w5323), .D(w6437), .nC(w5322), .C(w5357) );
	vdp_slatch g5243 (.Q(w5324), .D(w6438), .nC(w5322), .C(w5357) );
	vdp_slatch g5244 (.Q(w5325), .D(w5381), .nC(w5322), .C(w5357) );
	vdp_slatch g5245 (.Q(w6351), .D(w5379), .nC(w5322), .C(w5357) );
	vdp_slatch g5246 (.Q(w5287), .D(w5378), .nC(w5322), .C(w5357) );
	vdp_slatch g5247 (.Q(w5286), .D(w5377), .nC(w5322), .C(w5357) );
	vdp_slatch g5248 (.Q(w5285), .D(w5374), .nC(w5322), .C(w5357) );
	vdp_aon22 g5249 (.Z(w5411), .B2(w5328), .B1(w5362), .A1(w5355), .A2(w5334) );
	vdp_comp_we g5250 (.nZ(w5328), .A(w5361), .Z(w5334) );
	vdp_notif0 g5251 (.A(w5356), .nZ(DB[11]), .nE(w5373) );
	vdp_notif0 g5252 (.A(w5360), .nZ(DB[3]), .nE(w5373) );
	vdp_notif0 g5253 (.A(w5329), .nZ(DB[10]), .nE(w5373) );
	vdp_notif0 g5254 (.A(w5330), .nZ(DB[2]), .nE(w5373) );
	vdp_notif0 g5255 (.A(w5338), .nZ(DB[1]), .nE(w5373) );
	vdp_notif0 g5256 (.A(w5365), .nZ(DB[9]), .nE(w5373) );
	vdp_notif0 g5257 (.A(w5347), .nZ(DB[8]), .nE(w5373) );
	vdp_notif0 g5258 (.A(w5348), .nZ(DB[0]), .nE(w5373) );
	vdp_not g5259 (.nZ(w5353), .A(w5352) );
	vdp_aon22 g5260 (.Z(w5384), .B2(w5328), .B1(w5333), .A1(w5326), .A2(w5334) );
	vdp_aon22 g5261 (.Z(w5389), .B2(w5328), .B1(w5337), .A1(w5336), .A2(w5334) );
	vdp_aon22 g5262 (.Z(w5406), .B2(w5328), .B1(w5353), .A1(w5349), .A2(w5334) );
	vdp_comp_str g5263 (.nZ(w5322), .A(w5375), .Z(w5357) );
	vdp_not g5264 (.nZ(w5362), .A(w5363) );
	vdp_not g5265 (.nZ(w5333), .A(w5331) );
	vdp_not g5266 (.nZ(w5337), .A(w5335) );
	vdp_and3 g5267 (.Z(w5789), .B(w5387), .A(w5336), .C(w5335) );
	vdp_and3 g5268 (.Z(w5393), .B(w5407), .A(w5349), .C(w5352) );
	vdp_and3 g5269 (.Z(w5409), .B(w5385), .A(w5326), .C(w5331) );
	vdp_and3 g5270 (.Z(w5746), .B(w5355), .A(w5368), .C(w5363) );
	vdp_aon2222 g5271 (.Z(w5360), .B2(w5281), .B1(w5371), .A1(w5372), .A2(w5283), .D2(w5279), .D1(w5369), .C1(w5370), .C2(w5364) );
	vdp_aon2222 g5272 (.Z(w5356), .B2(w5282), .B1(w5371), .A1(w5372), .A2(w5284), .D2(w5358), .D1(w5369), .C1(w5370), .C2(w5359) );
	vdp_aon2222 g5273 (.Z(w5329), .B2(w5291), .B1(w5371), .A1(w5372), .A2(w5289), .D2(w5295), .D1(w5369), .C1(w5370), .C2(w5293) );
	vdp_aon2222 g5274 (.Z(w5330), .B2(w5292), .B1(w5371), .A1(w5372), .A2(w5290), .D2(w5296), .D1(w5369), .C1(w5370), .C2(w5294) );
	vdp_aon2222 g5275 (.Z(w5338), .B2(w5304), .B1(w5371), .A1(w5372), .A2(w5306), .D2(w5321), .D1(w5369), .C1(w5370), .C2(w5302) );
	vdp_aon2222 g5276 (.Z(w5365), .B2(w5305), .B1(w5371), .A1(w5372), .A2(w5307), .D2(w5301), .D1(w5369), .C1(w5370), .C2(w5303) );
	vdp_aon2222 g5277 (.Z(w5347), .B2(w5314), .B1(w5371), .A1(w5372), .A2(w5312), .D2(w5318), .D1(w5369), .C1(w5370), .C2(w5316) );
	vdp_aon2222 g5278 (.Z(w5348), .B2(w5315), .B1(w5371), .A1(w5372), .A2(w5313), .D2(w5350), .D1(w5369), .C1(w5370), .C2(w5317) );
	vdp_slatch g5279 (.Q(w5403), .D(w5424), .nC(w5423), .C(w5402) );
	vdp_comp_str g5280 (.nZ(w5423), .A(w5422), .Z(w5402) );
	vdp_slatch g5281 (.Q(w5401), .D(w5428), .nC(w5423), .C(w5402) );
	vdp_slatch g5282 (.Q(w5400), .D(w5429), .nC(w5423), .C(w5402) );
	vdp_slatch g5283 (.Q(w5399), .D(w5432), .nC(w5423), .C(w5402) );
	vdp_slatch g5284 (.Q(w5398), .D(w5437), .nC(w5438), .C(w5396) );
	vdp_comp_str g5285 (.nZ(w5438), .A(w5433), .Z(w5396) );
	vdp_slatch g5286 (.Q(w5397), .D(w5440), .nC(w5438), .C(w5396) );
	vdp_slatch g5287 (.Q(w5395), .D(w5441), .nC(w5438), .C(w5396) );
	vdp_slatch g5288 (.Q(w5391), .D(w5443), .nC(w5438), .C(w5396) );
	vdp_sr_bit g5289 (.Q(w5445), .D(w5332), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5290 (.nQ(w5390), .D(w5447), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5291 (.nQ(w5449), .D(w5388), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5292 (.nQ(w5386), .D(w5456), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5293 (.nQ(w5462), .D(w6394), .nC(nDCLK2), .C(DCLK2) );
	vdp_slatch g5294 (.Q(w5381), .D(w5424), .nC(w5464), .C(w5383) );
	vdp_slatch g5295 (.Q(w6436), .D(w5428), .nC(w5464), .C(w5383) );
	vdp_slatch g5296 (.Q(w6437), .D(w5429), .nC(w5464), .C(w5383) );
	vdp_slatch g5297 (.Q(w6438), .D(w5432), .nC(w5464), .C(w5383) );
	vdp_comp_str g5298 (.nZ(w5464), .A(w5463), .Z(w5383) );
	vdp_slatch g5299 (.Q(w5379), .D(w5437), .nC(w5475), .C(w5376) );
	vdp_slatch g5300 (.Q(w5378), .D(w5440), .nC(w5475), .C(w5376) );
	vdp_slatch g5301 (.Q(w5377), .D(w5441), .nC(w5475), .C(w5376) );
	vdp_slatch g5302 (.Q(w5374), .D(w5443), .nC(w5475), .C(w5376) );
	vdp_comp_str g5303 (.nZ(w5475), .A(w5480), .Z(w5376) );
	vdp_dlatch_inv g5304 (.nQ(w5473), .D(w5472), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5305 (.nQ(w5476), .D(w6393), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5306 (.nQ(w5410), .D(w5479), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5307 (.Z(w5478), .B(w5410), .A(w5415) );
	vdp_xor g5308 (.Z(w6432), .B(w5386), .A(w5415) );
	vdp_xor g5309 (.Z(w5446), .B(w5390), .A(w5415) );
	vdp_xor g5310 (.Z(w6360), .B(w6359), .A(w5415) );
	vdp_sr_bit g5311 (.Q(w6435), .D(w5351), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5312 (.nQ(w6359), .D(w5413), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5313 (.nQ(w6361), .D(w5405), .nC(nDCLK2), .C(DCLK2) );
	vdp_and g5314 (.Z(w5407), .B(w6360), .A(w5416) );
	vdp_and g5315 (.Z(w5408), .B(w6361), .A(DCLK1) );
	vdp_and g5316 (.Z(w5392), .B(w5449), .A(DCLK1) );
	vdp_and g5317 (.Z(w5387), .B(w5446), .A(w5416) );
	vdp_and g5318 (.Z(w5369), .B(w5451), .A(w5450) );
	vdp_and g5319 (.Z(w5370), .B(w81), .A(w5451) );
	vdp_and g5320 (.Z(w5371), .B(w82), .A(w5450) );
	vdp_and g5321 (.Z(w5372), .B(w81), .A(w82) );
	vdp_and g5322 (.Z(w5385), .B(w6432), .A(w82) );
	vdp_and g5323 (.Z(w5404), .B(w5462), .A(DCLK1) );
	vdp_and g5324 (.Z(w5394), .B(w5476), .A(DCLK1) );
	vdp_and g5325 (.Z(w5368), .B(w5478), .A(w5416) );
	vdp_sr_bit g5326 (.Q(w5454), .D(w5457), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5327 (.Q(w5465), .D(w5435), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_not g5328 (.nZ(w5375), .A(w5382) );
	vdp_not g5329 (.nZ(w5380), .A(w123) );
	vdp_not g5330 (.nZ(w5450), .A(w81) );
	vdp_not g5331 (.nZ(w5451), .A(w82) );
	vdp_aoi21 g5332 (.Z(w5405), .B(w5419), .A1(w5406), .A2(w5407) );
	vdp_aoi21 g5333 (.Z(w5388), .B(w5419), .A1(w5389), .A2(w5387) );
	vdp_aoi21 g5334 (.Z(w6394), .B(w5461), .A1(w5384), .A2(w5385) );
	vdp_oai21 g5335 (.Z(w5382), .B(DCLK2), .A1(w5466), .A2(w5465) );
	vdp_aoi21 g5336 (.Z(w6393), .B(w5461), .A1(w5368), .A2(w5411) );
	vdp_not g5337 (.nZ(w5373), .A(w116) );
	vdp_nand g5338 (.Z(w5435), .B(w5473), .A(w5380) );
	vdp_sr_bit g5339 (.Q(w5426), .D(w5482), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5340 (.Q(w5431), .D(w6362), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5341 (.Q(w5442), .D(w6434), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5342 (.Q(w5427), .D(w5444), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5343 (.Q(w5448), .D(w2699), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5344 (.Q(w5452), .D(w5453), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5345 (.Q(w6404), .D(w5469), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5346 (.Q(w5469), .D(w5481), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5347 (.Q(w5484), .D(w5280), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g5348 (.Z(w5481), .B2(w5280), .B1(w5488), .A1(w5487), .A2(w5484) );
	vdp_aon22 g5349 (.Z(w5453), .B2(w5457), .B1(w5488), .A1(w5487), .A2(w5454) );
	vdp_aon22 g5350 (.Z(w5444), .B2(w5332), .B1(w5488), .A1(w5487), .A2(w5445) );
	vdp_aon22 g5351 (.Z(w5482), .B2(w5351), .B1(w5488), .A1(w5487), .A2(w6435) );
	vdp_not g5352 (.nZ(w5425), .A(w5479) );
	vdp_not g5353 (.nZ(w5417), .A(w82) );
	vdp_not g5354 (.nZ(w5422), .A(w5500) );
	vdp_not g5355 (.nZ(w5430), .A(M5) );
	vdp_not g5356 (.nZ(w5433), .A(w5434) );
	vdp_not g5357 (.nZ(w5420), .A(w5493) );
	vdp_not g5358 (.nZ(w5414), .A(w5491) );
	vdp_not g5359 (.nZ(w5463), .A(w5460) );
	vdp_not g5360 (.nZ(w5480), .A(w5468) );
	vdp_not g5361 (.nZ(w5474), .A(w5469) );
	vdp_comp_we g5362 (.nZ(w5488), .A(M5), .Z(w5487) );
	vdp_and g5363 (.Z(w2817), .B(w5427), .A(w5426) );
	vdp_or g5364 (.Z(w6362), .B(w5426), .A(w5430) );
	vdp_or g5365 (.Z(w5436), .B(w5439), .A(w5435) );
	vdp_and g5366 (.Z(w6434), .B(w5427), .A(M5) );
	vdp_and g5367 (.Z(w2699), .B(w5452), .A(M5) );
	vdp_or g5368 (.Z(w5477), .B(w5435), .A(w5467) );
	vdp_not g5369 (.nZ(w5499), .A(SPR_PRIO) );
	vdp_bufif0 g5370 (.A(w6404), .Z(COL[0]), .nE(w5499) );
	vdp_oai21 g5371 (.Z(w5460), .B(DCLK2), .A1(w5436), .A2(w5459) );
	vdp_bufif0 g5372 (.A(w5448), .Z(COL[6]), .nE(w5499) );
	vdp_bufif0 g5373 (.A(w5442), .Z(COL[5]), .nE(w5499) );
	vdp_bufif0 g5374 (.A(w5431), .Z(COL[4]), .nE(w5499) );
	vdp_oai21 g5375 (.Z(w5434), .B(DCLK2), .A1(w5436), .A2(w5421) );
	vdp_oai21 g5376 (.Z(w5500), .B(DCLK2), .A1(w5494), .A2(w5421) );
	vdp_and3 g5377 (.Z(w5421), .B(w5498), .A(w5420), .C(w5497) );
	vdp_and3 g5378 (.Z(w5439), .B(w5498), .A(w5420), .C(w5485) );
	vdp_and3 g5379 (.Z(w5459), .B(w5497), .A(w5486), .C(w5420) );
	vdp_and3 g5380 (.Z(w5467), .B(w5485), .A(w5486), .C(w5420) );
	vdp_or4 g5381 (.Z(w2698), .B(w5490), .A(w5471), .D(w5469), .C(w5470) );
	vdp_and4 g5382 (.Z(w2757), .B(w5470), .A(w5490), .D(w5474), .C(w5471) );
	vdp_and4 g5383 (.Z(w2756), .B(w5470), .A(w5490), .D(w5469), .C(w5471) );
	vdp_oai21 g5384 (.Z(w5468), .B(DCLK2), .A1(w5459), .A2(w5477) );
	vdp_nand3 g5385 (.Z(w5413), .B(w5414), .A(w5425), .C(w5496) );
	vdp_nand3 g5386 (.Z(w5418), .B(w5495), .A(w115), .C(w5417) );
	vdp_nand3 g5387 (.Z(w5458), .B(w81), .A(w115), .C(w5417) );
	vdp_nand g5388 (.Z(w5461), .B(w5458), .A(w5489) );
	vdp_nand g5389 (.Z(w5455), .B(w5492), .A(w5491) );
	vdp_nand g5390 (.Z(w5456), .B(w5425), .A(w5455) );
	vdp_nand g5391 (.Z(w5447), .B(w5414), .A(w5425) );
	vdp_nand g5392 (.Z(w5419), .B(w5418), .A(w5489) );
	vdp_sr_bit g5393 (.Q(w6365), .D(w6364), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5394 (.Q(w6366), .D(w6365), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5395 (.Q(w5565), .D(w6366), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5396 (.Q(w5572), .D(w5565), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5397 (.Q(w5472), .D(w6367), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5398 (.Q(w6433), .D(w5573), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5399 (.Q(w5575), .D(w6471), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5400 (.Q(w5556), .D(w6363), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_dlatch_inv g5401 (.nQ(w5523), .D(w5515), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5402 (.nQ(w5528), .D(w5514), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5403 (.nQ(w5534), .D(w5513), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5404 (.nQ(w5539), .D(w5512), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5405 (.nQ(w5540), .D(w5511), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5406 (.nQ(w5543), .D(w5510), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5407 (.nQ(w5544), .D(w5509), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5408 (.nQ(w5547), .D(w5507), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5409 (.nQ(w5569), .D(w5570), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5410 (.nQ(w5567), .D(w5552), .nC(nDCLK1), .C(DCLK1) );
	vdp_cnt_bit_load g5411 (.Q(w5570), .D(w5571), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1), .R(1'b0), .CI(w6473), .L(w5504), .nL(w5549) );
	vdp_cnt_bit_load g5412 (.Q(w5552), .D(w5551), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1), .R(1'b0), .CI(w5505), .L(w5504), .nL(w5549), .CO(w6473) );
	vdp_aon22 g5413 (.Z(w5437), .B2(w5506), .B1(DB[11]), .A1(w5547), .A2(w5524) );
	vdp_aon22 g5414 (.Z(w5507), .B2(w5508), .B1(w5536), .A1(w5535), .A2(w5527) );
	vdp_aon22 g5415 (.Z(w5440), .B2(w5506), .B1(DB[12]), .A1(w5544), .A2(w5524) );
	vdp_aon22 g5416 (.Z(w5509), .B2(w5508), .B1(w5532), .A1(w5533), .A2(w5527) );
	vdp_aon22 g5417 (.Z(w5441), .B2(w5506), .B1(DB[13]), .A1(w5543), .A2(w5524) );
	vdp_aon22 g5418 (.Z(w5510), .B2(w5508), .B1(w5525), .A1(w5526), .A2(w5527) );
	vdp_aon22 g5419 (.Z(w5443), .B2(w5506), .B1(DB[14]), .A1(w5540), .A2(w5524) );
	vdp_aon22 g5420 (.Z(w5511), .B2(w5508), .B1(w5516), .A1(w5517), .A2(w5527) );
	vdp_aon22 g5421 (.Z(w5424), .B2(w5506), .B1(DB[3]), .A1(w5539), .A2(w5524) );
	vdp_aon22 g5422 (.Z(w5512), .B2(w5508), .B1(w5535), .A1(w5536), .A2(w5527) );
	vdp_aon22 g5423 (.Z(w5428), .B2(w5506), .B1(DB[4]), .A1(w5534), .A2(w5524) );
	vdp_aon22 g5424 (.Z(w5513), .B2(w5508), .B1(w5533), .A1(w5532), .A2(w5527) );
	vdp_aon22 g5425 (.Z(w5429), .B2(w5506), .B1(DB[5]), .A1(w5528), .A2(w5524) );
	vdp_aon22 g5426 (.Z(w5514), .B2(w5508), .B1(w5526), .A1(w5525), .A2(w5527) );
	vdp_aon22 g5427 (.Z(w5432), .B2(w5506), .B1(DB[6]), .A1(w5523), .A2(w5524) );
	vdp_aon22 g5428 (.Z(w5515), .B2(w5508), .B1(w5517), .A1(w5516), .A2(w5527) );
	vdp_slatch g5429 (.Q(w6363), .D(w5559), .nC(w5503), .C(w5560) );
	vdp_dlatch_inv g5430 (.nQ(w5557), .D(w5556), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5431 (.nQ(w5573), .D(w26), .nC(nHCLK1), .C(HCLK1) );
	vdp_xnor g5432 (.Z(w5486), .B(1'b0), .A(w5567) );
	vdp_xor g5433 (.Z(w5548), .B(w5556), .A(w5558) );
	vdp_aon22 g5434 (.Z(w6471), .B2(w5565), .B1(M5), .A1(w5572), .A2(w6472) );
	vdp_not g5435 (.nZ(w5574), .A(w5573) );
	vdp_not g5436 (.nZ(w6472), .A(M5) );
	vdp_not g5437 (.nZ(w5503), .A(w5560) );
	vdp_not g5438 (.nZ(w6364), .A(w5563) );
	vdp_not g5439 (.nZ(w5485), .A(w5557) );
	vdp_not g5440 (.nZ(w5493), .A(w5569) );
	vdp_not g5441 (.nZ(w5505), .A(w5560) );
	vdp_comp_we g5442 (.nZ(w5524), .A(w123), .Z(w5506) );
	vdp_comp_we g5443 (.nZ(w5527), .A(w5548), .Z(w5508) );
	vdp_comp_we g5444 (.nZ(w5549), .A(w5560), .Z(w5504) );
	vdp_and g5445 (.Z(w6367), .B(w6433), .A(w5574) );
	vdp_aoi21 g5446 (.Z(w5563), .B(w25), .A1(M5), .A2(w22) );
	vdp_sr_bit g5447 (.Q(w5558), .D(w5620), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_aon22 g5448 (.Z(w5628), .B2(w5622), .B1(w5621), .A1(w5618), .A2(w5566) );
	vdp_aon22 g5449 (.Z(w5627), .B2(w5622), .B1(w5625), .A1(w5623), .A2(w5566) );
	vdp_aon22 g5450 (.Z(w5624), .B2(w5622), .B1(w5623), .A1(w5625), .A2(w5566) );
	vdp_aon22 g5451 (.Z(w5629), .B2(w5622), .B1(w5618), .A1(w5621), .A2(w5566) );
	vdp_not g5452 (.nZ(w5585), .A(w5621) );
	vdp_not g5453 (.nZ(w5586), .A(w5625) );
	vdp_not g5454 (.nZ(w5591), .A(w5623) );
	vdp_not g5455 (.nZ(w5590), .A(w5618) );
	vdp_not g5456 (.nZ(w5519), .A(w5627) );
	vdp_not g5457 (.nZ(w5520), .A(w5628) );
	vdp_not g5458 (.nZ(w5521), .A(w5629) );
	vdp_not g5459 (.nZ(w5522), .A(w5624) );
	vdp_not g5460 (.nZ(w5564), .A(M5) );
	vdp_comp_we g5461 (.nZ(w5622), .A(w5558), .Z(w5566) );
	vdp_not g5462 (.nZ(w5560), .A(w5619) );
	vdp_not g5463 (.nZ(w5617), .A(w5616) );
	vdp_dlatch_inv g5464 (.nQ(w5616), .D(w5615), .nC(nHCLK1), .C(HCLK1) );
	vdp_aon2222 g5465 (.Z(w5518), .B2(w5520), .B1(w5579), .A1(w5578), .A2(w5519), .D2(w5522), .D1(w5596), .C1(w5595), .C2(w5521) );
	vdp_aon2222 g5466 (.Z(w5568), .B2(w5591), .B1(w5583), .A1(w5590), .A2(w5578), .D2(w5585), .D1(w5587), .C1(w5586), .C2(w5630) );
	vdp_aon2222 g5467 (.Z(w5538), .B2(w5520), .B1(w5584), .A1(w5583), .A2(w5519), .D2(w5522), .D1(w5588), .C1(w5631), .C2(w5521) );
	vdp_aon2222 g5468 (.Z(w5529), .B2(w5591), .B1(w5584), .A1(w5590), .A2(w5579), .D2(w5585), .D1(w5598), .C1(w5586), .C2(w5592) );
	vdp_aon2222 g5469 (.Z(w5546), .B2(w5520), .B1(w5592), .A1(w5630), .A2(w5519), .D2(w5522), .D1(w5594), .C1(w5593), .C2(w5521) );
	vdp_aon2222 g5470 (.Z(w5537), .B2(w5591), .B1(w5631), .A1(w5590), .A2(w5595), .D2(w5585), .D1(w5597), .C1(w5586), .C2(w5593) );
	vdp_aon2222 g5471 (.Z(w6392), .B2(w5520), .B1(w5598), .A1(w5587), .A2(w5519), .D2(w5522), .D1(w5599), .C1(w5597), .C2(w5521) );
	vdp_aon2222 g5472 (.Z(w5541), .B2(w5591), .B1(w5588), .A1(w5590), .A2(w5596), .D2(w5585), .D1(w5599), .C1(w5586), .C2(w5594) );
	vdp_aon2222 g5473 (.Z(w5530), .B2(w5520), .B1(w5601), .A1(w5600), .A2(w5519), .D2(w5522), .D1(w5613), .C1(w5602), .C2(w5521) );
	vdp_aon2222 g5474 (.Z(w5545), .B2(w5591), .B1(w5603), .A1(w5590), .A2(w5600), .D2(w5585), .D1(w5604), .C1(w5586), .C2(w5605) );
	vdp_aon2222 g5475 (.Z(w5542), .B2(w5520), .B1(w5607), .A1(w5603), .A2(w5519), .D2(w5522), .D1(w5606), .C1(w5608), .C2(w5521) );
	vdp_aon2222 g5476 (.Z(w5554), .B2(w5591), .B1(w5607), .A1(w5590), .A2(w5601), .D2(w5585), .D1(w5609), .C1(w5586), .C2(w5610) );
	vdp_aon2222 g5477 (.Z(w5553), .B2(w5520), .B1(w5610), .A1(w5605), .A2(w5519), .D2(w5522), .D1(w5611), .C1(w5612), .C2(w5521) );
	vdp_aon2222 g5478 (.Z(w5555), .B2(w5591), .B1(w5608), .A1(w5590), .A2(w5602), .D2(w5585), .D1(w5614), .C1(w5586), .C2(w5612) );
	vdp_aon2222 g5479 (.Z(w5562), .B2(w5520), .B1(w5609), .A1(w5604), .A2(w5519), .D2(w5522), .D1(w5626), .C1(w5614), .C2(w5521) );
	vdp_aon2222 g5480 (.Z(w5561), .B2(w5591), .B1(w5606), .A1(w5590), .A2(w5613), .D2(w5585), .D1(w5626), .C1(w5586), .C2(w5611) );
	vdp_aoi22 g5481 (.Z(w5516), .B2(w5577), .B1(w5518), .A1(w5531), .A2(w5568) );
	vdp_aoi22 g5482 (.Z(w5525), .B2(w5577), .B1(w5530), .A1(w5531), .A2(w5529) );
	vdp_aoi22 g5483 (.Z(w5532), .B2(w5577), .B1(w5538), .A1(w5531), .A2(w5537) );
	vdp_aoi22 g5484 (.Z(w5536), .B2(w5577), .B1(w5542), .A1(w5531), .A2(w5541) );
	vdp_aoi22 g5485 (.Z(w5517), .B2(w5577), .B1(w5546), .A1(w5531), .A2(w5545) );
	vdp_aoi22 g5486 (.Z(w5526), .B2(w5577), .B1(w5553), .A1(w5531), .A2(w5554) );
	vdp_aoi22 g5487 (.Z(w5533), .B2(w5577), .B1(w6392), .A1(w5531), .A2(w5555) );
	vdp_aoi22 g5488 (.Z(w5535), .B2(w5577), .B1(w5562), .A1(w5531), .A2(w5561) );
	vdp_nand g5489 (.Z(w5619), .B(w5617), .A(HCLK2) );
	vdp_nor g5490 (.Z(w5577), .B(w5564), .A(w5472) );
	vdp_nor g5491 (.Z(w5531), .B(M5), .A(w5472) );
	vdp_sr_bit g5492 (.Q(w5621), .D(w5625), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5493 (.Q(w5625), .D(w5623), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5494 (.Q(w5623), .D(w5618), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5495 (.Q(w5618), .D(w5619), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_dlatch_inv g5496 (.nQ(w5466), .D(w5621), .nC(nDCLK1), .C(DCLK1) );
	vdp_comp_str g5497 (.nZ(w5582), .A(w5633), .Z(w5635) );
	vdp_comp_str g5498 (.nZ(w5581), .A(w5633), .Z(w5638) );
	vdp_comp_str g5499 (.nZ(w5589), .A(w5633), .Z(w5639) );
	vdp_comp_str g5500 (.nZ(w5580), .A(w5633), .Z(w5634) );
	vdp_slatch g5501 (.D(w5648), .Q(w5578), .nC(w5580), .C(w5634) );
	vdp_slatch g5502 (.D(w6497), .Q(w5579), .nC(w5589), .C(w5639) );
	vdp_slatch g5503 (.D(w6496), .Q(w5595), .nC(w5581), .C(w5638) );
	vdp_slatch g5504 (.D(w6495), .Q(w5596), .nC(w5582), .C(w5635) );
	vdp_slatch g5505 (.D(w5647), .Q(w5583), .nC(w5580), .C(w5634) );
	vdp_slatch g5506 (.D(w6494), .Q(w5584), .nC(w5589), .C(w5639) );
	vdp_slatch g5507 (.D(w6493), .Q(w5631), .nC(w5581), .C(w5638) );
	vdp_slatch g5508 (.D(w6492), .Q(w5588), .nC(w5582), .C(w5635) );
	vdp_slatch g5509 (.D(w5646), .Q(w5630), .nC(w5580), .C(w5634) );
	vdp_slatch g5510 (.D(w6491), .Q(w5592), .nC(w5589), .C(w5639) );
	vdp_slatch g5511 (.D(w6490), .Q(w5593), .nC(w5581), .C(w5638) );
	vdp_slatch g5512 (.D(w6489), .Q(w5594), .nC(w5582), .C(w5635) );
	vdp_slatch g5513 (.D(w5645), .Q(w5587), .nC(w5580), .C(w5634) );
	vdp_slatch g5514 (.D(w6488), .Q(w5598), .nC(w5589), .C(w5639) );
	vdp_slatch g5515 (.D(w6487), .Q(w5597), .nC(w5581), .C(w5638) );
	vdp_slatch g5516 (.D(w6486), .Q(w5599), .nC(w5582), .C(w5635) );
	vdp_slatch g5517 (.D(w5644), .Q(w5600), .nC(w5580), .C(w5634) );
	vdp_slatch g5518 (.D(w6485), .Q(w5601), .nC(w5589), .C(w5639) );
	vdp_slatch g5519 (.D(w6484), .Q(w5602), .nC(w5581), .C(w5638) );
	vdp_slatch g5520 (.D(w6483), .Q(w5613), .nC(w5582), .C(w5635) );
	vdp_slatch g5521 (.D(w5643), .Q(w5603), .nC(w5580), .C(w5634) );
	vdp_slatch g5522 (.D(w6482), .Q(w5607), .nC(w5589), .C(w5639) );
	vdp_slatch g5523 (.D(w6481), .Q(w5608), .nC(w5581), .C(w5638) );
	vdp_slatch g5524 (.D(w6480), .Q(w5606), .nC(w5582), .C(w5635) );
	vdp_slatch g5525 (.D(w5642), .Q(w5605), .nC(w5580), .C(w5634) );
	vdp_slatch g5526 (.D(w6479), .Q(w5610), .nC(w5589), .C(w5639) );
	vdp_slatch g5527 (.D(w6478), .Q(w5612), .nC(w5581), .C(w5638) );
	vdp_slatch g5528 (.D(w6477), .Q(w5611), .nC(w5582), .C(w5635) );
	vdp_slatch g5529 (.D(w5641), .Q(w5604), .nC(w5580), .C(w5634) );
	vdp_slatch g5530 (.D(w6476), .Q(w5609), .nC(w5589), .C(w5639) );
	vdp_slatch g5531 (.D(w6475), .Q(w5614), .nC(w5581), .C(w5638) );
	vdp_slatch g5532 (.D(w6474), .nC(w5582), .C(w5635), .Q(w5626) );
	vdp_sr_bit g5533 (.Q(w5649), .D(w5650), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g5534 (.Q(w6368), .D(w5649), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g5535 (.Q(w5663), .D(w6368), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_comp_str g5536 (.nZ(w5653), .A(w5664), .Z(w5640) );
	vdp_comp_str g5537 (.nZ(w5656), .A(w5664), .Z(w5637) );
	vdp_comp_str g5538 (.nZ(w5658), .A(w5664), .Z(w5636) );
	vdp_dlatch_inv g5539 (.nQ(w5650), .D(w5659), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g5540 (.Z(w5633), .B(DCLK2), .A(w5663) );
	vdp_and g5541 (.Z(w5664), .B(DCLK2), .A(w5649) );
	vdp_and g5542 (.Z(w5665), .B(DCLK2), .A(w5650) );
	vdp_slatch g5543 (.Q(w6476), .D(w6500), .nC(w5653), .C(w5640) );
	vdp_slatch g5544 (.Q(w6475), .D(w6499), .nC(w5656), .C(w5637) );
	vdp_slatch g5545 (.Q(w6474), .D(w6498), .nC(w5658), .C(w5636) );
	vdp_slatch g5546 (.Q(w6479), .D(w6503), .nC(w5653), .C(w5640) );
	vdp_slatch g5547 (.Q(w6478), .D(w6502), .nC(w5656), .C(w5637) );
	vdp_slatch g5548 (.Q(w6477), .D(w6501), .nC(w5658), .C(w5636) );
	vdp_slatch g5549 (.Q(w6482), .D(w6506), .nC(w5653), .C(w5640) );
	vdp_slatch g5550 (.Q(w6481), .D(w6505), .nC(w5656), .C(w5637) );
	vdp_slatch g5551 (.Q(w6480), .D(w6504), .nC(w5658), .C(w5636) );
	vdp_slatch g5552 (.Q(w6485), .D(w6509), .nC(w5653), .C(w5640) );
	vdp_slatch g5553 (.Q(w6484), .D(w6508), .nC(w5656), .C(w5637) );
	vdp_slatch g5554 (.Q(w6483), .D(w6507), .nC(w5658), .C(w5636) );
	vdp_slatch g5555 (.Q(w6488), .D(w6512), .nC(w5653), .C(w5640) );
	vdp_slatch g5556 (.Q(w6487), .D(w6511), .nC(w5656), .C(w5637) );
	vdp_slatch g5557 (.Q(w6486), .D(w6510), .nC(w5658), .C(w5636) );
	vdp_slatch g5558 (.Q(w6491), .D(w6515), .nC(w5653), .C(w5640) );
	vdp_slatch g5559 (.Q(w6490), .D(w6514), .nC(w5656), .C(w5637) );
	vdp_slatch g5560 (.Q(w6489), .D(w6513), .nC(w5658), .C(w5636) );
	vdp_slatch g5561 (.Q(w6494), .D(w6518), .nC(w5653), .C(w5640) );
	vdp_slatch g5562 (.Q(w6493), .D(w6517), .nC(w5656), .C(w5637) );
	vdp_slatch g5563 (.Q(w6492), .D(w6516), .nC(w5658), .C(w5636) );
	vdp_slatch g5564 (.Q(w6497), .D(w6521), .nC(w5653), .C(w5640) );
	vdp_slatch g5565 (.Q(w6496), .D(w6520), .nC(w5656), .C(w5637) );
	vdp_slatch g5566 (.Q(w6495), .D(w6519), .nC(w5658), .C(w5636) );
	vdp_sr_bit g5567 (.Q(w5662), .D(w5661), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_dlatch_inv g5568 (.nQ(w5661), .D(w5660), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g5569 (.Z(w5672), .B(w5661), .A(DCLK2) );
	vdp_nand g5570 (.Z(w5660), .B(w5565), .A(HCLK1) );
	vdp_nand g5571 (.Z(w5659), .B(w5575), .A(HCLK1) );
	vdp_and g5572 (.Z(w5671), .B(w5662), .A(DCLK2) );
	vdp_comp_str g5573 (.nZ(w5657), .A(w5672), .Z(w5670) );
	vdp_comp_str g5574 (.nZ(w5655), .A(w5671), .Z(w5669) );
	vdp_comp_str g5575 (.nZ(w5654), .A(w5665), .Z(w5668) );
	vdp_comp_str g5576 (.nZ(w5652), .A(w5664), .Z(w5667) );
	vdp_slatch g5577 (.D(S[7]), .Q(w5648), .nC(w5652), .C(w5667) );
	vdp_slatch g5578 (.D(S[7]), .Q(w6521), .nC(w5654), .C(w5668) );
	vdp_slatch g5579 (.D(S[7]), .Q(w6520), .nC(w5655), .C(w5669) );
	vdp_slatch g5580 (.D(S[7]), .Q(w6519), .nC(w5657), .C(w5670) );
	vdp_slatch g5581 (.D(S[5]), .Q(w5647), .nC(w5652), .C(w5667) );
	vdp_slatch g5582 (.D(S[5]), .Q(w6518), .nC(w5654), .C(w5668) );
	vdp_slatch g5583 (.D(S[5]), .Q(w6517), .nC(w5655), .C(w5669) );
	vdp_slatch g5584 (.D(S[5]), .Q(w6516), .nC(w5657), .C(w5670) );
	vdp_slatch g5585 (.D(S[3]), .Q(w5646), .nC(w5652), .C(w5667) );
	vdp_slatch g5586 (.D(S[3]), .Q(w6515), .nC(w5654), .C(w5668) );
	vdp_slatch g5587 (.D(S[3]), .Q(w6514), .nC(w5655), .C(w5669) );
	vdp_slatch g5588 (.D(S[3]), .Q(w6513), .nC(w5657), .C(w5670) );
	vdp_slatch g5589 (.D(S[1]), .Q(w5645), .nC(w5652), .C(w5667) );
	vdp_slatch g5590 (.D(S[1]), .Q(w6512), .nC(w5654), .C(w5668) );
	vdp_slatch g5591 (.D(S[1]), .Q(w6511), .nC(w5655), .C(w5669) );
	vdp_slatch g5592 (.D(S[1]), .Q(w6510), .nC(w5657), .C(w5670) );
	vdp_slatch g5593 (.D(S[6]), .Q(w5644), .nC(w5652), .C(w5667) );
	vdp_slatch g5594 (.D(S[6]), .Q(w6509), .nC(w5654), .C(w5668) );
	vdp_slatch g5595 (.D(S[6]), .Q(w6508), .nC(w5655), .C(w5669) );
	vdp_slatch g5596 (.D(S[6]), .Q(w6507), .nC(w5657), .C(w5670) );
	vdp_slatch g5597 (.D(S[4]), .Q(w5643), .nC(w5652), .C(w5667) );
	vdp_slatch g5598 (.D(S[4]), .Q(w6506), .nC(w5654), .C(w5668) );
	vdp_slatch g5599 (.D(S[4]), .Q(w6505), .nC(w5655), .C(w5669) );
	vdp_slatch g5600 (.D(S[4]), .Q(w6504), .nC(w5657), .C(w5670) );
	vdp_slatch g5601 (.D(S[2]), .Q(w5642), .nC(w5652), .C(w5667) );
	vdp_slatch g5602 (.D(S[2]), .Q(w6503), .nC(w5654), .C(w5668) );
	vdp_slatch g5603 (.D(S[2]), .Q(w6502), .nC(w5655), .C(w5669) );
	vdp_slatch g5604 (.D(S[2]), .Q(w6501), .nC(w5657), .C(w5670) );
	vdp_slatch g5605 (.D(S[0]), .Q(w5641), .nC(w5652), .C(w5667) );
	vdp_slatch g5606 (.D(S[0]), .Q(w6500), .nC(w5654), .C(w5668) );
	vdp_slatch g5607 (.D(S[0]), .Q(w6499), .nC(w5655), .C(w5669) );
	vdp_slatch g5608 (.D(S[0]), .nC(w5657), .C(w5670), .Q(w6498) );
	vdp_aon21_sr g5609 (.Q(w5727), .A1(w5320), .A2(w6682), .B(w6408), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5610 (.Q(w6408), .A1(w5299), .A2(w6682), .B(w6409), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5611 (.Q(w6409), .A1(w5297), .A2(w6682), .B(w6410), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5612 (.Q(w6410), .A1(w5687), .A2(w6682), .B(w6411), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5613 (.Q(w6411), .A1(w5716), .A2(w6682), .B(w6412), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5614 (.Q(w6412), .A1(w5679), .A2(w6682), .B(w6407), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5615 (.Q(w6407), .A1(w5680), .A2(w6682), .B(w6406), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5616 (.Q(w6406), .A1(w5681), .A2(w6682), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5617 (.Q(w6419), .A1(w5683), .A2(w6683), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5618 (.Q(w6418), .A1(w5684), .A2(w6683), .B(w6419), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5619 (.Q(w6417), .A1(w5697), .A2(w6683), .B(w6418), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5620 (.Q(w6416), .A1(w5685), .A2(w6683), .B(w6417), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5621 (.Q(w6415), .A1(w5686), .A2(w6683), .B(w6416), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5622 (.Q(w6414), .A1(w5298), .A2(w6683), .B(w6415), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5623 (.Q(w6413), .A1(w5300), .A2(w6683), .B(w6414), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5624 (.Q(w5731), .A1(w5319), .A2(w6683), .B(w6413), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5625 (.Q(w5736), .A1(w5693), .A2(w6684), .B(w6426), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5626 (.Q(w6426), .A1(w5689), .A2(w6684), .B(w6425), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5627 (.Q(w6425), .A1(w5688), .A2(w6684), .B(w6424), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5628 (.Q(w6424), .A1(w5695), .A2(w6684), .B(w6423), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5629 (.Q(w6423), .A1(w5696), .A2(w6684), .B(w6422), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5630 (.Q(w6422), .A1(w5698), .A2(w6684), .B(w6421), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5631 (.Q(w6421), .A1(w5710), .A2(w6684), .B(w6420), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5632 (.Q(w6420), .A1(w5711), .A2(w6684), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_or4 g5633 (.Z(w5719), .B(w5716), .A(w5281), .C(w5685), .D(w5696) );
	vdp_or4 g5634 (.Z(w5363), .B(w5687), .A(w5359), .C(w5686), .D(w5695) );
	vdp_aon22 g5635 (.Z(w5706), .B2(w4497), .B1(w5713), .A1(w5741), .A2(DB[0]) );
	vdp_aon22 g5636 (.Z(w5705), .B2(w4498), .B1(w5713), .A1(w5741), .A2(DB[1]) );
	vdp_aon22 g5637 (.Z(w5704), .B2(w4506), .B1(w5713), .A1(w5741), .A2(DB[2]) );
	vdp_aon22 g5638 (.Z(w5703), .B2(w4497), .B1(w5713), .A1(w5741), .A2(DB[8]) );
	vdp_aon22 g5639 (.Z(w5702), .B2(w4498), .B1(w5713), .A1(w5741), .A2(DB[9]) );
	vdp_aon22 g5640 (.Z(w5701), .B2(w4506), .B1(w5713), .A1(w5741), .A2(DB[10]) );
	vdp_or4 g5641 (.Z(w5728), .B(w5677), .A(w5678), .C(w5682), .D(w5715) );
	vdp_or4 g5642 (.Z(w5720), .B(w5690), .A(w5718), .C(w5691), .D(w5717) );
	vdp_or4 g5643 (.Z(w5735), .B(w5680), .A(w5283), .C(w5684), .D(w5710) );
	vdp_or4 g5644 (.Z(w5732), .B(w5697), .A(w5698), .C(w5679), .D(w5282) );
	vdp_or4 g5645 (.Z(w5742), .B(w5692), .A(w5694), .C(w5700), .D(w5699) );
	vdp_or4 g5646 (.Z(w5733), .B(w5708), .A(w5709), .C(w5712), .D(w5707) );
	vdp_or4 g5647 (.Z(w5744), .B(w5681), .A(w5284), .C(w5683), .D(w5711) );
	vdp_comp_we g5648 (.nZ(w5713), .A(w123), .Z(w5741) );
	vdp_not g5649 (.nZ(w6682), .A(w5344) );
	vdp_not g5650 (.nZ(w6683), .A(w5344) );
	vdp_not g5651 (.nZ(w6684), .A(w5344) );
	vdp_slatch g5652 (.Q(w5717), .D(w5759), .nC(w5725), .C(w5758) );
	vdp_comp_str g5653 (.nZ(w5725), .A(w5375), .Z(w5758) );
	vdp_slatch g5654 (.Q(w5691), .D(w5761), .nC(w5725), .C(w5758) );
	vdp_slatch g5655 (.Q(w5690), .D(w5762), .nC(w5725), .C(w5758) );
	vdp_slatch g5656 (.Q(w5718), .D(w5763), .nC(w5725), .C(w5758) );
	vdp_slatch g5657 (.Q(w5678), .D(w5764), .nC(w5725), .C(w5758) );
	vdp_slatch g5658 (.Q(w5677), .D(w5766), .nC(w5725), .C(w5758) );
	vdp_slatch g5659 (.Q(w5682), .D(w5767), .nC(w5725), .C(w5758) );
	vdp_slatch g5660 (.Q(w5715), .D(w5768), .nC(w5725), .C(w5758) );
	vdp_slatch g5661 (.Q(w5707), .D(w5777), .nC(w5739), .C(w5776) );
	vdp_comp_str g5662 (.nZ(w5739), .A(w5375), .Z(w5776) );
	vdp_slatch g5663 (.Q(w5712), .D(w5779), .nC(w5739), .C(w5776) );
	vdp_slatch g5664 (.Q(w5708), .D(w5780), .nC(w5739), .C(w5776) );
	vdp_slatch g5665 (.Q(w5709), .D(w5781), .nC(w5739), .C(w5776) );
	vdp_slatch g5666 (.Q(w5694), .D(w5782), .nC(w5739), .C(w5776) );
	vdp_slatch g5667 (.Q(w5692), .D(w5784), .nC(w5739), .C(w5776) );
	vdp_slatch g5668 (.Q(w5700), .D(w5785), .nC(w5739), .C(w5776) );
	vdp_slatch g5669 (.Q(w5699), .D(w5786), .nC(w5739), .C(w5776) );
	vdp_comp_we g5670 (.nZ(w5722), .A(1'b0), .Z(w5361) );
	vdp_aon22 g5671 (.Z(w5788), .B2(w5722), .B1(w5743), .A1(w5742), .A2(w5361) );
	vdp_not g5672 (.nZ(w5344), .A(w4508) );
	vdp_not g5673 (.nZ(w5743), .A(w5744) );
	vdp_not g5674 (.nZ(w5734), .A(w5735) );
	vdp_not g5675 (.nZ(w5730), .A(w5732) );
	vdp_not g5676 (.nZ(w5721), .A(w5719) );
	vdp_and3 g5677 (.Z(w5748), .B(w5747), .A(w5720), .C(w5719) );
	vdp_aon22 g5678 (.Z(w5756), .B2(w5722), .B1(w5721), .A1(w5720), .A2(w5361) );
	vdp_notif0 g5679 (.A(w5723), .nZ(DB[4]), .nE(w5724) );
	vdp_aon2222 g5680 (.Z(w5723), .B2(w5716), .B1(w5754), .A1(w5755), .A2(w5680), .D2(w5320), .D1(w5752), .C1(w5753), .C2(w5297) );
	vdp_notif0 g5681 (.A(w5726), .nZ(DB[12]), .nE(w5724) );
	vdp_aon2222 g5682 (.Z(w5726), .B2(w5679), .B1(w5754), .A1(w5755), .A2(w5681), .D2(w5299), .D1(w5752), .C1(w5753), .C2(w5687) );
	vdp_notif0 g5683 (.A(w6403), .nZ(DB[13]), .nE(w5724) );
	vdp_aon2222 g5684 (.Z(w6403), .B2(w5697), .B1(w5754), .A1(w5755), .A2(w5683), .D2(w5300), .D1(w5752), .C1(w5753), .C2(w5686) );
	vdp_notif0 g5685 (.A(w5729), .nZ(DB[5]), .nE(w5724) );
	vdp_aon2222 g5686 (.Z(w5729), .B2(w5685), .B1(w5754), .A1(w5755), .A2(w5684), .D2(w5319), .D1(w5752), .C1(w5753), .C2(w5298) );
	vdp_notif0 g5687 (.A(w5738), .nZ(DB[14]), .nE(w5724) );
	vdp_aon2222 g5688 (.Z(w5738), .B2(w5698), .B1(w5754), .A1(w5755), .A2(w5711), .D2(w5689), .D1(w5752), .C1(w5753), .C2(w5695) );
	vdp_notif0 g5689 (.A(w5737), .nZ(DB[6]), .nE(w5724) );
	vdp_aon2222 g5690 (.Z(w5737), .B2(w5696), .B1(w5754), .A1(w5755), .A2(w5710), .D2(w5693), .D1(w5752), .C1(w5753), .C2(w5688) );
	vdp_aon22 g5691 (.Z(w5769), .B2(w5722), .B1(w5730), .A1(w5728), .A2(w5361) );
	vdp_aon22 g5692 (.Z(w5772), .B2(w5722), .B1(w5734), .A1(w5733), .A2(w5361) );
	vdp_and3 g5693 (.Z(w5750), .B(w5771), .A(w5728), .C(w5732) );
	vdp_and3 g5694 (.Z(w5751), .B(w5773), .A(w5733), .C(w5735) );
	vdp_and3 g5695 (.Z(w5749), .B(w5787), .A(w5742), .C(w5744) );
	vdp_not g5696 (.nZ(w5724), .A(w116) );
	vdp_slatch g5697 (.Q(w5782), .D(w5437), .nC(w5818), .C(w5783) );
	vdp_slatch g5698 (.Q(w5784), .D(w5440), .nC(w5818), .C(w5783) );
	vdp_slatch g5699 (.Q(w5785), .D(w5441), .nC(w5818), .C(w5783) );
	vdp_slatch g5700 (.Q(w5786), .D(w5443), .nC(w5818), .C(w5783) );
	vdp_comp_str g5701 (.nZ(w5818), .A(w5819), .Z(w5783) );
	vdp_slatch g5702 (.Q(w5777), .D(w5424), .nC(w5813), .C(w5778) );
	vdp_slatch g5703 (.Q(w5779), .D(w5428), .nC(w5813), .C(w5778) );
	vdp_slatch g5704 (.Q(w5780), .D(w5429), .nC(w5813), .C(w5778) );
	vdp_slatch g5705 (.Q(w5781), .D(w5432), .nC(w5813), .C(w5778) );
	vdp_comp_str g5706 (.nZ(w5813), .A(w5817), .Z(w5778) );
	vdp_slatch g5707 (.Q(w5764), .D(w5437), .nC(w5800), .C(w5765) );
	vdp_slatch g5708 (.Q(w5766), .D(w5440), .nC(w5800), .C(w5765) );
	vdp_slatch g5709 (.Q(w5767), .D(w5441), .nC(w5800), .C(w5765) );
	vdp_slatch g5710 (.Q(w5768), .D(w5443), .nC(w5800), .C(w5765) );
	vdp_comp_str g5711 (.nZ(w5800), .A(w6679), .Z(w5765) );
	vdp_slatch g5712 (.Q(w5759), .D(w5424), .nC(w5799), .C(w5760) );
	vdp_slatch g5713 (.Q(w5761), .D(w5428), .nC(w5799), .C(w5760) );
	vdp_slatch g5714 (.Q(w5762), .D(w5429), .nC(w5799), .C(w5760) );
	vdp_slatch g5715 (.Q(w5763), .D(w5432), .nC(w5799), .C(w5760) );
	vdp_comp_str g5716 (.nZ(w5799), .A(w5797), .Z(w5760) );
	vdp_dlatch_inv g5717 (.nQ(w6402), .D(w5792), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5718 (.Z(w5794), .B(w5415), .A(w6402) );
	vdp_sr_bit g5719 (.Q(w121), .D(w6400), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g5720 (.Q(w5791), .D(w5727), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5721 (.nQ(w5796), .D(w5757), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5722 (.nQ(w6395), .D(w5770), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5723 (.nQ(w6397), .D(w5806), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5724 (.Z(w6396), .B(w6397), .A(w5415) );
	vdp_sr_bit g5725 (.Q(w6405), .D(w5731), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5726 (.nQ(w5774), .D(w6677), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5727 (.Z(w6398), .B(w5774), .A(w5415) );
	vdp_sr_bit g5728 (.Q(w5810), .D(w5736), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5729 (.nQ(w5807), .D(w6401), .nC(nDCLK2), .C(DCLK2) );
	vdp_not g5730 (.nZ(w5823), .A(w5415) );
	vdp_not g5731 (.nZ(w5775), .A(w82) );
	vdp_not g5732 (.nZ(w5811), .A(w81) );
	vdp_dlatch_inv g5733 (.nQ(w5821), .D(w6399), .nC(nDCLK2), .C(DCLK2) );
	vdp_and g5734 (.Z(w5787), .B(w5823), .A(w5416) );
	vdp_aoi21 g5735 (.Z(w6399), .B(w5808), .A1(w5788), .A2(w5787) );
	vdp_and g5736 (.Z(w5674), .B(w5821), .A(DCLK1) );
	vdp_and g5737 (.Z(w5675), .B(w5807), .A(DCLK1) );
	vdp_and g5738 (.Z(w5773), .B(w6398), .A(w5416) );
	vdp_aoi21 g5739 (.Z(w6401), .B(w5808), .A1(w5772), .A2(w5773) );
	vdp_and g5740 (.Z(w5771), .B(w6396), .A(w5416) );
	vdp_aoi21 g5741 (.Z(w5770), .B(w5795), .A1(w5769), .A2(w5771) );
	vdp_and g5742 (.Z(w5747), .B(w5416), .A(w5794) );
	vdp_aoi21 g5743 (.Z(w5757), .B(w5795), .A1(w5756), .A2(w5747) );
	vdp_and g5744 (.Z(w5714), .B(DCLK1), .A(w5796) );
	vdp_and g5745 (.Z(w5676), .B(w6395), .A(DCLK1) );
	vdp_and g5746 (.Z(w5752), .B(w5775), .A(w5811) );
	vdp_and g5747 (.Z(w5754), .B(w82), .A(w5811) );
	vdp_and g5748 (.Z(w5753), .B(w5775), .A(w81) );
	vdp_and g5749 (.Z(w5755), .B(w82), .A(w81) );
	vdp_or8 g5750 (.Z(w6400), .B(w5748), .A(w5409), .C(w5749), .D(w5789), .F(w5751), .E(w5746), .G(w5393), .H(w5750) );
	vdp_sr_bit g5751 (.Q(w5471), .D(w5829), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5752 (.Q(w5793), .D(w5471), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5753 (.Q(w5470), .D(w5805), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5754 (.Q(w5824), .D(w5470), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5755 (.Q(w5490), .D(w6384), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5756 (.Q(w5812), .D(w5490), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_comp_we g5757 (.nZ(w5827), .A(M5), .Z(w5826) );
	vdp_not g5758 (.nZ(w5819), .A(w5820) );
	vdp_or g5759 (.Z(w5494), .B(w5822), .A(w5435) );
	vdp_and3 g5760 (.Z(w5822), .B(w5486), .A(w5493), .C(w5485) );
	vdp_and3 g5761 (.Z(w5815), .B(w5486), .A(w5493), .C(w5497) );
	vdp_and3 g5762 (.Z(w6677), .B(w5491), .A(w5479), .C(w5492) );
	vdp_and3 g5763 (.Z(w5802), .B(w5498), .A(w5493), .C(w5485) );
	vdp_and3 g5764 (.Z(w5804), .B(w5498), .A(w5493), .C(w5497) );
	vdp_aoi21 g5765 (.Z(w5792), .B(w5425), .A1(w5414), .A2(w5496) );
	vdp_aon22 g5766 (.Z(w5829), .B2(w5727), .B1(w5827), .A1(w5826), .A2(w5791) );
	vdp_aon22 g5767 (.Z(w5805), .B2(w5731), .B1(w5827), .A1(w5826), .A2(w6405) );
	vdp_aon22 g5768 (.Z(w6384), .B2(w5736), .B1(w5827), .A1(w5826), .A2(w5810) );
	vdp_bufif0 g5769 (.A(w5824), .Z(COL[2]), .nE(w5828) );
	vdp_oai21 g5770 (.Z(w5803), .B(DCLK2), .A1(w5816), .A2(w5804) );
	vdp_and g5771 (.Z(w5806), .B(w5491), .A(w5479) );
	vdp_or g5772 (.Z(w5816), .B(w5802), .A(w5435) );
	vdp_bufif0 g5773 (.A(w5812), .Z(COL[3]), .nE(w5828) );
	vdp_oai21 g5774 (.Z(w5814), .B(DCLK2), .A1(w5816), .A2(w5815) );
	vdp_oai21 g5775 (.Z(w5820), .B(DCLK2), .A1(w5815), .A2(w5494) );
	vdp_not g5776 (.nZ(w5497), .A(w5485) );
	vdp_not g5777 (.nZ(w5817), .A(w5814) );
	vdp_not g5778 (.nZ(w5495), .A(w81) );
	vdp_not g5779 (.nZ(w5498), .A(w5486) );
	vdp_not g5780 (.nZ(w6679), .A(w5803) );
	vdp_not g5781 (.nZ(w5496), .A(w5492) );
	vdp_not g5782 (.nZ(w5797), .A(w5798) );
	vdp_bufif0 g5783 (.A(w5793), .Z(COL[1]), .nE(w5828) );
	vdp_oai21 g5784 (.Z(w5798), .B(DCLK2), .A1(w5477), .A2(w5804) );
	vdp_not g5785 (.nZ(w5828), .A(SPR_PRIO) );
	vdp_nand3 g5786 (.Z(w5801), .B(w115), .A(w82), .C(w5495) );
	vdp_nand g5787 (.Z(w5795), .B(w5489), .A(w5801) );
	vdp_nand3 g5788 (.Z(w5809), .B(w115), .A(w82), .C(w81) );
	vdp_nand g5789 (.Z(w5808), .B(w5489), .A(w5809) );
	vdp_sr_bit g5790 (.Q(w5856), .D(w5897), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5791 (.Q(w5857), .D(w5895), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5792 (.Q(w5854), .D(w5902), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5793 (.Q(w5855), .D(w5894), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5794 (.Z(w4503), .B2(w5856), .B1(w5891), .A1(w5890), .A2(w80), .C1(w5845), .C2(w5857) );
	vdp_aon222 g5795 (.Z(w4502), .B2(w5854), .B1(w5891), .A1(w5890), .A2(w79), .C1(w5845), .C2(w5855) );
	vdp_sr_bit g5796 (.Q(w5852), .D(w5901), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5797 (.Q(w5853), .D(w5893), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5798 (.Z(w4501), .B2(w5852), .B1(w5891), .A1(w5890), .A2(w78), .C1(w5845), .C2(w5853) );
	vdp_sr_bit g5799 (.Q(w5850), .D(w5900), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5800 (.Q(w5851), .D(w5892), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5801 (.Z(w4500), .B2(w5850), .B1(w5891), .A1(w5890), .A2(w77), .C1(w5845), .C2(w5851) );
	vdp_sr_bit g5802 (.Q(w5846), .D(w5899), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5803 (.Q(w5849), .D(w5903), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5804 (.Z(w4499), .B2(w5846), .B1(w5891), .A1(w5890), .A2(w76), .C1(w5845), .C2(w5849) );
	vdp_sr_bit g5805 (.Q(w5847), .D(w5898), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5806 (.Q(w5848), .D(w5889), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5807 (.Z(w4504), .B2(w5847), .B1(w5891), .A1(w5890), .A2(w75), .C1(w5845), .C2(w5848) );
	vdp_sr_bit g5808 (.Q(w5479), .D(w6656), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_slatch g5809 (.Q(w6656), .D(w5571), .nC(w5881), .C(w5842) );
	vdp_sr_bit g5810 (.Q(w5491), .D(w6654), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_slatch g5811 (.Q(w6654), .D(w5551), .nC(w5881), .C(w5842) );
	vdp_sr_bit g5812 (.Q(w5492), .D(w6655), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_slatch g5813 (.Q(w6655), .D(w5559), .nC(w5881), .C(w5842) );
	vdp_sr_bit g5814 (.Q(w5858), .D(w26), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5815 (.Q(w5841), .D(w5858), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5816 (.Q(w5840), .D(w5886), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5817 (.Q(w5874), .D(w5884), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5818 (.Q(w5873), .D(w5883), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5819 (.Q(w5837), .D(w4508), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5820 (.Q(w5836), .D(w5869), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5821 (.Q(w5864), .D(w6429), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5822 (.Q(w6429), .D(w5905), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_xor g5823 (.Z(w5866), .B(w5864), .A(w5865) );
	vdp_dlatch_inv g5824 (.nQ(w5835), .D(w5869), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5825 (.nQ(w5867), .D(w5866), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5826 (.nQ(w5838), .D(w5839), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5827 (.nQ(w5872), .D(w5871), .nC(nHCLK1), .C(HCLK1) );
	vdp_comp_str g5828 (.nZ(w5881), .A(w5878), .Z(w5842) );
	vdp_oai21 g5829 (.Z(w6428), .B(w5868), .A1(w5905), .A2(w5864) );
	vdp_and g5830 (.Z(w4497), .B(w5862), .A(w5834) );
	vdp_not g5831 (.nZ(w5415), .A(w5867) );
	vdp_not g5832 (.nZ(w5869), .A(w6428) );
	vdp_and g5833 (.Z(w4498), .B(w5861), .A(w5834) );
	vdp_and g5834 (.Z(w4506), .B(w5860), .A(w5834) );
	vdp_or g5835 (.Z(w5870), .B(w5836), .A(w5869) );
	vdp_not g5836 (.nZ(w5888), .A(w123) );
	vdp_not g5837 (.nZ(w4508), .A(w5871) );
	vdp_not g5838 (.nZ(w5904), .A(M5) );
	vdp_not g5839 (.nZ(w5891), .A(w6647) );
	vdp_not g5840 (.nZ(w5843), .A(w5842) );
	vdp_not g5841 (.nZ(w5890), .A(w5888) );
	vdp_not g5842 (.nZ(w5845), .A(w5844) );
	vdp_or4 g5843 (.Z(w4505), .B(w4508), .A(w123), .C(w5837), .D(w5870) );
	vdp_or4 g5844 (.Z(w5871), .B(w5874), .A(w5834), .C(w5840), .D(w5873) );
	vdp_nand g5845 (.Z(w5839), .B(w5872), .A(HCLK2) );
	vdp_nand g5846 (.Z(w5489), .B(w5888), .A(w5838) );
	vdp_nor g5847 (.Z(w5416), .B(w5835), .A(w123) );
	vdp_nand g5848 (.Z(w5844), .B(w5888), .A(w5843) );
	vdp_nand g5849 (.Z(w6647), .B(w5888), .A(w5834) );
	vdp_aoi22 g5850 (.Z(w5834), .B2(w5904), .B1(w26), .A1(M5), .A2(w5841) );
	vdp_cnt_bit_load g5851 (.Q(w5934), .D(w5882), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w7), .CI(w5993), .L(w5880), .nL(w5927) );
	vdp_cnt_bit_load g5852 (.Q(w5879), .D(w5931), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w7), .CI(w5875), .L(w5880), .nL(w5927), .CO(w5993) );
	vdp_sr_bit g5853 (.Q(w5868), .D(w6391), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5854 (.SUM(w5886), .CO(w6635), .CI(1'b1), .A(HPOS[0]), .B(M5) );
	vdp_fa g5855 (.SUM(w5884), .CO(w6636), .CI(w6635), .A(HPOS[1]), .B(1'b0) );
	vdp_fa g5856 (.SUM(w5883), .CO(w6637), .CI(w6636), .A(HPOS[2]), .B(1'b1) );
	vdp_fa g5857 (.SUM(w5889), .CO(w6638), .CI(w6637), .A(HPOS[3]), .B(M5) );
	vdp_fa g5858 (.SUM(w5903), .CO(w6639), .CI(w6638), .A(HPOS[4]), .B(w5942) );
	vdp_fa g5859 (.SUM(w5892), .CO(w6640), .CI(w6639), .A(HPOS[5]), .B(1'b1) );
	vdp_fa g5860 (.SUM(w5893), .CO(w6641), .CI(w6640), .A(HPOS[6]), .B(1'b1) );
	vdp_fa g5861 (.SUM(w5894), .CO(w6642), .CI(w6641), .A(HPOS[7]), .B(1'b1) );
	vdp_fa g5862 (.SUM(w5895), .CI(w6642), .A(HPOS[8]), .B(1'b1) );
	vdp_not g5863 (.nZ(w5942), .A(M5) );
	vdp_aoi33 g5864 (.Z(w6391), .B2(w6653), .B1(w5897), .A1(H40), .A2(w5897), .A3(w5896), .B3(w6653) );
	vdp_not g5865 (.nZ(w6653), .A(H40) );
	vdp_or g5866 (.Z(w5896), .B(w5901), .A(w5902) );
	vdp_and g5867 (.Z(w5877), .B(w5875), .A(w5876) );
	vdp_sr_bit g5868 (.Q(w5875), .D(w6427), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5869 (.Q(w6427), .D(w5615), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5870 (.nQ(w5924), .D(w5466), .nC(nDCLK2), .C(DCLK2) );
	vdp_slatch g5871 (.Q(w5923), .D(w5910), .nC(w5863), .C(w5914) );
	vdp_slatch g5872 (.Q(w5862), .D(w5923), .nC(w5859), .C(w5916) );
	vdp_slatch g5873 (.Q(w5917), .D(w5908), .nC(w5863), .C(w5914) );
	vdp_slatch g5874 (.Q(w5860), .D(w5917), .nC(w5859), .C(w5916) );
	vdp_slatch g5875 (.Q(w5918), .D(w5909), .nC(w5863), .C(w5914) );
	vdp_slatch g5876 (.Q(w5861), .D(w5918), .nC(w5859), .C(w5916) );
	vdp_slatch g5877 (.Q(w6430), .D(w5620), .nC(w5863), .C(w5914) );
	vdp_sr_bit g5878 (.Q(w5865), .D(w6430), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_and g5879 (.Z(w5907), .B(DCLK2), .A(w5466) );
	vdp_comp_str g5880 (.nZ(w5859), .A(w5907), .Z(w5916) );
	vdp_comp_str g5881 (.nZ(w5863), .A(w5878), .Z(w5914) );
	vdp_not g5882 (.nZ(w5905), .A(w5924) );
	vdp_comp_we g5883 (.nZ(w5927), .A(w5877), .Z(w5880) );
	vdp_and3 g5884 (.Z(w5878), .B(HCLK1), .A(w5876), .C(w5875) );
	vdp_nand g5885 (.Z(w5931), .B(w5912), .A(M5) );
	vdp_nand g5886 (.Z(w5882), .B(w5911), .A(M5) );
	vdp_nor g5887 (.Z(w5876), .B(w5934), .A(w5879) );
	vdp_fa g5888 (.SUM(w5897), .CI(w5952), .A(w5951), .B(w5963) );
	vdp_aon22 g5889 (.Z(w5951), .B2(w5955), .B1(w5950), .A1(w5986), .A2(w5920) );
	vdp_sr_bit g5890 (.Q(w5950), .D(w5897), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5891 (.Q(w5986), .D(w5987), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5892 (.SUM(w5987), .CI(w5948), .A(w5949), .B(w5982) );
	vdp_aon22 g5893 (.Z(w5949), .B2(w5960), .B1(w5985), .A1(1'b0), .A2(w5913) );
	vdp_fa g5894 (.SUM(w5902), .CO(w5952), .CI(w5947), .A(w5946), .B(w5963) );
	vdp_aon22 g5895 (.Z(w5946), .B2(w5955), .B1(w5945), .A1(w5983), .A2(w5920) );
	vdp_sr_bit g5896 (.Q(w5945), .D(w5902), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5897 (.Q(w5983), .D(w5989), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5898 (.SUM(w5989), .CO(w5948), .CI(w5944), .A(w5943), .B(w5982) );
	vdp_aon22 g5899 (.Z(w5943), .B2(w5960), .B1(w5980), .A1(w5981), .A2(w5913) );
	vdp_fa g5900 (.SUM(w5901), .CO(w5947), .CI(w5941), .A(w5940), .B(w5963) );
	vdp_aon22 g5901 (.Z(w5940), .B2(w5955), .B1(w5939), .A1(w5979), .A2(w5920) );
	vdp_fa g5902 (.SUM(w5990), .CO(w5944), .CI(w5938), .A(w5937), .B(w5966) );
	vdp_aon22 g5903 (.Z(w5937), .B2(w5960), .B1(w5977), .A1(w5978), .A2(w5913) );
	vdp_sr_bit g5904 (.Q(w5939), .D(w5901), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5905 (.Q(w5979), .D(w5990), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5906 (.SUM(w5900), .CO(w5941), .CI(w5953), .A(w5936), .B(w5963) );
	vdp_aon22 g5907 (.Z(w5936), .B2(w5955), .B1(w5935), .A1(w5976), .A2(w5920) );
	vdp_sr_bit g5908 (.Q(w5935), .D(w5900), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5909 (.Q(w5976), .D(w5975), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5910 (.SUM(w5975), .CO(w5938), .CI(w5932), .A(w5933), .B(w5966) );
	vdp_aon22 g5911 (.Z(w5933), .B2(w5960), .B1(w6650), .A1(w5974), .A2(w5913) );
	vdp_fa g5912 (.SUM(w5899), .CO(w5953), .CI(w5929), .A(w5930), .B(w5963) );
	vdp_aon22 g5913 (.Z(w5930), .B2(w5955), .B1(w5928), .A1(w5973), .A2(w5920) );
	vdp_sr_bit g5914 (.Q(w5928), .D(w5899), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5915 (.Q(w5973), .D(w6643), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5916 (.SUM(w6643), .CO(w5932), .CI(w5926), .A(w5925), .B(w5972) );
	vdp_aon22 g5917 (.Z(w5925), .B2(w5960), .B1(w5991), .A1(w5971), .A2(w5913) );
	vdp_fa g5918 (.SUM(w5898), .CO(w5929), .CI(w5922), .A(w5921), .B(w5963) );
	vdp_aon22 g5919 (.Z(w5921), .B2(w5955), .B1(w5919), .A1(w5970), .A2(w5920) );
	vdp_sr_bit g5920 (.Q(w5919), .D(w5898), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5921 (.Q(w5970), .D(w5969), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5922 (.SUM(w5969), .CO(w5926), .CI(w5620), .A(w5915), .B(w5965) );
	vdp_aon22 g5923 (.Z(w5915), .B2(w5960), .B1(w5967), .A1(w5968), .A2(w5913) );
	vdp_aon22 g5924 (.Z(w5571), .B2(w5960), .B1(w5964), .A1(w5988), .A2(w5913) );
	vdp_aon22 g5925 (.Z(w5551), .B2(w5960), .B1(w5959), .A1(w5962), .A2(w5913) );
	vdp_aon22 g5926 (.Z(w5559), .B2(w5960), .B1(w5958), .A1(w5961), .A2(w5913) );
	vdp_and g5927 (.Z(w5922), .B(w5957), .A(w6649) );
	vdp_comp_we g5928 (.nZ(w5913), .A(M5), .Z(w5960) );
	vdp_comp_we g5929 (.nZ(w5955), .A(w6648), .Z(w5920) );
	vdp_sr_bit g5930 (.Q(w6648), .D(w5878), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5931 (.Q(w5956), .D(w5924), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5932 (.Q(w6003), .D(w6006), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5933 (.Q(w6006), .D(w6007), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5934 (.Q(w6007), .D(w6011), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5935 (.Q(w6011), .D(w6012), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5936 (.Q(w6012), .D(w6013), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5937 (.nQ(w6013), .D(w6016), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5938 (.nZ(w5964), .A(w6003) );
	vdp_sr_bit g5939 (.Q(w6017), .D(w6018), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5940 (.Q(w6018), .D(w6022), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5941 (.Q(w6022), .D(w6023), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5942 (.Q(w6023), .D(w6025), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5943 (.Q(w6025), .D(w6028), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5944 (.nQ(w6028), .D(w6027), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5945 (.nZ(w5967), .A(w6017) );
	vdp_sr_bit g5946 (.Q(w6029), .D(w6431), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5947 (.Q(w6431), .D(w6032), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5948 (.Q(w6032), .D(w6034), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5949 (.Q(w6034), .D(w6035), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5950 (.Q(w6035), .D(w6036), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5951 (.nQ(w6036), .D(w6040), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5952 (.nZ(w5991), .A(w6029) );
	vdp_sr_bit g5953 (.Q(w6041), .D(w6044), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5954 (.Q(w6044), .D(w6048), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5955 (.Q(w6048), .D(w6047), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5956 (.Q(w6047), .D(w6049), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5957 (.Q(w6049), .D(w6052), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5958 (.nQ(w6052), .D(w6053), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5959 (.nZ(w6650), .A(w6041) );
	vdp_sr_bit g5960 (.Q(w6056), .D(w6059), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5961 (.Q(w6059), .D(w6060), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5962 (.Q(w6060), .D(w6061), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5963 (.Q(w6061), .D(w6085), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5964 (.Q(w6085), .D(w6086), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5965 (.nQ(w6086), .D(w6066), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5966 (.nZ(w5977), .A(w6056) );
	vdp_sr_bit g5967 (.Q(w6087), .D(w6081), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5968 (.Q(w6081), .D(w6080), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5969 (.Q(w6080), .D(w6078), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5970 (.Q(w6078), .D(w6077), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5971 (.Q(w6077), .D(w6075), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5972 (.nQ(w6075), .D(w6065), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5973 (.nZ(w5980), .A(w6087) );
	vdp_sr_bit g5974 (.Q(w6651), .D(w6071), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5975 (.Q(w6071), .D(w6072), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5976 (.Q(w6072), .D(w6068), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5977 (.Q(w6068), .D(w6067), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5978 (.Q(w6067), .D(w6063), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5979 (.nQ(w6063), .D(w6064), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5980 (.nZ(w5985), .A(w6651) );
	vdp_and g5981 (.Z(w5963), .B(w5957), .A(w5865) );
	vdp_and g5982 (.Z(w5999), .B(w5620), .A(w5912) );
	vdp_and g5983 (.Z(w6000), .B(w5620), .A(w5911) );
	vdp_or g5984 (.Z(w5965), .B(w5999), .A(w5966) );
	vdp_and g5985 (.B(w6002), .A(M5), .Z(w5620) );
	vdp_or g5986 (.Z(w5972), .B(w6000), .A(w5966) );
	vdp_and g5987 (.Z(w5966), .B(w23), .A(w6660) );
	vdp_or g5988 (.Z(w5982), .B(w5966), .A(M5) );
	vdp_not g5989 (.nZ(w6660), .A(M5) );
	vdp_not g5990 (.nZ(w6649), .A(w5865) );
	vdp_nor g5991 (.Z(w5957), .B(w6648), .A(w5956) );
	vdp_sr_bit g5992 (.Q(w6015), .D(w6019), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5993 (.Q(w6019), .D(w6020), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5994 (.Q(w6020), .D(w6021), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5995 (.Q(w6021), .D(w6024), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5996 (.Q(w6024), .D(w6652), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5997 (.nQ(w6652), .D(w6094), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5998 (.nZ(w5909), .A(w6015) );
	vdp_sr_bit g5999 (.Q(w6004), .D(w6005), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6000 (.Q(w6005), .D(w6008), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6001 (.Q(w6008), .D(w6009), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6002 (.Q(w6009), .D(w6010), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6003 (.Q(w6010), .D(w6014), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6004 (.nQ(w6014), .D(w6093), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6005 (.nZ(w5910), .A(w6004) );
	vdp_sr_bit g6006 (.Q(w5994), .D(w5995), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6007 (.Q(w5995), .D(w5996), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6008 (.Q(w5996), .D(w5998), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6009 (.Q(w5998), .D(w5997), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6010 (.Q(w5997), .D(w6001), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6011 (.nQ(w6001), .D(w6092), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6012 (.nZ(w6002), .A(w5994) );
	vdp_sr_bit g6013 (.Q(w6026), .D(w6030), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6014 (.Q(w6030), .D(w6031), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6015 (.Q(w6031), .D(w6033), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6016 (.Q(w6033), .D(w6037), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6017 (.Q(w6037), .D(w6038), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6018 (.nQ(w6038), .D(w6099), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6019 (.nZ(w5908), .A(w6026) );
	vdp_sr_bit g6020 (.Q(w6039), .D(w6042), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6021 (.Q(w6042), .D(w6043), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6022 (.Q(w6043), .D(w6045), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6023 (.Q(w6045), .D(w6046), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6024 (.Q(w6046), .D(w6050), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6025 (.nQ(w6050), .D(w6095), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6026 (.nZ(w5912), .A(w6039) );
	vdp_sr_bit g6027 (.Q(w6051), .D(w6054), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6028 (.Q(w6054), .D(w6055), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6029 (.Q(w6055), .D(w6057), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6030 (.Q(w6057), .D(w6058), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6031 (.Q(w6058), .D(w6062), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6032 (.nQ(w6062), .D(w6096), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6033 (.nZ(w5911), .A(w6051) );
	vdp_sr_bit g6034 (.Q(w6083), .D(w6084), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6035 (.Q(w6084), .D(w6088), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6036 (.Q(w6088), .D(w6089), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6037 (.Q(w6089), .D(w6082), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6038 (.Q(w6082), .D(w6079), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6039 (.nQ(w6079), .D(w6097), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6040 (.nZ(w5958), .A(w6083) );
	vdp_sr_bit g6041 (.Q(w6074), .D(w6076), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6042 (.Q(w6076), .D(w6073), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6043 (.Q(w6073), .D(w6070), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6044 (.Q(w6070), .D(w6069), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6045 (.Q(w6069), .D(w6090), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6046 (.nQ(w6090), .D(w6098), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6047 (.nZ(w5959), .A(w6074) );
	vdp_slatch g6048 (.D(w6124), .nC(w6162), .C(w6102), .nQ(w5961) );
	vdp_slatch g6049 (.D(S[1]), .nC(w6163), .C(w6106), .Q(w6123) );
	vdp_slatch g6050 (.D(S[1]), .nC(w6164), .C(w6105), .Q(w6122) );
	vdp_aoi22 g6051 (.Z(w6121), .B2(w6168), .B1(w6123), .A1(w6122), .A2(w6103) );
	vdp_slatch g6052 (.D(S[0]), .nC(w6163), .C(w6106), .Q(w6126) );
	vdp_slatch g6053 (.D(S[0]), .nC(w6164), .C(w6105), .Q(w6125) );
	vdp_aoi22 g6054 (.Z(w6124), .B2(w6168), .B1(w6126), .A1(w6125), .A2(w6103) );
	vdp_slatch g6055 (.D(w6121), .nC(w6162), .C(w6102), .nQ(w5962) );
	vdp_slatch g6056 (.D(S[2]), .nC(w6163), .C(w6106), .Q(w6120) );
	vdp_slatch g6057 (.D(S[2]), .nC(w6164), .C(w6105), .Q(w6119) );
	vdp_aoi22 g6058 (.Z(w6205), .B2(w6168), .B1(w6120), .A1(w6119), .A2(w6103) );
	vdp_slatch g6059 (.D(w6205), .nC(w6162), .C(w6102), .nQ(w5988) );
	vdp_slatch g6060 (.D(S[3]), .nC(w6163), .C(w6106), .Q(w6118) );
	vdp_slatch g6061 (.D(S[3]), .nC(w6164), .C(w6105), .Q(w6117) );
	vdp_aoi22 g6062 (.Z(w6116), .B2(w6168), .B1(w6118), .A1(w6117), .A2(w6103) );
	vdp_slatch g6063 (.D(w6116), .nC(w6162), .C(w6102), .nQ(w5968) );
	vdp_slatch g6064 (.D(S[4]), .nC(w6163), .C(w6106), .Q(w6115) );
	vdp_slatch g6065 (.D(S[4]), .nC(w6164), .C(w6105), .Q(w6114) );
	vdp_aoi22 g6066 (.Z(w6113), .B2(w6168), .B1(w6115), .A1(w6114), .A2(w6103) );
	vdp_slatch g6067 (.D(w6113), .nC(w6162), .C(w6102), .nQ(w5971) );
	vdp_slatch g6068 (.D(S[5]), .nC(w6163), .C(w6106), .Q(w6112) );
	vdp_slatch g6069 (.D(S[5]), .nC(w6164), .C(w6105), .Q(w6111) );
	vdp_aoi22 g6070 (.Z(w6110), .B2(w6168), .B1(w6112), .A1(w6111), .A2(w6103) );
	vdp_slatch g6071 (.D(w6110), .nC(w6162), .C(w6102), .nQ(w5974) );
	vdp_slatch g6072 (.D(S[6]), .nC(w6163), .C(w6106), .Q(w6109) );
	vdp_slatch g6073 (.D(S[6]), .nC(w6164), .C(w6105), .Q(w6107) );
	vdp_aoi22 g6074 (.Z(w6108), .B2(w6168), .B1(w6109), .A1(w6107), .A2(w6103) );
	vdp_slatch g6075 (.D(w6108), .nC(w6162), .C(w6102), .nQ(w5978) );
	vdp_slatch g6076 (.D(S[7]), .nC(w6163), .C(w6106), .Q(w6104) );
	vdp_slatch g6077 (.D(S[7]), .nC(w6164), .C(w6105), .Q(w6100) );
	vdp_aoi22 g6078 (.Z(w6101), .B2(w6168), .B1(w6104), .A1(w6100), .A2(w6103) );
	vdp_slatch g6079 (.D(w6101), .nC(w6162), .C(w6102), .nQ(w5981) );
	vdp_comp_str g6080 (.nZ(w6162), .A(w5615), .Z(w6102) );
	vdp_comp_str g6081 (.nZ(w6163), .A(w4958), .Z(w6106) );
	vdp_comp_str g6082 (.nZ(w6164), .A(w4962), .Z(w6105) );
	vdp_comp_we g6083 (.nZ(w6168), .A(w6161), .Z(w6103) );
	vdp_sr_bit g6084 (.Q(w6159), .D(w6155), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6085 (.Z(w6155), .B(w6160), .A(w6127) );
	vdp_fa g6086 (.SUM(w6160), .CI(w6129), .A(w6159), .B(1'b0) );
	vdp_sr_bit g6087 (.Q(w6194), .D(w6150), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6088 (.Z(w6150), .B(w6156), .A(w6127) );
	vdp_fa g6089 (.SUM(w6156), .CO(w6129), .CI(w6130), .A(w6194), .B(1'b0) );
	vdp_sr_bit g6090 (.Q(w6151), .D(w6174), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6091 (.Z(w6174), .B(w6152), .A(w6127) );
	vdp_fa g6092 (.SUM(w6152), .CO(w6130), .CI(w6132), .A(w6151), .B(w6131) );
	vdp_sr_bit g6093 (.Q(w6147), .D(w6146), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6094 (.Z(w6146), .B(w6148), .A(w6127) );
	vdp_fa g6095 (.SUM(w6148), .CO(w6132), .CI(w6134), .A(w6147), .B(w6133) );
	vdp_sr_bit g6096 (.Q(w6137), .D(w6657), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6097 (.Q(w6657), .D(w22), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6098 (.nQ(w6135), .D(w6137), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g6099 (.nQ(w6127), .D(w6136), .nC(nHCLK1), .C(HCLK1) );
	vdp_and g6100 (.Z(w6131), .B(w6134), .A(w6143) );
	vdp_and g6101 (.Z(w6133), .B(w6134), .A(w6142) );
	vdp_and g6102 (.Z(w4584), .B(w6657), .A(w6219) );
	vdp_or g6103 (.Z(w6136), .B(w6140), .A(w6206) );
	vdp_not g6104 (.nZ(w6139), .A(M5) );
	vdp_not g6105 (.nZ(w6134), .A(w6135) );
	vdp_fa g6106 (.SUM(w6179), .CO(w6182), .CI(w6180), .A(w6233), .B(w6153) );
	vdp_aoi22 g6107 (.Z(w6245), .B2(w6165), .B1(w6181), .A1(w6179), .A2(w6229) );
	vdp_notif0 g6108 (.A(w6245), .nZ(VRAMA[9]), .nE(w6222) );
	vdp_fa g6109 (.SUM(w6170), .CO(w6180), .CI(w6176), .A(w6232), .B(w6157) );
	vdp_aoi22 g6110 (.Z(w6178), .B2(w6165), .B1(w6179), .A1(w6170), .A2(w6229) );
	vdp_notif0 g6111 (.A(w6178), .nZ(VRAMA[8]), .nE(w6222) );
	vdp_fa g6112 (.SUM(w6166), .CO(w6176), .CI(w6169), .A(w6231), .B(w6149) );
	vdp_aoi22 g6113 (.Z(w6177), .B2(w6165), .B1(w6170), .A1(w6166), .A2(w6229) );
	vdp_notif0 g6114 (.A(w6177), .nZ(VRAMA[7]), .nE(w6222) );
	vdp_fa g6115 (.SUM(w6172), .CO(w6169), .CI(1'b0), .A(w6230), .B(w6145) );
	vdp_aoi22 g6116 (.Z(w6167), .B2(w6165), .B1(w6166), .A1(w6172), .A2(w6229) );
	vdp_notif0 g6117 (.A(w6167), .nZ(VRAMA[6]), .nE(w6222) );
	vdp_not g6118 (.nZ(w6222), .A(w6236) );
	vdp_ha g6119 (.SUM(w6181), .B(w6234), .A(w6182), .CO(w6183) );
	vdp_aoi22 g6120 (.Z(w6185), .B2(w6165), .B1(w6184), .A1(w6181), .A2(w6229) );
	vdp_notif0 g6121 (.A(w6185), .nZ(VRAMA[10]), .nE(w6239) );
	vdp_ha g6122 (.SUM(w6184), .B(w6235), .A(w6183), .CO(w6186) );
	vdp_aoi22 g6123 (.Z(w6187), .B2(w6165), .B1(w6195), .A1(w6184), .A2(w6229) );
	vdp_notif0 g6124 (.A(w6187), .nZ(VRAMA[11]), .nE(w6239) );
	vdp_ha g6125 (.SUM(w6195), .B(w6238), .A(w6186), .CO(w6188) );
	vdp_aoi22 g6126 (.Z(w6190), .B2(w6165), .B1(w6189), .A1(w6195), .A2(w6229) );
	vdp_notif0 g6127 (.A(w6190), .nZ(VRAMA[12]), .nE(w6239) );
	vdp_ha g6128 (.SUM(w6189), .B(w6237), .A(w6188), .CO(w6192) );
	vdp_aoi22 g6129 (.Z(w6193), .B2(w6165), .B1(w6191), .A1(w6189), .A2(w6229) );
	vdp_notif0 g6130 (.A(w6193), .nZ(VRAMA[13]), .nE(w6239) );
	vdp_ha g6131 (.SUM(w6191), .B(w6241), .A(w6192), .CO(w6198) );
	vdp_aoi22 g6132 (.Z(w6196), .B2(w6165), .B1(w6197), .A1(w6191), .A2(w6229) );
	vdp_notif0 g6133 (.A(w6196), .nZ(VRAMA[14]), .nE(w6239) );
	vdp_ha g6134 (.SUM(w6197), .B(w6240), .A(w6198), .CO(w6199) );
	vdp_aoi22 g6135 (.Z(w6202), .B2(w6165), .B1(w6203), .A1(w6197), .A2(w6229) );
	vdp_notif0 g6136 (.A(w6202), .nZ(VRAMA[15]), .nE(w6239) );
	vdp_ha g6137 (.SUM(w6203), .B(w6243), .A(w6199) );
	vdp_aoi22 g6138 (.Z(w6201), .B2(w6165), .B1(w5232), .A1(w6203), .A2(w6229) );
	vdp_notif0 g6139 (.A(w6201), .nZ(VRAMA[16]), .nE(w6239) );
	vdp_not g6140 (.nZ(w6239), .A(w6236) );
	vdp_sr_bit g6141 (.Q(w6236), .D(w6390), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6142 (.nQ(w4507), .D(w6200), .nC(nHCLK2), .C(HCLK2) );
	vdp_and g6143 (.Z(w6390), .B(M5), .A(w22) );
	vdp_or9 g6144 (.Z(w6200), .B(w6098), .A(w6097), .C(w6016), .D(w6027), .F(w6053), .E(w6040), .G(w6066), .H(w6065), .I(w6064) );
	vdp_sr_bit g6145 (.Q(w4578), .D(w6536), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_sr_bit g6146 (.D(w6658), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_fa g6147 (.SUM(w6145), .CO(w6644), .CI(1'b0), .A(w6217), .B(w6146) );
	vdp_fa g6148 (.SUM(w6149), .CO(w6645), .CI(w6644), .A(w6218), .B(w6174) );
	vdp_fa g6149 (.SUM(w6157), .CO(w6646), .CI(w6645), .A(1'b0), .B(w6150) );
	vdp_fa g6150 (.SUM(w6153), .CI(w6646), .A(1'b0), .B(w6155) );
	vdp_notif0 g6151 (.A(1'b1), .nZ(VRAMA[0]), .nE(w6222) );
	vdp_notif0 g6152 (.A(1'b1), .nZ(VRAMA[1]), .nE(w6222) );
	vdp_not g6153 (.nZ(w6154), .A(w6223) );
	vdp_notif0 g6154 (.A(w6154), .nZ(VRAMA[2]), .nE(w6222) );
	vdp_not g6155 (.nZ(w6158), .A(w6225) );
	vdp_notif0 g6156 (.A(w6158), .nZ(VRAMA[3]), .nE(w6222) );
	vdp_not g6157 (.nZ(w6171), .A(w6224) );
	vdp_notif0 g6158 (.A(w6171), .nZ(VRAMA[4]), .nE(w6222) );
	vdp_notif0 g6159 (.A(w6173), .nZ(VRAMA[5]), .nE(w6222) );
	vdp_aoi22 g6160 (.Z(w6173), .B2(w6165), .B1(w6172), .A1(w6215), .A2(w6229) );
	vdp_comp_we g6161 (.nZ(w6165), .A(w1), .Z(w6229) );
	vdp_aon22 g6162 (.Z(w6217), .B2(w6141), .B1(w6215), .A1(w6213), .A2(w6216) );
	vdp_aon22 g6163 (.Z(w6218), .B2(w6141), .B1(w6213), .A1(w6212), .A2(w6216) );
	vdp_comp_we g6164 (.nZ(w6141), .A(w1), .Z(w6216) );
	vdp_or g6165 (.Z(w6658), .B(w6206), .A(w4584) );
	vdp_nor g6166 (.Z(w6536), .B(w6140), .A(w6139) );
	vdp_comp_str g6167 (.nZ(w6269), .A(w6226), .Z(w6242) );
	vdp_slatch g6168 (.D(w6272), .nC(w6269), .C(w6242), .Q(w6097) );
	vdp_aon22 g6169 (.Z(w6273), .B2(w6246), .B1(w6125), .A1(DB[0]), .A2(w6227) );
	vdp_slatch g6170 (.D(w6274), .nC(w6269), .C(w6242), .Q(w6098) );
	vdp_aon22 g6171 (.Z(w6275), .B2(w6246), .B1(w6122), .A1(DB[1]), .A2(w6227) );
	vdp_slatch g6172 (.D(w6276), .nC(w6269), .C(w6242), .Q(w6016) );
	vdp_aon22 g6173 (.Z(w6277), .B2(w6246), .B1(w6119), .A1(DB[2]), .A2(w6227) );
	vdp_slatch g6174 (.D(w6278), .nC(w6269), .C(w6242), .Q(w6027) );
	vdp_aon22 g6175 (.Z(w6279), .B2(w6246), .B1(w6117), .A1(DB[3]), .A2(w6227) );
	vdp_slatch g6176 (.D(w6280), .nC(w6269), .C(w6242), .Q(w6040) );
	vdp_aon22 g6177 (.Z(w6281), .B2(w6246), .B1(w6114), .A1(DB[4]), .A2(w6227) );
	vdp_slatch g6178 (.D(w6282), .nC(w6269), .C(w6242), .Q(w6053) );
	vdp_aon22 g6179 (.Z(w6283), .B2(w6246), .B1(w6111), .A1(DB[5]), .A2(w6227) );
	vdp_slatch g6180 (.D(w6284), .nC(w6269), .C(w6242), .Q(w6066) );
	vdp_aon22 g6181 (.Z(w6285), .B2(w6246), .B1(w6107), .A1(DB[6]), .A2(w6227) );
	vdp_slatch g6182 (.D(w6287), .nC(w6269), .C(w6242), .Q(w6065) );
	vdp_aon22 g6183 (.Z(w6288), .B2(w6246), .B1(w6100), .A1(DB[7]), .A2(w6227) );
	vdp_slatch g6184 (.D(w6286), .nC(w6269), .C(w6242), .Q(w6064) );
	vdp_aon22 g6185 (.Z(w6289), .B2(w6246), .B1(w5073), .A1(DB[8]), .A2(w6227) );
	vdp_slatch g6186 (.D(w6260), .nC(w6257), .C(w6228), .Q(w6232) );
	vdp_aon22 g6187 (.Z(w6296), .B2(w6246), .B1(w6120), .A1(DB[2]), .A2(w6227) );
	vdp_slatch g6188 (.D(w6259), .nC(w6257), .C(w6228), .Q(w6233) );
	vdp_aon22 g6189 (.Z(w6291), .B2(w6246), .B1(w6118), .A1(DB[3]), .A2(w6227) );
	vdp_slatch g6190 (.D(w6266), .nC(w6257), .C(w6228), .Q(w6234) );
	vdp_aon22 g6191 (.Z(w6292), .B2(w6246), .B1(w6115), .A1(DB[4]), .A2(w6227) );
	vdp_slatch g6192 (.D(w6265), .nC(w6257), .C(w6228), .Q(w6235) );
	vdp_aon22 g6193 (.Z(w6295), .B2(w6246), .B1(w6112), .A1(DB[5]), .A2(w6227) );
	vdp_slatch g6194 (.D(w6263), .nC(w6257), .C(w6228), .Q(w6238) );
	vdp_aon22 g6195 (.Z(w6297), .B2(w6246), .B1(w6109), .A1(DB[6]), .A2(w6227) );
	vdp_slatch g6196 (.D(w6264), .nC(w6257), .C(w6228), .Q(w6237) );
	vdp_aon22 g6197 (.Z(w6298), .B2(w6246), .B1(w6104), .A1(DB[7]), .A2(w6227) );
	vdp_slatch g6198 (.D(w6262), .nC(w6257), .C(w6228), .Q(w6241) );
	vdp_aon22 g6199 (.Z(w6299), .B2(w6246), .B1(w5013), .A1(DB[8]), .A2(w6227) );
	vdp_slatch g6200 (.D(w6255), .nC(w6257), .C(w6228), .Q(w6240) );
	vdp_aon22 g6201 (.Z(w6254), .B2(w6246), .B1(w5074), .A1(DB[9]), .A2(w6227) );
	vdp_slatch g6202 (.D(w6270), .nC(w6257), .C(w6228), .Q(w6243) );
	vdp_aon22 g6203 (.Z(w6271), .B2(w6246), .B1(w5082), .A1(DB[10]), .A2(w6227) );
	vdp_slatch g6204 (.D(w6258), .nC(w6257), .C(w6228), .Q(w6230) );
	vdp_aon22 g6205 (.Z(w6293), .B2(w6246), .B1(w6126), .A1(DB[0]), .A2(w6227) );
	vdp_slatch g6206 (.D(w6301), .nC(w6257), .C(w6228), .Q(w6231) );
	vdp_aon22 g6207 (.Z(w6294), .B2(w6246), .B1(w6123), .A1(DB[1]), .A2(w6227) );
	vdp_comp_str g6208 (.nZ(w6257), .A(w6226), .Z(w6228) );
	vdp_not g6209 (.nZ(w6226), .A(w6385) );
	vdp_oai21 g6210 (.Z(w6385), .B(HCLK1), .A1(w6140), .A2(w117) );
	vdp_sr_bit g6211 (.Q(w6386), .D(w6388), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6212 (.Q(w5615), .D(w6387), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6213 (.Q(w6161), .D(w6389), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6214 (.Q(w6290), .D(w5575), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g6215 (.Q(w6209), .D(w6214), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w6206), .CI(w22), .L(w6211), .nL(w6249), .CO(w6250) );
	vdp_cnt_bit_load g6216 (.Q(w6248), .D(w6210), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w6206), .CI(w6250), .L(w6211), .nL(w6249) );
	vdp_comp_we g6217 (.nZ(w6249), .A(w6140), .Z(w6211) );
	vdp_not g6218 (.nZ(w6214), .A(w6251) );
	vdp_not g6219 (.nZ(w6210), .A(w6247) );
	vdp_not g6220 (.nZ(w6207), .A(w120) );
	vdp_nand g6221 (.Z(w6302), .B(w120), .A(w4578) );
	vdp_nand g6222 (.Z(w6208), .B(w6207), .A(w4578) );
	vdp_not g6223 (.nZ(w6246), .A(w6208) );
	vdp_nor g6224 (.Z(w6219), .B(w6248), .A(w6209) );
	vdp_and g6225 (.Z(w6140), .B(w6219), .A(w22) );
	vdp_rs_ff g6226 (.Q(w6388), .R(w6220), .S(w6206) );
	vdp_and3 g6227 (.Z(w6387), .B(w5575), .A(w4585), .C(w6386) );
	vdp_cnt_bit g6228 (.Q(w6389), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w7), .CI(w6290) );
	vdp_not g6229 (.nZ(w6227), .A(w6302) );
	vdp_not g6230 (.nZ(w6253), .A(w4542) );
	vdp_not g6231 (.nZ(w6256), .A(w4543) );
	vdp_comp_str g6232 (.nZ(w6252), .A(w6226), .Z(w6304) );
	vdp_not g6233 (.nZ(w6312), .A(w117) );
	vdp_aon22 g6234 (.Z(w6314), .B2(w6246), .B1(w5134), .A1(DB[0]), .A2(w6227) );
	vdp_slatch g6235 (.D(w6303), .nC(w6252), .C(w6304), .Q(w6092) );
	vdp_bufif0 g6236 (.A(w6311), .Z(DB[0]), .nE(w6312) );
	vdp_aon222 g6237 (.Z(w6311), .B2(w4544), .B1(w6097), .A1(w6092), .A2(w6253), .C1(w6230), .C2(w6256) );
	vdp_aon22 g6238 (.Z(w6317), .B2(w6246), .B1(w5213), .A1(DB[1]), .A2(w6227) );
	vdp_slatch g6239 (.D(w6313), .nC(w6252), .C(w6304), .Q(w6093) );
	vdp_bufif0 g6240 (.A(w6315), .Z(DB[1]), .nE(w6312) );
	vdp_aon222 g6241 (.Z(w6315), .B2(w4544), .B1(w6098), .A1(w6093), .A2(w6253), .C1(w6231), .C2(w6256) );
	vdp_aon22 g6242 (.Z(w6319), .B2(w6246), .B1(w5233), .A1(DB[2]), .A2(w6227) );
	vdp_slatch g6243 (.D(w6316), .nC(w6252), .C(w6304), .Q(w6094) );
	vdp_bufif0 g6244 (.A(w6318), .Z(DB[2]), .nE(w6312) );
	vdp_aon222 g6245 (.Z(w6318), .B2(w4544), .B1(w6016), .A1(w6094), .A2(w6253), .C1(w6232), .C2(w6256) );
	vdp_aon22 g6246 (.Z(w6328), .B2(w6246), .B1(w5198), .A1(DB[3]), .A2(w6227) );
	vdp_slatch g6247 (.D(w6320), .nC(w6252), .C(w6304), .Q(w6099) );
	vdp_bufif0 g6248 (.A(w6327), .Z(DB[3]), .nE(w6312) );
	vdp_aon222 g6249 (.Z(w6327), .B2(w4544), .B1(w6027), .A1(w6099), .A2(w6253), .C1(w6233), .C2(w6256) );
	vdp_aon22 g6250 (.Z(w6325), .B2(w6246), .B1(w4523), .A1(DB[4]), .A2(w6227) );
	vdp_slatch g6251 (.D(w6251), .nC(w6252), .C(w6304), .Q(w6095) );
	vdp_bufif0 g6252 (.A(w6326), .Z(DB[4]), .nE(w6312) );
	vdp_aon222 g6253 (.Z(w6326), .B2(w4544), .B1(w6040), .A1(w6095), .A2(w6253), .C1(w6234), .C2(w6256) );
	vdp_aon22 g6254 (.Z(w6323), .B2(w6246), .B1(w4568), .A1(DB[5]), .A2(w6227) );
	vdp_slatch g6255 (.D(w6247), .nC(w6252), .C(w6304), .Q(w6096) );
	vdp_bufif0 g6256 (.A(w6324), .Z(DB[5]), .nE(w6312) );
	vdp_aon222 g6257 (.Z(w6324), .B2(w4544), .B1(w6053), .A1(w6096), .A2(w6253), .C1(w6235), .C2(w6256) );
	vdp_aon22 g6258 (.Z(w6321), .B2(w6246), .B1(w4524), .A1(DB[6]), .A2(w6227) );
	vdp_slatch g6259 (.D(w6322), .nC(w6252), .C(w6304), .Q(w6142) );
	vdp_bufif0 g6260 (.A(w6344), .Z(DB[6]), .nE(w6312) );
	vdp_aon222 g6261 (.Z(w6344), .B2(w4544), .B1(w6066), .A1(w6142), .A2(w6253), .C1(w6238), .C2(w6256) );
	vdp_aon22 g6262 (.Z(w6340), .B2(w6246), .B1(w4520), .A1(DB[7]), .A2(w6227) );
	vdp_slatch g6263 (.D(w6341), .nC(w6261), .C(w6342), .Q(w6143) );
	vdp_bufif0 g6264 (.A(w6343), .Z(DB[7]), .nE(w6312) );
	vdp_aon222 g6265 (.Z(w6343), .B2(w4544), .B1(w6065), .A1(w6143), .A2(w6253), .C1(w6237), .C2(w6256) );
	vdp_aon22 g6266 (.Z(w6338), .B2(w6246), .B1(w6305), .A1(DB[8]), .A2(w6227) );
	vdp_slatch g6267 (.D(w6339), .nC(w6261), .C(w6342), .Q(w6223) );
	vdp_bufif0 g6268 (.A(w6659), .Z(DB[8]), .nE(w6312) );
	vdp_aon222 g6269 (.Z(w6659), .B2(w4544), .B1(w6064), .A1(w6223), .A2(w6253), .C1(w6241), .C2(w6256) );
	vdp_aon22 g6270 (.Z(w6336), .B2(w6246), .B1(w6310), .A1(DB[9]), .A2(w6227) );
	vdp_slatch g6271 (.D(w6337), .nC(w6261), .C(w6342), .Q(w6225) );
	vdp_bufif0 g6272 (.A(w6345), .Z(DB[9]), .nE(w6312) );
	vdp_aon222 g6273 (.Z(w6345), .B2(w4544), .B1(1'b0), .A1(w6225), .A2(w6253), .C1(w6240), .C2(w6256) );
	vdp_aon22 g6274 (.Z(w6334), .B2(w6246), .B1(w6309), .A1(DB[10]), .A2(w6227) );
	vdp_slatch g6275 (.D(w6335), .nC(w6261), .C(w6342), .Q(w6224) );
	vdp_bufif0 g6276 (.A(w6346), .Z(DB[10]), .nE(w6312) );
	vdp_aon222 g6277 (.Z(w6346), .B2(w4544), .B1(1'b0), .A1(w6224), .A2(w6253), .C1(w6243), .C2(w6256) );
	vdp_aon22 g6278 (.Z(w6332), .B2(w6246), .B1(w6308), .A1(DB[11]), .A2(w6227) );
	vdp_slatch g6279 (.D(w6333), .nC(w6261), .C(w6342), .Q(w6215) );
	vdp_bufif0 g6280 (.A(w6215), .Z(DB[11]), .nE(w6312) );
	vdp_aon22 g6281 (.Z(w6331), .B2(w6246), .B1(w6307), .A1(DB[12]), .A2(w6227) );
	vdp_slatch g6282 (.D(w6347), .nC(w6261), .C(w6342), .Q(w6213) );
	vdp_bufif0 g6283 (.A(w6213), .Z(DB[12]), .nE(w6312) );
	vdp_aon22 g6284 (.Z(w6329), .B2(w6246), .B1(w6306), .A1(DB[13]), .A2(w6227) );
	vdp_slatch g6285 (.D(w6330), .nC(w6261), .C(w6342), .Q(w6212) );
	vdp_bufif0 g6286 (.A(w6212), .Z(DB[13]), .nE(w6312) );
	vdp_comp_str g6287 (.nZ(w6261), .A(w6226), .Z(w6342) );
	vdp_sr_bit g6288 (.Q(w4687), .D(w126), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6289 (.Q(w4688), .D(VRAMA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6290 (.Q(w6356), .D(w6349), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6291 (.Q(w4680), .D(VRAMA[3]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6292 (.Q(w4682), .D(VRAMA[4]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6293 (.Q(w4683), .D(VRAMA[5]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6294 (.Q(w4684), .D(VRAMA[6]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6295 (.Q(w4685), .D(VRAMA[7]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6296 (.Q(w4686), .D(VRAMA[8]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6297 (.Q(w4627), .D(w6353), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6298 (.Q(w4626), .D(w6354), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_and g6299 (.Z(w6353), .B(w129), .A(w6355) );
	vdp_and g6300 (.Z(w6354), .B(w128), .A(w6355) );
	vdp_sr_bit g6301 (.Q(w6369), .D(RD_DATA[0]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6302 (.Q(w6370), .D(RD_DATA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6303 (.Q(w6372), .D(w321), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6304 (.Q(w6371), .D(RD_DATA[2]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_V_PLA g6305 (.o[0](w1878), .o[1](w1879), .o[2](w1880), .o[3](w1881), .o[4](w1882), .o[5](w1883), .o[6](w1884), .o[7](w1885), .o[8](w1886), .o[9](w1887), .o[10](w1888), .o[11](w1889), .o[12](w1890), .o[13](w1891), .o[14](w1892), .o[15](w6777), .o[16](w6778), .o[17](w6779), .o[18](w1893), .o[19](w1894), .o[20](w1895), .o[21](w1896), .o[22](w6780), .o[23](w1897), .o[24](w1971), .o[25](w1898), .o[26](w1899), .o[27](w1972), .o[28](w1986), .o[29](w1985), .o[30](w2006), .o[31](w1915), .o[32](w1877), .o[33](w1876), .o[34](w1916), .o[35](w1900), .o[36](w1917), .o[37](w1918), .o[38](w1875), .o[39](w1874), .o[40](w1921), .o[41](w1919), .o[42](w1920), .o[43](w1872), .o[44](w1871), .o[45](w1870), .o[46](w1869), .o[47](w6666), .Vcnt[0](w1695), .Vcnt[1](w1837), .Vcnt[2](w1929), .Vcnt[3](w1822), .Vcnt[4](w1928), .Vcnt[5](w1776), .Vcnt[6](w1739), .Vcnt[7](w1811), .Vcnt[8](w1838), .ODD_EVEN(ODD_EVEN), .LS0(LS0), .PAL(PAL), .nPAL(w1830), .2(w1829), .3(w1818), .M5(M5) );
	vdp_not g6306 (.A(w588), .nZ(w6664) );
	vdp_not g6307 (.A(w961), .nZ(w6665) );
	vdp_not g6308 (.nZ(w2444), .A(w6664) );
	vdp_not g6309 (.nZ(w2445), .A(w6665) );
	vdp_cram g6310 (.q[8](w2743), .D[8](w2744), .q[7](w2845), .D[7](w2745), .q[6](w2742), .D[6](w2746), .q[5](w2748), .D[5](w2747), .q[4](w2741), .D[4](w2749), .q[3](w2750), .D[3](w2974), .q[2](w2740), .D[2](w2751), .q[1](w2739), .D[1](w2752), .q[0](w2737), .D[0](w2753), .A[0](w2772), .A[1](w2776), .CLK(HCLK1), .A[2](w2782), .A[3](w2792), .A[4](w2813), .A[5](w2812), .B(w2819), .A(w2818) );
	vdp_linebuf_ram g6311 (.q[0](w5315), .D[0](w5706), .q[1](w5304), .D[1](w5705), .q[2](w5292), .D[2](w5704), .q[3](w5281), .D[3](w5717), .q[4](w5716), .D[4](w5691), .q[5](w5685), .D[5](w5690), .q[6](w5696), .D[6](w5718), .q[7](w5314), .D[7](w5703), .q[8](w5305), .D[8](w5702), .q[9](w5291), .D[9](w5701), .q[10](w5282), .D[10](w5678), .q[11](w5679), .D[11](w5677), .q[12](w5697), .D[12](w5682), .q[13](w5698), .D[13](w5715), .q[14](w5313), .D[14](w5706), .q[15](w5306), .D[15](w5705), .q[16](w5290), .D[16](w5704), .q[17](w5283), .D[17](w5707), .q[18](w5680), .D[18](w5712), .q[19](w5684), .D[19](w5708), .q[20](w5710), .D[20](w5709), .q[21](w5312), .D[21](w5703), .q[22](w5307), .D[22](w5702), .q[23](w5289), .D[23](w5701), .q[24](w5284), .D[24](w5694), .q[25](w5681), .D[25](w5692), .q[26](w5683), .D[26](w5700), .q[27](w5711), .D[27](w5699), .CLK(w4505), .A[5](w4499), .A[4](w4500), .A[3](w4501), .A[2](w4502), .A[1](w4503), .A[0](w4504), .A(w5714), .B(w5676), .C(w5675), .D(w5674) );
	vdp_linebuf_ram g6312 (.q[0](w5350), .D[0](w5706), .q[1](w5321), .D[1](w5705), .q[2](w5296), .D[2](w5704), .q[3](w5279), .D[3](w5345), .q[4](w5320), .D[4](w5311), .q[5](w5319), .D[5](w5310), .q[6](w5693), .D[6](w5367), .q[7](w5318), .D[7](w5703), .q[8](w5301), .D[8](w5702), .q[9](w5295), .D[9](w5701), .q[10](w5358), .D[10](w5343), .q[11](w5299), .D[11](w5309), .q[12](w5300), .D[12](w5308), .q[13](w5689), .D[13](w5339), .q[14](w5317), .D[14](w5706), .q[15](w5302), .D[15](w5705), .q[16](w5294), .D[16](w5704), .q[17](w5364), .D[17](w5325), .q[18](w5297), .D[18](w5288), .q[19](w5298), .D[19](w5323), .q[20](w5688), .D[20](w5324), .q[21](w5316), .D[21](w5703), .q[22](w5303), .D[22](w5702), .q[23](w5293), .D[23](w5701), .q[24](w5359), .D[24](w6351), .q[25](w5687), .D[25](w5287), .q[26](w5686), .D[26](w5286), .q[27](w5695), .D[27](w5285), .A[0](w4504), .CLK(w4505), .A[5](w4499), .A[3](w4501), .A[4](w4500), .A[2](w4502), .A[1](w4503), .A(w5408), .B(w5392), .C(w5404), .D(w5394) );
	vdp_att_cashe_ram2 g6313 (.q[0](w4704), .D[0](FIFOo[0]), .q[1](w4703), .D[1](FIFOo[1]), .q[2](w4702), .D[2](FIFOo[2]), .q[3](w4701), .D[3](FIFOo[3]), .q[4](w4677), .D[4](FIFOo[4]), .q[5](w4676), .D[5](FIFOo[5]), .q[6](w4671), .D[6](FIFOo[6]), .q[7](w4847), .D[7](w6369), .q[8](w4885), .D[8](w6370), .q[9](w4870), .D[9](w6371), .q[10](w4867), .D[10](w6372), .CLK(HCLK1), .A[6](w6377), .A[5](w6378), .A[1](w6383), .A[0](w6382), .A[4](w6379), .A[3](w6380), .A[2](w6381), .A(w6374), .B(w4690) );
	vdp_att_cashe_ram1 g6314 (.q[0](w4736), .D[0](FIFOo[0]), .q[1](w4739), .D[1](FIFOo[1]), .q[2](w4732), .D[2](FIFOo[2]), .q[3](w4733), .D[3](FIFOo[3]), .q[4](w4715), .D[4](FIFOo[4]), .q[5](w4707), .D[5](FIFOo[5]), .q[6](w4708), .D[6](FIFOo[6]), .q[7](w4706), .D[7](FIFOo[7]), .q[8](w4705), .D[8](w6369), .q[9](w4700), .D[9](w6370), .CLK(HCLK1), .A[0](w6382), .A[1](w6383), .A[2](w6381), .A[3](w6380), .A[4](w6379), .A[5](w6378), .A[6](w6377), .A(w6376), .B(w6375) );
	vdp_att_temp_ram g6315 (.A[4](w4602), .A[0](w4606), .A[1](w4605), .A[2](w4604), .A[3](w4603), .q[0](w6258), .D[0](w6293), .q[1](w6301), .D[1](w6294), .q[2](w6260), .D[2](w6296), .q[3](w6259), .D[3](w6291), .q[4](w6266), .D[4](w6292), .q[5](w6265), .D[5](w6295), .q[6](w6263), .D[6](w6297), .q[7](w6264), .D[7](w6298), .q[8](w6262), .D[8](w6299), .q[9](w6255), .D[9](w6254), .q[10](w6270), .D[10](w6271), .q[11](w6272), .D[11](w6273), .q[12](w6274), .D[12](w6275), .q[13](w6276), .D[13](w6277), .q[14](w6278), .D[14](w6279), .q[15](w6280), .D[15](w6281), .q[16](w6282), .D[16](w6283), .q[17](w6284), .D[17](w6285), .q[18](w6287), .D[18](w6288), .q[19](w6286), .D[19](w6289), .q[20](w6303), .D[20](w6314), .q[21](w6313), .D[21](w6317), .q[22](w6316), .D[22](w6319), .q[23](w6320), .D[23](w6328), .q[24](w6251), .D[24](w6325), .q[25](w6247), .D[25](w6323), .q[26](w6322), .D[26](w6321), .q[26](w6341), .D[26](w6340), .q[27](w6339), .D[27](w6338), .q[28](w6337), .D[28](w6336), .q[29](w6335), .D[29](w6334), .q[30](w6333), .D[30](w6332), .q[31](w6347), .D[31](w6331), .q[32](w6330), .D[32](w6329), .CLK(HCLK1), .A(w4569), .B(w4570), .C(w4574) );
	vdp_vsram g6316 (.CLK(HCLK1), .D[10](w3992), .q[10](w3950), .D[9](w3996), .q[9](w3943), .D[8](w3994), .q[8](w3969), .D[7](w3993), .q[7](w3935), .D[6](w3981), .q[6](w3931), .D[5](w3979), .q[5](w3923), .D[4](w3986), .q[4](w3919), .D[3](w3988), .q[3](w3916), .D[2](w3991), .q[2](w3974), .D[1](w3949), .q[1](w3911), .D[0](w3967), .q[0](w3906), .A[1](w3723), .A[2](w3695), .A[3](w3694), .A[4](w3693), .A[5](w3692), .A[0](w3724), .A(w3691), .B(w3690) );
	vdp_not g6317 (.nZ(w1812), .A(w6666) );
	vdp_not g6318 (.nZ(PAL), .A(w6667) );
	vdp_H_PLA g6319 (.HPLA[0](w1931), .HPLA[1](w1912), .HPLA[2](w1904), .HPLA[3](w1740), .HPLA[4](w1902), .HPLA[5](w1905), .HPLA[7](w1741), .HPLA[8](w1742), .HPLA[9](w1862), .HPLA[6](w1743), .HPLA[10](w1865), .HPLA[11](w1908), .HPLA[16](w1866), .HPLA[15](w1910), .HPLA[14](w1909), .HPLA[13](w1913), .HPLA[12](w1914), .i0(w59), .HPLA[17](w1763), .HPLA[18](w1762), .HPLA[19](w1864), .HPLA[20](w1863), .HPLA[21](w1906), .HPLA[22](w1901), .Hcnt[0](w1932), .Hcnt[1](w1679), .Hcnt[2](w1684), .Hcnt[3](w1683), .Hcnt[4](w1728), .Hcnt[5](w1760), .Hcnt[6](w1907), .Hcnt[7](w1737), .Hcnt[8](w1765), .H40(H40), .M5(M5), .B(w1764), .C(w1663), .A(w1733), .HPLA[23](w1682), .HPLA[24](w1680), .HPLA[25](w1681), .HPLA[26](w1678), .HPLA[27](w1867), .HPLA[28](w1860), .HPLA[29](w1664), .HPLA[30](w1717), .HPLA[31](w1665), .HPLA[32](w1903), .HPLA[33](w1757), .3(w1911), .HPLA[35](w1793), .HPLA[36](w1755), .HPLA[34](w1933) );
	vdp_slatch g5073 (.D(S[4]), .nC(w5018), .C(w5019), .Q(w5212) );
endmodule // VDP

// Module Definitions [It is possible to wrap here on your primitives]

module vdp_slatch (  nQ, D, C, nC);

	output wire nQ;
	input wire D;
	input wire C;
	input wire nC;

endmodule // vdp_slatch

module vdp_sr_bit (  D, C2, C1, Q, nC2, nC1);

	input wire D;
	input wire C2;
	input wire C1;
	output wire Q;
	input wire nC2;
	input wire nC1;

endmodule // vdp_sr_bit

module vdp_notif0 (  A, nZ, nE);

	input wire A;
	output wire nZ;
	input wire nE;

endmodule // vdp_notif0

module vdp_aon22 (  Z, A1, A2, B1, B2);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire B1;
	input wire B2;

endmodule // vdp_aon22

module vdp_not (  A, nZ);

	input wire A;
	output wire nZ;

endmodule // vdp_not

module vdp_comp_str (  A, Z, nZ);

	input wire A;
	output wire Z;
	output wire nZ;

endmodule // vdp_comp_str

module vdp_comp_we (  A, Z, nZ);

	input wire A;
	output wire Z;
	output wire nZ;

endmodule // vdp_comp_we

module vdp_and (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_and

module vdp_nand (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_nand

module vdp_and3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_and3

module vdp_fa (  SUM, A, B, CO, CI);

	output wire SUM;
	input wire A;
	input wire B;
	output wire CO;
	input wire CI;

endmodule // vdp_fa

module vdp_comp_dff (  D, C2, C1, Q, nC2, nC1);

	input wire D;
	input wire C2;
	input wire C1;
	output wire Q;
	input wire nC2;
	input wire nC1;

endmodule // vdp_comp_dff

module vdp_or (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_or

module vdp_xor (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_xor

module vdp_aoi21 (  Z, B, A1, A2);

	output wire Z;
	input wire B;
	input wire A1;
	input wire A2;

endmodule // vdp_aoi21

module vdp_nor (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_nor

module vdp_and5 (  Z, A, B, C, D, E);

	output wire Z;
	input wire A;
	input wire B;
	input wire C;
	input wire D;
	input wire E;

endmodule // vdp_and5

module vdp_aon2222 (  C2, B2, A2, C1, B1, A1, Z, D2, D1);

	input wire C2;
	input wire B2;
	input wire A2;
	input wire C1;
	input wire B1;
	input wire A1;
	output wire Z;
	input wire D2;
	input wire D1;

endmodule // vdp_aon2222

module vdp_cnt_bit (  R, Q, C1, C2, nC1, nC2, CI);

	input wire R;
	output wire Q;
	input wire C1;
	input wire C2;
	input wire nC1;
	input wire nC2;
	input wire CI;

endmodule // vdp_cnt_bit

module vdp_oai21 (  A1, Z, A2, B);

	input wire A1;
	output wire Z;
	input wire A2;
	input wire B;

endmodule // vdp_oai21

module vdp_comb1 (  Z, A1, B, A2, C);

	output wire Z;
	input wire A1;
	input wire B;
	input wire A2;
	input wire C;

endmodule // vdp_comb1

module vdp_rs_ff (  Q, R, S);

	output wire Q;
	input wire R;
	input wire S;

endmodule // vdp_rs_ff

module vdp_and4 (  A, Z, B, C, D);

	input wire A;
	output wire Z;
	input wire B;
	input wire C;
	input wire D;

endmodule // vdp_and4

module vdp_or3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_or3

module vdp_bufif0 (  A, Z, nE);

	input wire A;
	output wire Z;
	input wire nE;

endmodule // vdp_bufif0

module vdp_aoi221 (  Z, A2, B1, B2, A1, C);

	output wire Z;
	input wire A2;
	input wire B1;
	input wire B2;
	input wire A1;
	input wire C;

endmodule // vdp_aoi221

module vdp_aon33 (  Z, A2, B1, B2, A1, A3, B3);

	output wire Z;
	input wire A2;
	input wire B1;
	input wire B2;
	input wire A1;
	input wire A3;
	input wire B3;

endmodule // vdp_aon33

module vdp_dlatch_inv (  D, C, Q, nC);

	input wire D;
	input wire C;
	output wire Q;
	input wire nC;

endmodule // vdp_dlatch_inv

module vdp_cnt_bit_load (  D, nL, L, R, Q, C1, C2, nC1, nC2, CI, CO);

	input wire D;
	input wire nL;
	input wire L;
	input wire R;
	output wire Q;
	input wire C1;
	input wire C2;
	input wire nC1;
	input wire nC2;
	input wire CI;
	output wire CO;

endmodule // vdp_cnt_bit_load

module vdp_nand3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_nand3

module vdp_nor3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_nor3

module vdp_dff (  Q, R, C, D);

	output wire Q;
	input wire R;
	input wire C;
	input wire D;

endmodule // vdp_dff

module vdp_ha (  SUM, A, B, CO);

	output wire SUM;
	input wire A;
	input wire B;
	output wire CO;

endmodule // vdp_ha

module vdp_slatch_r (  Q, D, R, C, nC);

	output wire Q;
	input wire D;
	input wire R;
	input wire C;
	input wire nC;

endmodule // vdp_slatch_r

module vdp_or5 (  C, A, B, Z, D, E);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;
	input wire E;

endmodule // vdp_or5

module vdp_2a3oi (  A1, B, Z, A2, C);

	input wire A1;
	input wire B;
	output wire Z;
	input wire A2;
	input wire C;

endmodule // vdp_2a3oi

module vdp_nor5 (  C, A, B, Z, D, E);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;
	input wire E;

endmodule // vdp_nor5

module vdp_or4 (  C, A, B, Z, D);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;

endmodule // vdp_or4

module vdp_aoi22 (  Z, A1, A2, B1, B2);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire B1;
	input wire B2;

endmodule // vdp_aoi22

module vdp_aon222 (  C2, B2, A2, C1, B1, A1, Z);

	input wire C2;
	input wire B2;
	input wire A2;
	input wire C1;
	input wire B1;
	input wire A1;
	output wire Z;

endmodule // vdp_aon222

module vdp_dlatch (  D, C, Q, nC);

	input wire D;
	input wire C;
	output wire Q;
	input wire nC;

endmodule // vdp_dlatch

module vdp_nor4 (  C, A, B, Z, D);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;

endmodule // vdp_nor4

module vdp_and6 (  C, A, B, Z, D, E, F);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;
	input wire E;
	input wire F;

endmodule // vdp_and6

module vdp_n_fet (  Z, A);

	output wire Z;
	input wire A;

endmodule // vdp_n_fet

module vdp_2A3OI (  Z, A1, A2, C, B);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire C;
	input wire B;

endmodule // vdp_2A3OI

module vdp_tff (  C2, C1, nC2, nC1, CI, R, A, Q);

	input wire C2;
	input wire C1;
	input wire nC2;
	input wire nC1;
	input wire CI;
	input wire R;
	input wire A;
	output wire Q;

endmodule // vdp_tff

module vdp_SDELAY8 (  Q, D, nC1, C1, nC2, C2, nC3, C3, nC4, C4, nC5, C5, nC6, C6, nC7, C7, nC8, C8, nC9, C9, nC10, C10, nC11, C11, nC12, C12, nC13, C13, nC14, C14, nC15, C15, nC16, C16);

	output wire Q;
	input wire D;
	input wire nC1;
	input wire C1;
	input wire nC2;
	input wire C2;
	input wire nC3;
	input wire C3;
	input wire nC4;
	input wire C4;
	input wire nC5;
	input wire C5;
	input wire nC6;
	input wire C6;
	input wire nC7;
	input wire C7;
	input wire nC8;
	input wire C8;
	input wire nC9;
	input wire C9;
	input wire nC10;
	input wire C10;
	input wire nC11;
	input wire C11;
	input wire nC12;
	input wire C12;
	input wire nC13;
	input wire C13;
	input wire nC14;
	input wire C14;
	input wire nC15;
	input wire C15;
	input wire nC16;
	input wire C16;

endmodule // vdp_SDELAY8

module vdp_SDELAY7 (  Q, D, C1, nC1, C2, nC2, nC3, C4, nC4, C5, nC5, C6, nC6, C7, nC7, C8, nC8, C9, nC9, C10, nC10, C11, nC11, C12, nC12, C13, nC13, C14, nC14, C3);

	output wire Q;
	input wire D;
	input wire C1;
	input wire nC1;
	input wire C2;
	input wire nC2;
	input wire nC3;
	input wire C4;
	input wire nC4;
	input wire C5;
	input wire nC5;
	input wire C6;
	input wire nC6;
	input wire C7;
	input wire nC7;
	input wire C8;
	input wire nC8;
	input wire C9;
	input wire nC9;
	input wire C10;
	input wire nC10;
	input wire C11;
	input wire nC11;
	input wire C12;
	input wire nC12;
	input wire C13;
	input wire nC13;
	input wire C14;
	input wire nC14;
	input wire C3;

endmodule // vdp_SDELAY7

module vdp_or8 (  Z, A, B, C, D, E, F, G, H);

	output wire Z;
	input wire A;
	input wire B;
	input wire C;
	input wire D;
	input wire E;
	input wire F;
	input wire G;
	input wire H;

endmodule // vdp_or8

module vdp_or7 (  Z, A, B, C, D, E, F, G);

	output wire Z;
	input wire A;
	input wire B;
	input wire C;
	input wire D;
	input wire E;
	input wire F;
	input wire G;

endmodule // vdp_or7

module vdp_clkgen (  PH, CLK1, nCLK1, CLK2, nCLK2);

	input wire PH;
	output wire CLK1;
	output wire nCLK1;
	output wire CLK2;
	output wire nCLK2;

endmodule // vdp_clkgen

module vdp_cgi2a (  Z, A, C, B);

	output wire Z;
	input wire A;
	input wire C;
	input wire B;

endmodule // vdp_cgi2a

module vdp_nand4 (  Z, A, B, D, C);

	output wire Z;
	input wire A;
	input wire B;
	input wire D;
	input wire C;

endmodule // vdp_nand4

module vdp_lfsr_bit (  Q, A, C2, C1, nC2, nC1, C, B);

	output wire Q;
	input wire A;
	input wire C2;
	input wire C1;
	input wire nC2;
	input wire nC1;
	input wire C;
	input wire B;

endmodule // vdp_lfsr_bit

module vdp_aoi222 (  Z, A1, B1, B2, A2, C1, C2);

	output wire Z;
	input wire A1;
	input wire B1;
	input wire B2;
	input wire A2;
	input wire C1;
	input wire C2;

endmodule // vdp_aoi222

module vdp_aon333 (  Z, A1, A2, A3, B1, B2, B3, C1, C2, C3);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire A3;
	input wire B1;
	input wire B2;
	input wire B3;
	input wire C1;
	input wire C2;
	input wire C3;

endmodule // vdp_aon333

module vdp_aoi33 (  Z, A1, A2, A3, B1, B2, B3);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire A3;
	input wire B1;
	input wire B2;
	input wire B3;

endmodule // vdp_aoi33

module vdp_comp_strong (  nZ, Z, A);

	output wire nZ;
	output wire Z;
	input wire A;

endmodule // vdp_comp_strong

module vdp_neg_dff (  Q, C, D, R);

	output wire Q;
	input wire C;
	input wire D;
	input wire R;

endmodule // vdp_neg_dff

module vdp_buf (  Z, A);

	output wire Z;
	input wire A;

endmodule // vdp_buf

module vdp_aon2x8 (  Z, A1, B1, C1, D2, A2, B2, C2, D1, E2, F1, E1, F2, G1, H2, G2, H1);

	output wire Z;
	input wire A1;
	input wire B1;
	input wire C1;
	input wire D2;
	input wire A2;
	input wire B2;
	input wire C2;
	input wire D1;
	input wire E2;
	input wire F1;
	input wire E1;
	input wire F2;
	input wire G1;
	input wire H2;
	input wire G2;
	input wire H1;

endmodule // vdp_aon2x8

module vdp_xnor (  Z, A, B);

	output wire Z;
	input wire A;
	input wire B;

endmodule // vdp_xnor

module vdp_oai211 (  Z, A1, A2, B, C);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire B;
	input wire C;

endmodule // vdp_oai211

module vdp_aoi31 (  Z, B3, B2, B1, A);

	output wire Z;
	input wire B3;
	input wire B2;
	input wire B1;
	input wire A;

endmodule // vdp_aoi31

module vdp_AOI222 (  Z, B1, A1, B2, A2, C1, C2);

	output wire Z;
	input wire B1;
	input wire A1;
	input wire B2;
	input wire A2;
	input wire C1;
	input wire C2;

endmodule // vdp_AOI222

module vdp_cnt_bit_rev (  nC2, nC1, C2, C1, Q, CI, B, A);

	input wire nC2;
	input wire nC1;
	input wire C2;
	input wire C1;
	output wire Q;
	input wire CI;
	input wire B;
	input wire A;

endmodule // vdp_cnt_bit_rev

module vdp_2x_sr_bit (  Q, D, nC2, nC1, C2, C1, nC4, nC3, C4, C3);

	output wire Q;
	input wire D;
	input wire nC2;
	input wire nC1;
	input wire C2;
	input wire C1;
	input wire nC4;
	input wire nC3;
	input wire C4;
	input wire C3;

endmodule // vdp_2x_sr_bit

module vdp_and9 (  Z, B, A, C, D, F, E, G, H, I);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;
	input wire I;

endmodule // vdp_and9

module vdp_nor12 (  Z, B, A, C, D, F, E, G, H, J, I, K, L);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;
	input wire J;
	input wire I;
	input wire K;
	input wire L;

endmodule // vdp_nor12

module vdp_nor8 (  Z, B, A, C, D, F, E, G, H);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;

endmodule // vdp_nor8

module vdp_aon21_sr (  Q, A1, A2, B, nC2, nC1, C2, C1);

	output wire Q;
	input wire A1;
	input wire A2;
	input wire B;
	input wire nC2;
	input wire nC1;
	input wire C2;
	input wire C1;

endmodule // vdp_aon21_sr

module vdp_or9 (  Z, B, A, C, D, F, E, G, H, I);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;
	input wire I;

endmodule // vdp_or9

module vdp_V_PLA (  o[0], o[1], o[2], o[3], o[4], o[5], o[6], o[7], o[8], o[9], o[10], o[11], o[12], o[13], o[14], o[15], o[16], o[17], o[18], o[19], o[20], o[21], o[22], o[23], o[24], o[25], o[26], o[27], o[28], o[29], o[30], o[31], o[32], o[33], o[34], o[35], o[36], o[37], o[38], o[39], o[40], o[41], o[42], o[43], o[44], o[45], o[46], o[47], Vcnt[0], Vcnt[1], Vcnt[2], Vcnt[3], Vcnt[4], Vcnt[5], Vcnt[6], Vcnt[7], Vcnt[8], ODD_EVEN, LS0, PAL, nPAL, 2, 3, M5);

	output wire o[0];
	output wire o[1];
	output wire o[2];
	output wire o[3];
	output wire o[4];
	output wire o[5];
	output wire o[6];
	output wire o[7];
	output wire o[8];
	output wire o[9];
	output wire o[10];
	output wire o[11];
	output wire o[12];
	output wire o[13];
	output wire o[14];
	output wire o[15];
	output wire o[16];
	output wire o[17];
	output wire o[18];
	output wire o[19];
	output wire o[20];
	output wire o[21];
	output wire o[22];
	output wire o[23];
	output wire o[24];
	output wire o[25];
	output wire o[26];
	output wire o[27];
	output wire o[28];
	output wire o[29];
	output wire o[30];
	output wire o[31];
	output wire o[32];
	output wire o[33];
	output wire o[34];
	output wire o[35];
	output wire o[36];
	output wire o[37];
	output wire o[38];
	output wire o[39];
	output wire o[40];
	output wire o[41];
	output wire o[42];
	output wire o[43];
	output wire o[44];
	output wire o[45];
	output wire o[46];
	output wire o[47];
	input wire Vcnt[0];
	input wire Vcnt[1];
	input wire Vcnt[2];
	input wire Vcnt[3];
	input wire Vcnt[4];
	input wire Vcnt[5];
	input wire Vcnt[6];
	input wire Vcnt[7];
	input wire Vcnt[8];
	input wire ODD_EVEN;
	input wire LS0;
	input wire PAL;
	input wire nPAL;
	input wire 2;
	input wire 3;
	input wire M5;

endmodule // vdp_V_PLA

module vdp_cram (  q[8], D[8], q[7], D[7], q[6], D[6], q[5], D[5], q[4], D[4], q[3], D[3], q[2], D[2], q[1], D[1], q[0], D[0], A[0], A[1], CLK, A[2], A[3], A[4], A[5], B, A);

	output wire q[8];
	input wire D[8];
	output wire q[7];
	input wire D[7];
	output wire q[6];
	input wire D[6];
	output wire q[5];
	input wire D[5];
	output wire q[4];
	input wire D[4];
	output wire q[3];
	input wire D[3];
	output wire q[2];
	input wire D[2];
	output wire q[1];
	input wire D[1];
	output wire q[0];
	input wire D[0];
	input wire A[0];
	input wire A[1];
	input wire CLK;
	input wire A[2];
	input wire A[3];
	input wire A[4];
	input wire A[5];
	input wire B;
	input wire A;

endmodule // vdp_cram

module vdp_linebuf_ram (  q[0], D[0], q[1], D[1], q[2], D[2], q[3], D[3], q[4], D[4], q[5], D[5], q[6], D[6], q[7], D[7], q[8], D[8], q[9], D[9], q[10], D[10], q[11], D[11], q[12], D[12], q[13], D[13], q[14], D[14], q[15], D[15], q[16], D[16], q[17], D[17], q[18], D[18], q[19], D[19], q[20], D[20], q[21], D[21], q[22], D[22], q[23], D[23], q[24], D[24], q[25], D[25], q[26], D[26], q[27], D[27], CLK, A[5], A[4], A[3], A[2], A[1], A[0], A, B, C, D);

	output wire q[0];
	input wire D[0];
	output wire q[1];
	input wire D[1];
	output wire q[2];
	input wire D[2];
	output wire q[3];
	input wire D[3];
	output wire q[4];
	input wire D[4];
	output wire q[5];
	input wire D[5];
	output wire q[6];
	input wire D[6];
	output wire q[7];
	input wire D[7];
	output wire q[8];
	input wire D[8];
	output wire q[9];
	input wire D[9];
	output wire q[10];
	input wire D[10];
	output wire q[11];
	input wire D[11];
	output wire q[12];
	input wire D[12];
	output wire q[13];
	input wire D[13];
	output wire q[14];
	input wire D[14];
	output wire q[15];
	input wire D[15];
	output wire q[16];
	input wire D[16];
	output wire q[17];
	input wire D[17];
	output wire q[18];
	input wire D[18];
	output wire q[19];
	input wire D[19];
	output wire q[20];
	input wire D[20];
	output wire q[21];
	input wire D[21];
	output wire q[22];
	input wire D[22];
	output wire q[23];
	input wire D[23];
	output wire q[24];
	input wire D[24];
	output wire q[25];
	input wire D[25];
	output wire q[26];
	input wire D[26];
	output wire q[27];
	input wire D[27];
	input wire CLK;
	input wire A[5];
	input wire A[4];
	input wire A[3];
	input wire A[2];
	input wire A[1];
	input wire A[0];
	input wire A;
	input wire B;
	input wire C;
	input wire D;

endmodule // vdp_linebuf_ram

module vdp_att_cashe_ram2 (  q[0], D[0], q[1], D[1], q[2], D[2], q[3], D[3], q[4], D[4], q[5], D[5], q[6], D[6], q[7], D[7], q[8], D[8], q[9], D[9], q[10], D[10], CLK, A[6], A[5], A[1], A[0], A[4], A[3], A[2], A, B);

	output wire q[0];
	input wire D[0];
	output wire q[1];
	input wire D[1];
	output wire q[2];
	input wire D[2];
	output wire q[3];
	input wire D[3];
	output wire q[4];
	input wire D[4];
	output wire q[5];
	input wire D[5];
	output wire q[6];
	input wire D[6];
	output wire q[7];
	input wire D[7];
	output wire q[8];
	input wire D[8];
	output wire q[9];
	input wire D[9];
	output wire q[10];
	input wire D[10];
	input wire CLK;
	input wire A[6];
	input wire A[5];
	input wire A[1];
	input wire A[0];
	input wire A[4];
	input wire A[3];
	input wire A[2];
	input wire A;
	input wire B;

endmodule // vdp_att_cashe_ram2

module vdp_att_cashe_ram1 (  q[0], D[0], q[1], D[1], q[2], D[2], q[3], D[3], q[4], D[4], q[5], D[5], q[6], D[6], q[7], D[7], q[8], D[8], q[9], D[9], CLK, A[0], A[1], A[2], A[3], A[4], A[5], A[6], A, B);

	output wire q[0];
	input wire D[0];
	output wire q[1];
	input wire D[1];
	output wire q[2];
	input wire D[2];
	output wire q[3];
	input wire D[3];
	output wire q[4];
	input wire D[4];
	output wire q[5];
	input wire D[5];
	output wire q[6];
	input wire D[6];
	output wire q[7];
	input wire D[7];
	output wire q[8];
	input wire D[8];
	output wire q[9];
	input wire D[9];
	input wire CLK;
	input wire A[0];
	input wire A[1];
	input wire A[2];
	input wire A[3];
	input wire A[4];
	input wire A[5];
	input wire A[6];
	input wire A;
	input wire B;

endmodule // vdp_att_cashe_ram1

module vdp_att_temp_ram (  A[4], A[0], A[1], A[2], A[3], q[0], D[0], q[1], D[1], q[2], D[2], q[3], D[3], q[4], D[4], q[5], D[5], q[6], D[6], q[7], D[7], q[8], D[8], q[9], D[9], q[10], D[10], q[11], D[11], q[12], D[12], q[13], D[13], q[14], D[14], q[15], D[15], q[16], D[16], q[17], D[17], q[18], D[18], q[19], D[19], q[20], D[20], q[21], D[21], q[22], D[22], q[23], D[23], q[24], D[24], q[25], D[25], q[26], D[26], q[26], D[26], q[27], D[27], q[28], D[28], q[29], D[29], q[30], D[30], q[31], D[31], q[32], D[32], CLK, A, B, C);

	input wire A[4];
	input wire A[0];
	input wire A[1];
	input wire A[2];
	input wire A[3];
	output wire q[0];
	input wire D[0];
	output wire q[1];
	input wire D[1];
	output wire q[2];
	input wire D[2];
	output wire q[3];
	input wire D[3];
	output wire q[4];
	input wire D[4];
	output wire q[5];
	input wire D[5];
	output wire q[6];
	input wire D[6];
	output wire q[7];
	input wire D[7];
	output wire q[8];
	input wire D[8];
	output wire q[9];
	input wire D[9];
	output wire q[10];
	input wire D[10];
	output wire q[11];
	input wire D[11];
	output wire q[12];
	input wire D[12];
	output wire q[13];
	input wire D[13];
	output wire q[14];
	input wire D[14];
	output wire q[15];
	input wire D[15];
	output wire q[16];
	input wire D[16];
	output wire q[17];
	input wire D[17];
	output wire q[18];
	input wire D[18];
	output wire q[19];
	input wire D[19];
	output wire q[20];
	input wire D[20];
	output wire q[21];
	input wire D[21];
	output wire q[22];
	input wire D[22];
	output wire q[23];
	input wire D[23];
	output wire q[24];
	input wire D[24];
	output wire q[25];
	input wire D[25];
	output wire q[26];
	input wire D[26];
	output wire q[26];
	input wire D[26];
	output wire q[27];
	input wire D[27];
	output wire q[28];
	input wire D[28];
	output wire q[29];
	input wire D[29];
	output wire q[30];
	input wire D[30];
	output wire q[31];
	input wire D[31];
	output wire q[32];
	input wire D[32];
	input wire CLK;
	input wire A;
	input wire B;
	input wire C;

endmodule // vdp_att_temp_ram

module vdp_vsram (  CLK, D[10], q[10], D[9], q[9], D[8], q[8], D[7], q[7], D[6], q[6], D[5], q[5], D[4], q[4], D[3], q[3], D[2], q[2], D[1], q[1], D[0], q[0], A[1], A[2], A[3], A[4], A[5], A[0], A, B);

	input wire CLK;
	input wire D[10];
	output wire q[10];
	input wire D[9];
	output wire q[9];
	input wire D[8];
	output wire q[8];
	input wire D[7];
	output wire q[7];
	input wire D[6];
	output wire q[6];
	input wire D[5];
	output wire q[5];
	input wire D[4];
	output wire q[4];
	input wire D[3];
	output wire q[3];
	input wire D[2];
	output wire q[2];
	input wire D[1];
	output wire q[1];
	input wire D[0];
	output wire q[0];
	input wire A[1];
	input wire A[2];
	input wire A[3];
	input wire A[4];
	input wire A[5];
	input wire A[0];
	input wire A;
	input wire B;

endmodule // vdp_vsram

module vdp_H_PLA (  HPLA[0], HPLA[1], HPLA[2], HPLA[3], HPLA[4], HPLA[5], HPLA[7], HPLA[8], HPLA[9], HPLA[6], HPLA[10], HPLA[11], HPLA[16], HPLA[15], HPLA[14], HPLA[13], HPLA[12], i0, HPLA[17], HPLA[18], HPLA[19], HPLA[20], HPLA[21], HPLA[22], Hcnt[0], Hcnt[1], Hcnt[2], Hcnt[3], Hcnt[4], Hcnt[5], Hcnt[6], Hcnt[7], Hcnt[8], H40, M5, B, C, A, HPLA[23], HPLA[24], HPLA[25], HPLA[26], HPLA[27], HPLA[28], HPLA[29], HPLA[30], HPLA[31], HPLA[32], HPLA[33], 3, HPLA[35], HPLA[36], HPLA[34]);

	output wire HPLA[0];
	output wire HPLA[1];
	output wire HPLA[2];
	output wire HPLA[3];
	output wire HPLA[4];
	output wire HPLA[5];
	output wire HPLA[7];
	output wire HPLA[8];
	output wire HPLA[9];
	output wire HPLA[6];
	output wire HPLA[10];
	output wire HPLA[11];
	output wire HPLA[16];
	output wire HPLA[15];
	output wire HPLA[14];
	output wire HPLA[13];
	output wire HPLA[12];
	input wire i0;
	output wire HPLA[17];
	output wire HPLA[18];
	output wire HPLA[19];
	output wire HPLA[20];
	output wire HPLA[21];
	output wire HPLA[22];
	input wire Hcnt[0];
	input wire Hcnt[1];
	input wire Hcnt[2];
	input wire Hcnt[3];
	input wire Hcnt[4];
	input wire Hcnt[5];
	input wire Hcnt[6];
	input wire Hcnt[7];
	input wire Hcnt[8];
	input wire H40;
	input wire M5;
	input wire B;
	input wire C;
	input wire A;
	output wire HPLA[23];
	output wire HPLA[24];
	output wire HPLA[25];
	output wire HPLA[26];
	output wire HPLA[27];
	output wire HPLA[28];
	output wire HPLA[29];
	output wire HPLA[30];
	output wire HPLA[31];
	output wire HPLA[32];
	output wire HPLA[33];
	input wire 3;
	output wire HPLA[35];
	output wire HPLA[36];
	output wire HPLA[34];

endmodule // vdp_H_PLA



// ERROR: conflicting wire AD_DATA[7]
// ERROR: conflicting wire AD_DATA[6]
// ERROR: conflicting wire AD_DATA[4]
// ERROR: conflicting wire RD_DATA[2]
// ERROR: conflicting wire RD_DATA[1]
// ERROR: conflicting wire RD_DATA[0]
// ERROR: conflicting wire AD_DATA[5]
// ERROR: conflicting wire DB[0]
// ERROR: conflicting wire DB[1]
// ERROR: conflicting wire DB[2]
// ERROR: conflicting wire DB[3]
// ERROR: conflicting wire DB[4]
// ERROR: conflicting wire DB[5]
// ERROR: conflicting wire DB[6]
// ERROR: conflicting wire DB[7]
// ERROR: conflicting wire DB[8]
// ERROR: conflicting wire DB[9]
// ERROR: conflicting wire AD_DATA[3]
// ERROR: conflicting wire AD_DATA[2]
// ERROR: conflicting wire AD_DATA[1]
// ERROR: conflicting wire AD_DATA[0]
// ERROR: conflicting wire DB[14]
// ERROR: conflicting wire DB[13]
// ERROR: conflicting wire DB[12]
// ERROR: conflicting wire DB[11]
// ERROR: conflicting wire DB[10]
// ERROR: floating wire w188
// ERROR: conflicting wire RD_DATA[4]
// ERROR: floating wire w219
// ERROR: conflicting wire RD_DATA[6]
// ERROR: floating wire w235
// ERROR: conflicting wire w237
// ERROR: conflicting wire w245
// ERROR: conflicting wire w254
// ERROR: conflicting wire w262
// ERROR: conflicting wire w279
// ERROR: conflicting wire w288
// ERROR: conflicting wire w297
// ERROR: conflicting wire w305
// ERROR: conflicting wire w321
// ERROR: floating wire w334
// ERROR: conflicting wire RD_DATA[5]
// ERROR: floating wire w350
// ERROR: conflicting wire DB[15]
// ERROR: conflicting wire w355
// ERROR: floating wire w457
// ERROR: conflicting wire VRAMA[0]
// ERROR: floating wire w572
// ERROR: conflicting wire VRAMA[8]
// ERROR: conflicting wire VRAMA[7]
// ERROR: conflicting wire VRAMA[9]
// ERROR: conflicting wire VRAMA[10]
// ERROR: conflicting wire VRAMA[6]
// ERROR: conflicting wire VRAMA[5]
// ERROR: conflicting wire VRAMA[11]
// ERROR: conflicting wire VRAMA[12]
// ERROR: conflicting wire VRAMA[4]
// ERROR: conflicting wire VRAMA[13]
// ERROR: conflicting wire VRAMA[3]
// ERROR: conflicting wire VRAMA[14]
// ERROR: conflicting wire VRAMA[2]
// ERROR: conflicting wire CA[14]
// ERROR: conflicting wire VRAMA[15]
// ERROR: conflicting wire VRAMA[1]
// ERROR: conflicting wire VRAMA[16]
// ERROR: floating wire w795
// ERROR: floating wire w797
// ERROR: floating wire w810
// ERROR: floating wire w811
// ERROR: floating wire w1070
// ERROR: conflicting wire COL[0]
// ERROR: conflicting wire COL[1]
// ERROR: conflicting wire COL[2]
// ERROR: conflicting wire COL[3]
// ERROR: conflicting wire COL[4]
// ERROR: conflicting wire COL[5]
// ERROR: conflicting wire COL[6]
// ERROR: floating wire w1092
// ERROR: floating wire w1093
// ERROR: floating wire w1219
// ERROR: floating wire w1292
// ERROR: floating wire w1299
// ERROR: floating wire w1307
// ERROR: floating wire w1324
// ERROR: floating wire w1355
// ERROR: floating wire w1379
// ERROR: floating wire w1600
// ERROR: floating wire w1677
// ERROR: floating wire w1778
// ERROR: floating wire w1808
// ERROR: floating wire w1821
// ERROR: floating wire w1831
// ERROR: floating wire w1975
// ERROR: floating wire w2066
// ERROR: floating wire w2252
// ERROR: floating wire w2287
// ERROR: floating wire w2409
// ERROR: floating wire w2476
// ERROR: floating wire w2622
// ERROR: floating wire w2628
// ERROR: floating wire w2789
// ERROR: floating wire w3104
// ERROR: floating wire w3114
// ERROR: floating wire w3449
// ERROR: floating wire w3519
// ERROR: floating wire w3599
// ERROR: floating wire w3656
// ERROR: floating wire w3697
// ERROR: floating wire w3740
// ERROR: floating wire w3745
// ERROR: floating wire w3800
// ERROR: floating wire w3802
// ERROR: floating wire w3878
// ERROR: floating wire w3904
// ERROR: floating wire w3959
// ERROR: floating wire w4047
// ERROR: floating wire w4079
// ERROR: floating wire w4412
// ERROR: floating wire w4424
// ERROR: floating wire w4579
// ERROR: floating wire w4648
// ERROR: floating wire w4653
// ERROR: floating wire w4691
// ERROR: floating wire w4749
// ERROR: floating wire w4754
// ERROR: floating wire w4783
// ERROR: floating wire w4828
// ERROR: floating wire w4887
// ERROR: floating wire w4902
// ERROR: floating wire w4947
// ERROR: floating wire w5139
// ERROR: floating wire w5195
// ERROR: floating wire w5327
// ERROR: floating wire w5342
// ERROR: floating wire w5346
// ERROR: floating wire w5354
// ERROR: floating wire w5502
// ERROR: floating wire w5550
// ERROR: floating wire w5740
// ERROR: floating wire w5885
// ERROR: floating wire w5887
// ERROR: floating wire w5984
// ERROR: floating wire w6128
// ERROR: floating wire w6144
// ERROR: floating wire w6175
// ERROR: floating wire w6221
// ERROR: floating wire w6267
// ERROR: floating wire w6268
// ERROR: floating wire w6563
// ERROR: floating wire w6678
// ERROR: floating wire w6680
// ERROR: floating wire w6681
// WARNING: Cell vdp_fa:g385 port CO not connected.
// WARNING: Cell vdp_and:g527 port Z not connected.
// WARNING: Cell vdp_cnt_bit_load:g871 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g873 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g1405 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g1406 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1407 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1408 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1409 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1410 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1411 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1412 port Q not connected.
// WARNING: Cell vdp_or:g1576 port Z not connected.
// WARNING: Cell vdp_cnt_bit_load:g1959 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g1960 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2145 port CO not connected.
// WARNING: Cell vdp_ha:g2278 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2280 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2282 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2284 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2286 port CO not connected.
// WARNING: Cell vdp_rs_ff:g2380 port nQ not connected.
// WARNING: Cell vdp_rs_ff:g2381 port nQ not connected.
// WARNING: Cell vdp_comp_we:g2612 port nZ not connected.
// WARNING: Cell vdp_fa:g3842 port CO not connected.
// WARNING: Cell vdp_fa:g4058 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g4437 port CO not connected.
// WARNING: Cell vdp_fa:g4453 port CO not connected.
// WARNING: Cell vdp_fa:g4463 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g5851 port CO not connected.
// WARNING: Cell vdp_fa:g5862 port CO not connected.
// WARNING: Cell vdp_fa:g5888 port CO not connected.
// WARNING: Cell vdp_fa:g5892 port CO not connected.
// WARNING: Cell vdp_fa:g6086 port CO not connected.
// WARNING: Cell vdp_ha:g6137 port CO not connected.
// WARNING: Cell vdp_sr_bit:g6146 port Q not connected.
// WARNING: Cell vdp_fa:g6150 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g6216 port CO not connected.
