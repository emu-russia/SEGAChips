module VDP (  CH0_EN, CH0VOL[0], CH0VOL[1], CH1_EN, CH1VOL[0], CH1VOL[1], CH2_EN, CH2VOL[0], CH2VOL[1], CH3_EN, CH3VOL[0], CH3VOL[1], PSGDAC0[0], PSGDAC0[1], PSGDAC0[2], PSGDAC0[3], PSGDAC0[4], PSGDAC0[5], PSGDAC0[6], PSGDAC0[7], PSGDAC1[0], PSGDAC1[1], PSGDAC1[2], PSGDAC1[3], PSGDAC1[4], PSGDAC1[5], PSGDAC1[6], PSGDAC1[7], PSGDAC2[0], PSGDAC2[1], PSGDAC2[2], PSGDAC2[3], PSGDAC2[4], PSGDAC2[5], PSGDAC2[6], PSGDAC2[7], PSGDAC3[0], PSGDAC3[1], PSGDAC3[2], PSGDAC3[3], PSGDAC3[4], PSGDAC3[5], PSGDAC3[6], PSGDAC3[7], CAi[22], CAo[22], CA[19], DTACK_OUT, Z80_INT, RA[7], RA[6], RA[5], RA[4], RA[2], RA[1], RA[0], nRAS0, RA[3], nCAS0, nOE0, nLWR, nUWR, DTACK_IN, RnW, nLDS, nUDS, nAS, nM1, nWR, nRD, nIORQ, nILP2, nILP1, nINTAK, nMREQ, nBG, BGACK_OUT, BGACK_IN, nBR, VSYNC, nCSYNC, nCSYNC_IN, nHSYNC, nHSYNC_IN, DB[15], DB[14], DB[13], DB[12], DB[11], DB[10], DB[9], DB[8], DB[7], DB[6], DB[5], DB[4], DB[3], DB[2], DB[1], DB[0], CA[0], CA[1], CA[2], CA[3], CA[4], CA[5], CA[6], CA[7], CA[8], CA[9], CA[10], CA[11], CA[12], CA[13], CA[14], CA[15], CA[16], CA[17], CA[18], CA[20], CA[21], R_DAC[0], R_DAC[1], R_DAC[2], R_DAC[3], R_DAC[4], R_DAC[5], R_DAC[6], R_DAC[7], R_DAC[8], G_DAC[0], G_DAC[1], G_DAC[2], G_DAC[3], G_DAC[4], G_DAC[5], G_DAC[6], G_DAC[7], G_DAC[8], R_DAC[9], R_DAC[10], R_DAC[11], R_DAC[12], R_DAC[13], R_DAC[14], R_DAC[15], R_DAC[16], B_DAC[0], B_DAC[1], B_DAC[2], B_DAC[3], B_DAC[4], B_DAC[5], B_DAC[6], B_DAC[7], B_DAC[8], G_DAC[9], G_DAC[10], G_DAC[11], G_DAC[12], G_DAC[13], G_DAC[14], G_DAC[15], G_DAC[16], B_DAC[9], B_DAC[10], B_DAC[11], B_DAC[12], B_DAC[13], B_DAC[14], B_DAC[15], B_DAC[16], nOE1, nWE0, nWE1, nCAS1, nRAS1, AD_RD_DIR, nYS, nSC, nSE0_1, ADo[7], ADo[6], ADo[5], ADo[4], ADo[3], ADo[2], ADo[1], ADo[0], RDo[6], RDo[5], RDo[4], RDo[3], RDo[2], RDo[1], RDo[0], RDi[6], RDi[7], RDi[4], RDi[5], RDi[2], RDi[3], RDi[0], RDi[1], ADi[6], ADi[7], ADi[4], ADi[5], ADi[2], ADi[3], ADi[0], ADi[1], RDo[7], SD[7], SD[6], SD[5], SD[4], SD[3], SD[2], SD[1], SD[0], CLK1, CLK0, EDCLKi, EDCLKo, MCLK, SUB_CLK, nRES_PAD, M68kCLKi, EDCLKd, CA_PAD_DIR, DB_PAD_DIR, SEL0_M3, nPAL, nHL, SPA_Bo, SPA_Bi);

	output wire CH0_EN;
	output wire CH0VOL[0];
	output wire CH0VOL[1];
	output wire CH1_EN;
	output wire CH1VOL[0];
	output wire CH1VOL[1];
	output wire CH2_EN;
	output wire CH2VOL[0];
	output wire CH2VOL[1];
	output wire CH3_EN;
	output wire CH3VOL[0];
	output wire CH3VOL[1];
	output wire PSGDAC0[0];
	output wire PSGDAC0[1];
	output wire PSGDAC0[2];
	output wire PSGDAC0[3];
	output wire PSGDAC0[4];
	output wire PSGDAC0[5];
	output wire PSGDAC0[6];
	output wire PSGDAC0[7];
	output wire PSGDAC1[0];
	output wire PSGDAC1[1];
	output wire PSGDAC1[2];
	output wire PSGDAC1[3];
	output wire PSGDAC1[4];
	output wire PSGDAC1[5];
	output wire PSGDAC1[6];
	output wire PSGDAC1[7];
	output wire PSGDAC2[0];
	output wire PSGDAC2[1];
	output wire PSGDAC2[2];
	output wire PSGDAC2[3];
	output wire PSGDAC2[4];
	output wire PSGDAC2[5];
	output wire PSGDAC2[6];
	output wire PSGDAC2[7];
	output wire PSGDAC3[0];
	output wire PSGDAC3[1];
	output wire PSGDAC3[2];
	output wire PSGDAC3[3];
	output wire PSGDAC3[4];
	output wire PSGDAC3[5];
	output wire PSGDAC3[6];
	output wire PSGDAC3[7];
	input wire CAi[22];
	output wire CAo[22];
	output wire CA[19];
	output wire DTACK_OUT;
	output wire Z80_INT;
	output wire RA[7];
	output wire RA[6];
	output wire RA[5];
	output wire RA[4];
	output wire RA[2];
	output wire RA[1];
	output wire RA[0];
	output wire nRAS0;
	output wire RA[3];
	output wire nCAS0;
	output wire nOE0;
	output wire nLWR;
	output wire nUWR;
	input wire DTACK_IN;
	input wire RnW;
	input wire nLDS;
	input wire nUDS;
	input wire nAS;
	input wire nM1;
	input wire nWR;
	input wire nRD;
	input wire nIORQ;
	output wire nILP2;
	output wire nILP1;
	input wire nINTAK;
	input wire nMREQ;
	input wire nBG;
	output wire BGACK_OUT;
	input wire BGACK_IN;
	output wire nBR;
	output wire VSYNC;
	output wire nCSYNC;
	input wire nCSYNC_IN;
	output wire nHSYNC;
	input wire nHSYNC_IN;
	inout wire DB[15];
	inout wire DB[14];
	inout wire DB[13];
	inout wire DB[12];
	inout wire DB[11];
	inout wire DB[10];
	inout wire DB[9];
	inout wire DB[8];
	inout wire DB[7];
	inout wire DB[6];
	inout wire DB[5];
	inout wire DB[4];
	inout wire DB[3];
	inout wire DB[2];
	inout wire DB[1];
	inout wire DB[0];
	inout wire CA[0];
	inout wire CA[1];
	inout wire CA[2];
	inout wire CA[3];
	inout wire CA[4];
	inout wire CA[5];
	inout wire CA[6];
	inout wire CA[7];
	inout wire CA[8];
	inout wire CA[9];
	inout wire CA[10];
	inout wire CA[11];
	inout wire CA[12];
	inout wire CA[13];
	inout wire CA[14];
	inout wire CA[15];
	inout wire CA[16];
	inout wire CA[17];
	output wire CA[18];
	inout wire CA[20];
	inout wire CA[21];
	output wire R_DAC[0];
	output wire R_DAC[1];
	output wire R_DAC[2];
	output wire R_DAC[3];
	output wire R_DAC[4];
	output wire R_DAC[5];
	output wire R_DAC[6];
	output wire R_DAC[7];
	output wire R_DAC[8];
	output wire G_DAC[0];
	output wire G_DAC[1];
	output wire G_DAC[2];
	output wire G_DAC[3];
	output wire G_DAC[4];
	output wire G_DAC[5];
	output wire G_DAC[6];
	output wire G_DAC[7];
	output wire G_DAC[8];
	output wire R_DAC[9];
	output wire R_DAC[10];
	output wire R_DAC[11];
	output wire R_DAC[12];
	output wire R_DAC[13];
	output wire R_DAC[14];
	output wire R_DAC[15];
	output wire R_DAC[16];
	output wire B_DAC[0];
	output wire B_DAC[1];
	output wire B_DAC[2];
	output wire B_DAC[3];
	output wire B_DAC[4];
	output wire B_DAC[5];
	output wire B_DAC[6];
	output wire B_DAC[7];
	output wire B_DAC[8];
	output wire G_DAC[9];
	output wire G_DAC[10];
	output wire G_DAC[11];
	output wire G_DAC[12];
	output wire G_DAC[13];
	output wire G_DAC[14];
	output wire G_DAC[15];
	output wire G_DAC[16];
	output wire B_DAC[9];
	output wire B_DAC[10];
	output wire B_DAC[11];
	output wire B_DAC[12];
	output wire B_DAC[13];
	output wire B_DAC[14];
	output wire B_DAC[15];
	output wire B_DAC[16];
	output wire nOE1;
	output wire nWE0;
	output wire nWE1;
	output wire nCAS1;
	output wire nRAS1;
	output wire AD_RD_DIR;
	output wire nYS;
	output wire nSC;
	output wire nSE0_1;
	output wire ADo[7];
	output wire ADo[6];
	output wire ADo[5];
	output wire ADo[4];
	output wire ADo[3];
	output wire ADo[2];
	output wire ADo[1];
	output wire ADo[0];
	output wire RDo[6];
	output wire RDo[5];
	output wire RDo[4];
	output wire RDo[3];
	output wire RDo[2];
	output wire RDo[1];
	output wire RDo[0];
	input wire RDi[6];
	input wire RDi[7];
	input wire RDi[4];
	input wire RDi[5];
	input wire RDi[2];
	input wire RDi[3];
	input wire RDi[0];
	input wire RDi[1];
	input wire ADi[6];
	input wire ADi[7];
	input wire ADi[4];
	input wire ADi[5];
	input wire ADi[2];
	input wire ADi[3];
	input wire ADi[0];
	input wire ADi[1];
	output wire RDo[7];
	input wire SD[7];
	input wire SD[6];
	input wire SD[5];
	input wire SD[4];
	input wire SD[3];
	input wire SD[2];
	input wire SD[1];
	input wire SD[0];
	output wire CLK1;
	output wire CLK0;
	input wire EDCLKi;
	output wire EDCLKo;
	input wire MCLK;
	output wire SUB_CLK;
	input wire nRES_PAD;
	input wire M68kCLKi;
	output wire EDCLKd;
	output wire CA_PAD_DIR;
	output wire DB_PAD_DIR;
	input wire SEL0_M3;
	input wire nPAL;
	input wire nHL;
	output wire SPA_Bo;
	input wire SPA_Bi;

	// Wires

	wire w1;
	wire H40;
	wire w3;
	wire w4;
	wire w5;
	wire w6;
	wire w7;
	wire w8;
	wire w9;
	wire w10;
	wire w11;
	wire w12;
	wire w13;
	wire w14;
	wire w15;
	wire w16;
	wire w17;
	wire w18;
	wire w19;
	wire w20;
	wire w21;
	wire w22;
	wire w23;
	wire w24;
	wire w25;
	wire w26;
	wire w27;
	wire w28;
	wire w29;
	wire w30;
	wire w31;
	wire w32;
	wire w33;
	wire w34;
	wire w35;
	wire w36;
	wire w37;
	wire w38;
	wire w39;
	wire w40;
	wire w41;
	wire w42;
	wire w43;
	wire VSCR;
	wire w45;
	wire w46;
	wire w47;
	wire w48;
	wire ODD_EVEN;
	wire w50;
	wire w51;
	wire w52;
	wire w53;
	wire w54;
	wire w55;
	wire w56;
	wire w57;
	wire w58;
	wire w59;
	wire FIFOo[7];
	wire FIFOo[6];
	wire FIFOo[5];
	wire FIFOo[4];
	wire FIFOo[3];
	wire FIFOo[2];
	wire FIFOo[1];
	wire FIFOo[0];
	wire w68;
	wire w69;
	wire w70;
	wire w71;
	wire w72;
	wire w73;
	wire w74;
	wire w75;
	wire w76;
	wire S_TE;
	wire w78;
	wire LSCR;
	wire w80;
	wire HSCR;
	wire w82;
	wire w83;
	wire w84;
	wire w85;
	wire w86;
	wire w87;
	wire w88;
	wire w89;
	wire VPOS[9];
	wire w91;
	wire w92;
	wire w93;
	wire w94;
	wire HPOS[0];
	wire w96;
	wire w97;
	wire w98;
	wire V_INT_HAPPENED;
	wire w100;
	wire w101;
	wire w102;
	wire w103;
	wire VPOS[8];
	wire w105;
	wire w106;
	wire w107;
	wire COLLISION;
	wire w109;
	wire w110;
	wire w111;
	wire w112;
	wire SPRITE_OVF;
	wire w114;
	wire w115;
	wire w116;
	wire w117;
	wire COL[7];
	wire w119;
	wire w120;
	wire w121;
	wire w122;
	wire AD_DATA[7];
	wire AD_DATA[6];
	wire AD_DATA[4];
	wire RD_DATA[2];
	wire RD_DATA[1];
	wire RD_DATA[0];
	wire AD_DATA[5];
	wire DCLK1;
	wire DCLK2;
	wire nDCLK1;
	wire nDCLK2;
	wire HCLK1;
	wire HCLK2;
	wire nHCLK1;
	wire nHCLK2;
	wire SYSRES;
	wire DB[0];
	wire DB[1];
	wire DB[2];
	wire DB[3];
	wire DB[4];
	wire DB[5];
	wire DB[6];
	wire DB[7];
	wire DB[8];
	wire DB[9];
	wire AD_DATA[3];
	wire AD_DATA[2];
	wire AD_DATA[1];
	wire AD_DATA[0];
	wire DB[14];
	wire DB[13];
	wire DB[12];
	wire DB[11];
	wire DB[10];
	wire M5;
	wire w159;
	wire w160;
	wire w161;
	wire w162;
	wire w163;
	wire w164;
	wire w165;
	wire w166;
	wire w167;
	wire w168;
	wire w169;
	wire w170;
	wire w171;
	wire w172;
	wire w173;
	wire VPOS_80;
	wire HPOS[1];
	wire w176;
	wire w177;
	wire w178;
	wire w179;
	wire w180;
	wire w181;
	wire w182;
	wire w183;
	wire w184;
	wire w185;
	wire w186;
	wire w187;
	wire w188;
	wire VPOS[2];
	wire HPOS[3];
	wire w191;
	wire w192;
	wire w193;
	wire w194;
	wire w195;
	wire w196;
	wire w197;
	wire w198;
	wire w199;
	wire w200;
	wire w201;
	wire w202;
	wire w203;
	wire VPOS[4];
	wire w205;
	wire RD_DATA[4];
	wire HPOS[5];
	wire w208;
	wire w209;
	wire w210;
	wire w211;
	wire w212;
	wire w213;
	wire w214;
	wire w215;
	wire w216;
	wire w217;
	wire w218;
	wire w219;
	wire w220;
	wire RD_DATA[6];
	wire HPOS[7];
	wire w223;
	wire w224;
	wire w225;
	wire w226;
	wire w227;
	wire w228;
	wire w229;
	wire w230;
	wire w231;
	wire w232;
	wire w233;
	wire w234;
	wire w235;
	wire w236;
	wire w237;
	wire w238;
	wire w239;
	wire w240;
	wire w241;
	wire w242;
	wire w243;
	wire w244;
	wire w245;
	wire w246;
	wire w247;
	wire w248;
	wire w249;
	wire w250;
	wire w251;
	wire w252;
	wire w253;
	wire w254;
	wire w255;
	wire w256;
	wire w257;
	wire w258;
	wire w259;
	wire w260;
	wire w261;
	wire w262;
	wire w263;
	wire w264;
	wire w265;
	wire w266;
	wire w267;
	wire w268;
	wire w269;
	wire w270;
	wire w271;
	wire w272;
	wire w273;
	wire w274;
	wire w275;
	wire w276;
	wire w277;
	wire w278;
	wire w279;
	wire w280;
	wire w281;
	wire w282;
	wire w283;
	wire w284;
	wire w285;
	wire w286;
	wire w287;
	wire w288;
	wire w289;
	wire w290;
	wire w291;
	wire w292;
	wire w293;
	wire w294;
	wire w295;
	wire w296;
	wire w297;
	wire w298;
	wire w299;
	wire w300;
	wire w301;
	wire w302;
	wire w303;
	wire w304;
	wire w305;
	wire w306;
	wire HPOS[2];
	wire VPOS[1];
	wire w309;
	wire w310;
	wire w311;
	wire w312;
	wire w313;
	wire w314;
	wire w315;
	wire w316;
	wire w317;
	wire w318;
	wire w319;
	wire VPOS[3];
	wire w321;
	wire HPOS[4];
	wire w323;
	wire w324;
	wire w325;
	wire w326;
	wire w327;
	wire w328;
	wire w329;
	wire w330;
	wire w331;
	wire w332;
	wire w333;
	wire w334;
	wire w335;
	wire VPOS[5];
	wire RD_DATA[5];
	wire HPOS[6];
	wire w339;
	wire w340;
	wire w341;
	wire w342;
	wire w343;
	wire w344;
	wire w345;
	wire w346;
	wire w347;
	wire w348;
	wire w349;
	wire w350;
	wire w351;
	wire HPOS[8];
	wire VPOS[7];
	wire DB[15];
	wire w355;
	wire w356;
	wire w357;
	wire w358;
	wire w359;
	wire w360;
	wire w361;
	wire w362;
	wire w363;
	wire w364;
	wire w365;
	wire w366;
	wire w367;
	wire w368;
	wire w369;
	wire w370;
	wire w371;
	wire w372;
	wire w373;
	wire w374;
	wire w375;
	wire w376;
	wire w377;
	wire w378;
	wire w379;
	wire w380;
	wire w381;
	wire w382;
	wire w383;
	wire w384;
	wire w385;
	wire w386;
	wire w387;
	wire w388;
	wire w389;
	wire w390;
	wire w391;
	wire w392;
	wire w393;
	wire w394;
	wire SEL0_M3;
	wire w396;
	wire w397;
	wire w398;
	wire w399;
	wire w400;
	wire w401;
	wire w402;
	wire w403;
	wire w404;
	wire w405;
	wire w406;
	wire w407;
	wire w408;
	wire w409;
	wire w410;
	wire w411;
	wire w412;
	wire w413;
	wire w414;
	wire w415;
	wire w416;
	wire w417;
	wire w418;
	wire w419;
	wire w420;
	wire w421;
	wire w422;
	wire w423;
	wire w424;
	wire VRAM128k;
	wire w426;
	wire w427;
	wire w428;
	wire w429;
	wire w430;
	wire w431;
	wire w432;
	wire w433;
	wire w434;
	wire w435;
	wire w436;
	wire w437;
	wire w438;
	wire w439;
	wire w440;
	wire w441;
	wire w442;
	wire w443;
	wire w444;
	wire w445;
	wire w446;
	wire w447;
	wire w448;
	wire w449;
	wire w450;
	wire w451;
	wire w452;
	wire w453;
	wire w454;
	wire w455;
	wire w456;
	wire w457;
	wire w458;
	wire w459;
	wire w460;
	wire CA[0];
	wire w462;
	wire M3;
	wire w464;
	wire w465;
	wire w466;
	wire w467;
	wire w468;
	wire w469;
	wire w470;
	wire w471;
	wire w472;
	wire w473;
	wire w474;
	wire w475;
	wire w476;
	wire w477;
	wire w478;
	wire w479;
	wire w480;
	wire w481;
	wire w482;
	wire w483;
	wire w484;
	wire w485;
	wire w486;
	wire w487;
	wire w488;
	wire w489;
	wire w490;
	wire w491;
	wire w492;
	wire w493;
	wire w494;
	wire w495;
	wire w496;
	wire w497;
	wire w498;
	wire w499;
	wire w500;
	wire w501;
	wire w502;
	wire w503;
	wire w504;
	wire w505;
	wire w506;
	wire w507;
	wire w508;
	wire w509;
	wire w510;
	wire w511;
	wire w512;
	wire w513;
	wire w514;
	wire w515;
	wire w516;
	wire w517;
	wire w518;
	wire w519;
	wire w520;
	wire w521;
	wire w522;
	wire w523;
	wire w524;
	wire w525;
	wire w526;
	wire w527;
	wire w528;
	wire w529;
	wire w530;
	wire w531;
	wire w532;
	wire w533;
	wire w534;
	wire w535;
	wire w536;
	wire w537;
	wire w538;
	wire w539;
	wire w540;
	wire w541;
	wire w542;
	wire w543;
	wire w544;
	wire w545;
	wire w546;
	wire w547;
	wire w548;
	wire w549;
	wire VRAMA[0];
	wire w551;
	wire w552;
	wire w553;
	wire w554;
	wire w555;
	wire w556;
	wire w557;
	wire w558;
	wire w559;
	wire w560;
	wire w561;
	wire w562;
	wire w563;
	wire w564;
	wire w565;
	wire w566;
	wire w567;
	wire w568;
	wire w569;
	wire w570;
	wire w571;
	wire w572;
	wire w573;
	wire w574;
	wire FIFO_EMPTY;
	wire w576;
	wire w577;
	wire w578;
	wire w579;
	wire w580;
	wire w581;
	wire w582;
	wire w583;
	wire w584;
	wire w585;
	wire DMA_BUSY;
	wire w587;
	wire w588;
	wire w589;
	wire w590;
	wire w591;
	wire w592;
	wire w593;
	wire REG_BUS[0];
	wire w595;
	wire w596;
	wire w597;
	wire REG_BUS[7];
	wire VRAMA[8];
	wire w600;
	wire w601;
	wire w602;
	wire w603;
	wire w604;
	wire w605;
	wire w606;
	wire w607;
	wire w608;
	wire w609;
	wire w610;
	wire w611;
	wire w612;
	wire w613;
	wire w614;
	wire w615;
	wire w616;
	wire w617;
	wire w618;
	wire w619;
	wire w620;
	wire w621;
	wire w622;
	wire w623;
	wire CA[8];
	wire CA[7];
	wire w626;
	wire w627;
	wire w628;
	wire w629;
	wire w630;
	wire w631;
	wire w632;
	wire w633;
	wire w634;
	wire w635;
	wire w636;
	wire w637;
	wire CA[9];
	wire w639;
	wire VRAMA[7];
	wire w641;
	wire REG_BUS[6];
	wire VRAMA[9];
	wire w644;
	wire CA[6];
	wire w646;
	wire w647;
	wire w648;
	wire w649;
	wire w650;
	wire w651;
	wire w652;
	wire w653;
	wire w654;
	wire w655;
	wire w656;
	wire w657;
	wire w658;
	wire w659;
	wire REG_BUS[5];
	wire VRAMA[10];
	wire VRAMA[6];
	wire w663;
	wire REG_BUS[1];
	wire w665;
	wire w666;
	wire w667;
	wire w668;
	wire CA[10];
	wire w670;
	wire w671;
	wire w672;
	wire w673;
	wire w674;
	wire w675;
	wire REG_BUS[2];
	wire w677;
	wire CA[11];
	wire w679;
	wire w680;
	wire w681;
	wire w682;
	wire w683;
	wire w684;
	wire w685;
	wire w686;
	wire w687;
	wire w688;
	wire VRAMA[5];
	wire w690;
	wire w691;
	wire VRAMA[11];
	wire CA[5];
	wire w694;
	wire w695;
	wire REG_BUS[3];
	wire VRAMA[12];
	wire VRAMA[4];
	wire w699;
	wire w700;
	wire w701;
	wire REG_BUS[4];
	wire w703;
	wire CA[12];
	wire w705;
	wire w706;
	wire CA[4];
	wire w708;
	wire w709;
	wire w710;
	wire w711;
	wire CA[19];
	wire w713;
	wire w714;
	wire w715;
	wire w716;
	wire VRAMA[13];
	wire w718;
	wire w719;
	wire w720;
	wire VRAMA[3];
	wire CA[3];
	wire w723;
	wire w724;
	wire CA[13];
	wire CA[20];
	wire w727;
	wire w728;
	wire w729;
	wire w730;
	wire w731;
	wire VRAMA[14];
	wire VRAMA[2];
	wire w734;
	wire w735;
	wire w736;
	wire w737;
	wire w738;
	wire CA[2];
	wire w740;
	wire CA[21];
	wire w742;
	wire w743;
	wire w744;
	wire w745;
	wire w746;
	wire CA[14];
	wire w748;
	wire w749;
	wire VRAMA[15];
	wire CA[15];
	wire VRAMA[1];
	wire w753;
	wire w754;
	wire w755;
	wire w756;
	wire w757;
	wire w758;
	wire w759;
	wire w760;
	wire w761;
	wire w762;
	wire w763;
	wire CA[17];
	wire CA[1];
	wire VRAMA[16];
	wire w767;
	wire w768;
	wire CA[16];
	wire w770;
	wire w771;
	wire w772;
	wire w773;
	wire w774;
	wire w775;
	wire w776;
	wire w777;
	wire w778;
	wire w779;
	wire w780;
	wire w781;
	wire w782;
	wire w783;
	wire w784;
	wire w785;
	wire w786;
	wire w787;
	wire w788;
	wire w789;
	wire w790;
	wire w791;
	wire w792;
	wire w793;
	wire w794;
	wire w795;
	wire w796;
	wire w797;
	wire w798;
	wire w799;
	wire w800;
	wire w801;
	wire w802;
	wire w803;
	wire w804;
	wire w805;
	wire w806;
	wire w807;
	wire w808;
	wire w809;
	wire w810;
	wire w811;
	wire w812;
	wire w813;
	wire w814;
	wire w815;
	wire w816;
	wire w817;
	wire w818;
	wire w819;
	wire w820;
	wire w821;
	wire w822;
	wire w823;
	wire w824;
	wire w825;
	wire w826;
	wire w827;
	wire w828;
	wire w829;
	wire w830;
	wire w831;
	wire w832;
	wire w833;
	wire w834;
	wire w835;
	wire w836;
	wire w837;
	wire w838;
	wire w839;
	wire w840;
	wire w841;
	wire w842;
	wire w843;
	wire w844;
	wire w845;
	wire w846;
	wire w847;
	wire w848;
	wire w849;
	wire w850;
	wire w851;
	wire w852;
	wire w853;
	wire w854;
	wire w855;
	wire w856;
	wire w857;
	wire w858;
	wire w859;
	wire w860;
	wire w861;
	wire w862;
	wire w863;
	wire w864;
	wire w865;
	wire w866;
	wire w867;
	wire w868;
	wire w869;
	wire w870;
	wire w871;
	wire w872;
	wire w873;
	wire w874;
	wire w875;
	wire w876;
	wire w877;
	wire w878;
	wire w879;
	wire w880;
	wire w881;
	wire w882;
	wire w883;
	wire w884;
	wire w885;
	wire w886;
	wire w887;
	wire w888;
	wire w889;
	wire w890;
	wire w891;
	wire w892;
	wire w893;
	wire w894;
	wire w895;
	wire w896;
	wire w897;
	wire w898;
	wire w899;
	wire w900;
	wire w901;
	wire w902;
	wire w903;
	wire w904;
	wire w905;
	wire w906;
	wire w907;
	wire w908;
	wire w909;
	wire w910;
	wire w911;
	wire w912;
	wire w913;
	wire w914;
	wire w915;
	wire w916;
	wire w917;
	wire w918;
	wire w919;
	wire w920;
	wire w921;
	wire w922;
	wire w923;
	wire w924;
	wire w925;
	wire w926;
	wire w927;
	wire w928;
	wire w929;
	wire w930;
	wire w931;
	wire w932;
	wire w933;
	wire w934;
	wire w935;
	wire w936;
	wire w937;
	wire w938;
	wire w939;
	wire w940;
	wire w941;
	wire w942;
	wire w943;
	wire w944;
	wire w945;
	wire w946;
	wire w947;
	wire w948;
	wire w949;
	wire w950;
	wire w951;
	wire w952;
	wire w953;
	wire w954;
	wire w955;
	wire w956;
	wire w957;
	wire w958;
	wire w959;
	wire w960;
	wire w961;
	wire w962;
	wire w963;
	wire w964;
	wire w965;
	wire w966;
	wire w967;
	wire w968;
	wire w969;
	wire w970;
	wire w971;
	wire w972;
	wire w973;
	wire w974;
	wire w975;
	wire w976;
	wire w977;
	wire w978;
	wire w979;
	wire w980;
	wire w981;
	wire w982;
	wire w983;
	wire w984;
	wire w985;
	wire w986;
	wire w987;
	wire w988;
	wire w989;
	wire w990;
	wire w991;
	wire w992;
	wire w993;
	wire w994;
	wire w995;
	wire w996;
	wire w997;
	wire w998;
	wire w999;
	wire w1000;
	wire w1001;
	wire w1002;
	wire w1003;
	wire FIFO_FULL;
	wire w1005;
	wire w1006;
	wire w1007;
	wire w1008;
	wire w1009;
	wire w1010;
	wire w1011;
	wire w1012;
	wire w1013;
	wire w1014;
	wire w1015;
	wire w1016;
	wire w1017;
	wire w1018;
	wire w1019;
	wire w1020;
	wire w1021;
	wire w1022;
	wire PSG_Z80_CLK;
	wire LSM0;
	wire w1025;
	wire VPOS[0];
	wire w1027;
	wire w1028;
	wire w1029;
	wire w1030;
	wire w1031;
	wire w1032;
	wire w1033;
	wire w1034;
	wire w1035;
	wire w1036;
	wire w1037;
	wire w1038;
	wire w1039;
	wire w1040;
	wire w1041;
	wire w1042;
	wire w1043;
	wire w1044;
	wire w1045;
	wire COL[1];
	wire COL[0];
	wire COL[2];
	wire COL[3];
	wire COL[4];
	wire COL[6];
	wire w1052;
	wire w1053;
	wire LSM1;
	wire w1055;
	wire w1056;
	wire COL[5];
	wire w1058;
	wire w1059;
	wire w1060;
	wire w1061;
	wire w1062;
	wire w1063;
	wire w1064;
	wire w1065;
	wire w1066;
	wire w1067;
	wire w1068;
	wire w1069;
	wire w1070;
	wire DISP;
	wire w1072;
	wire w1073;
	wire w1074;
	wire w1075;
	wire w1076;
	wire w1077;
	wire LSM0;
	wire w1079;
	wire M2;
	wire w1081;
	wire w1082;
	wire w1083;
	wire w1084;
	wire w1085;
	wire w1086;
	wire w1087;
	wire w1088;
	wire w1089;
	wire w1090;
	wire w1091;
	wire LSM1;
	wire w1093;
	wire w1094;
	wire w1095;
	wire w1096;
	wire w1097;
	wire w1098;
	wire w1099;
	wire w1100;
	wire w1101;
	wire w1102;
	wire w1103;
	wire w1104;
	wire w1105;
	wire w1106;
	wire IE2;
	wire IE0;
	wire M1;
	wire w1110;
	wire RS0;
	wire PSG_TEST_OE;
	wire w1113;
	wire w1114;
	wire w1115;
	wire w1116;
	wire w1117;
	wire w1118;
	wire w1119;
	wire w1120;
	wire w1121;
	wire w1122;
	wire w1123;
	wire w1124;
	wire w1125;
	wire w1126;
	wire w1127;
	wire w1128;
	wire w1129;
	wire w1130;
	wire w1131;
	wire w1132;
	wire w1133;
	wire w1134;
	wire w1135;
	wire w1136;
	wire w1137;
	wire w1138;
	wire w1139;
	wire w1140;
	wire w1141;
	wire w1142;
	wire w1143;
	wire w1144;
	wire w1145;
	wire w1146;
	wire w1147;
	wire w1148;
	wire w1149;
	wire w1150;
	wire w1151;
	wire w1152;
	wire w1153;
	wire w1154;
	wire w1155;
	wire w1156;
	wire w1157;
	wire w1158;
	wire w1159;
	wire w1160;
	wire PAL;
	wire w1162;
	wire w1163;
	wire w1164;
	wire w1165;
	wire w1166;
	wire w1167;
	wire w1168;
	wire w1169;
	wire w1170;
	wire w1171;
	wire w1172;
	wire w1173;
	wire w1174;
	wire w1175;
	wire w1176;
	wire w1177;
	wire w1178;
	wire w1179;
	wire w1180;
	wire w1181;
	wire w1182;
	wire w1183;
	wire w1184;
	wire w1185;
	wire w1186;
	wire w1187;
	wire w1188;
	wire w1189;
	wire w1190;
	wire w1191;
	wire w1192;
	wire w1193;
	wire w1194;
	wire w1195;
	wire w1196;
	wire w1197;
	wire w1198;
	wire w1199;
	wire w1200;
	wire w1201;
	wire w1202;
	wire w1203;
	wire w1204;
	wire w1205;
	wire w1206;
	wire w1207;
	wire w1208;
	wire w1209;
	wire w1210;
	wire w1211;
	wire w1212;
	wire w1213;
	wire w1214;
	wire w1215;
	wire w1216;
	wire w1217;
	wire w1218;
	wire w1219;
	wire w1220;
	wire w1221;
	wire w1222;
	wire w1223;
	wire w1224;
	wire w1225;
	wire w1226;
	wire w1227;
	wire w1228;
	wire w1229;
	wire w1230;
	wire w1231;
	wire w1232;
	wire w1233;
	wire w1234;
	wire w1235;
	wire w1236;
	wire w1237;
	wire w1238;
	wire w1239;
	wire w1240;
	wire w1241;
	wire w1242;
	wire w1243;
	wire w1244;
	wire w1245;
	wire w1246;
	wire w1247;
	wire w1248;
	wire w1249;
	wire w1250;
	wire w1251;
	wire w1252;
	wire w1253;
	wire w1254;
	wire w1255;
	wire w1256;
	wire w1257;
	wire w1258;
	wire w1259;
	wire w1260;
	wire w1261;
	wire w1262;
	wire w1263;
	wire w1264;
	wire w1265;
	wire w1266;
	wire w1267;
	wire w1268;
	wire w1269;
	wire w1270;
	wire w1271;
	wire w1272;
	wire w1273;
	wire w1274;
	wire w1275;
	wire w1276;
	wire w1277;
	wire w1278;
	wire w1279;
	wire w1280;
	wire w1281;
	wire w1282;
	wire w1283;
	wire w1284;
	wire w1285;
	wire w1286;
	wire w1287;
	wire w1288;
	wire w1289;
	wire w1290;
	wire w1291;
	wire w1292;
	wire w1293;
	wire w1294;
	wire w1295;
	wire w1296;
	wire w1297;
	wire w1298;
	wire w1299;
	wire w1300;
	wire w1301;
	wire w1302;
	wire w1303;
	wire w1304;
	wire w1305;
	wire w1306;
	wire w1307;
	wire w1308;
	wire w1309;
	wire w1310;
	wire w1311;
	wire w1312;
	wire w1313;
	wire w1314;
	wire w1315;
	wire w1316;
	wire w1317;
	wire w1318;
	wire w1319;
	wire w1320;
	wire w1321;
	wire w1322;
	wire w1323;
	wire w1324;
	wire w1325;
	wire w1326;
	wire w1327;
	wire w1328;
	wire w1329;
	wire w1330;
	wire w1331;
	wire w1332;
	wire w1333;
	wire w1334;
	wire w1335;
	wire w1336;
	wire w1337;
	wire w1338;
	wire w1339;
	wire w1340;
	wire w1341;
	wire w1342;
	wire VRAM_REFRESH;
	wire w1344;
	wire w1345;
	wire w1346;
	wire w1347;
	wire w1348;
	wire w1349;
	wire w1350;
	wire w1351;
	wire w1352;
	wire w1353;
	wire w1354;
	wire w1355;
	wire w1356;
	wire w1357;
	wire w1358;
	wire w1359;
	wire w1360;
	wire w1361;
	wire w1362;
	wire w1363;
	wire w1364;
	wire w1365;
	wire w1366;
	wire w1367;
	wire w1368;
	wire w1369;
	wire w1370;
	wire w1371;
	wire w1372;
	wire w1373;
	wire w1374;
	wire w1375;
	wire w1376;
	wire w1377;
	wire w1378;
	wire w1379;
	wire w1380;
	wire w1381;
	wire w1382;
	wire w1383;
	wire w1384;
	wire w1385;
	wire w1386;
	wire w1387;
	wire w1388;
	wire w1389;
	wire w1390;
	wire w1391;
	wire w1392;
	wire w1393;
	wire w1394;
	wire w1395;
	wire w1396;
	wire w1397;
	wire w1398;
	wire w1399;
	wire w1400;
	wire w1401;
	wire w1402;
	wire w1403;
	wire w1404;
	wire w1405;
	wire w1406;
	wire w1407;
	wire w1408;
	wire w1409;
	wire w1410;
	wire w1411;
	wire w1412;
	wire w1413;
	wire w1414;
	wire w1415;
	wire w1416;
	wire w1417;
	wire w1418;
	wire w1419;
	wire w1420;
	wire w1421;
	wire w1422;
	wire w1423;
	wire w1424;
	wire w1425;
	wire w1426;
	wire w1427;
	wire w1428;
	wire w1429;
	wire w1430;
	wire w1431;
	wire w1432;
	wire w1433;
	wire w1434;
	wire w1435;
	wire w1436;
	wire w1437;
	wire w1438;
	wire w1439;
	wire w1440;
	wire w1441;
	wire w1442;
	wire w1443;
	wire w1444;
	wire w1445;
	wire w1446;
	wire w1447;
	wire w1448;
	wire w1449;
	wire w1450;
	wire w1451;
	wire w1452;
	wire w1453;
	wire w1454;
	wire CA[18];
	wire w1456;
	wire w1457;
	wire w1458;
	wire w1459;
	wire w1460;
	wire w1461;
	wire w1462;
	wire w1463;
	wire w1464;
	wire w1465;
	wire w1466;
	wire w1467;
	wire w1468;
	wire w1469;
	wire w1470;
	wire w1471;
	wire w1472;
	wire w1473;
	wire w1474;
	wire w1475;
	wire w1476;
	wire w1477;
	wire w1478;
	wire w1479;
	wire w1480;
	wire w1481;
	wire w1482;
	wire w1483;
	wire w1484;
	wire w1485;
	wire w1486;
	wire w1487;
	wire w1488;
	wire w1489;
	wire w1490;
	wire w1491;
	wire w1492;
	wire w1493;
	wire w1494;
	wire w1495;
	wire w1496;
	wire w1497;
	wire w1498;
	wire w1499;
	wire w1500;
	wire w1501;
	wire w1502;
	wire w1503;
	wire w1504;
	wire w1505;
	wire w1506;
	wire w1507;
	wire w1508;
	wire w1509;
	wire w1510;
	wire w1511;
	wire w1512;
	wire w1513;
	wire w1514;
	wire w1515;
	wire w1516;
	wire VPOS[6];
	wire w1518;
	wire w1519;
	wire w1520;
	wire w1521;
	wire w1522;
	wire w1523;
	wire w1524;
	wire w1525;
	wire w1526;
	wire w1527;
	wire w1528;
	wire w1529;
	wire w1530;
	wire w1531;
	wire w1532;
	wire w1533;
	wire w1534;
	wire w1535;
	wire w1536;
	wire w1537;
	wire w1538;
	wire w1539;
	wire w1540;
	wire w1541;
	wire w1542;
	wire w1543;
	wire w1544;
	wire w1545;
	wire w1546;
	wire w1547;
	wire w1548;
	wire w1549;
	wire w1550;
	wire w1551;
	wire w1552;
	wire w1553;
	wire w1554;
	wire w1555;
	wire w1556;
	wire w1557;
	wire w1558;
	wire w1559;
	wire w1560;
	wire w1561;
	wire w1562;
	wire w1563;
	wire w1564;
	wire w1565;
	wire w1566;
	wire w1567;
	wire w1568;
	wire w1569;
	wire w1570;
	wire w1571;
	wire w1572;
	wire w1573;
	wire w1574;
	wire w1575;
	wire w1576;
	wire w1577;
	wire w1578;
	wire w1579;
	wire w1580;
	wire w1581;
	wire w1582;
	wire w1583;
	wire w1584;
	wire w1585;
	wire w1586;
	wire w1587;
	wire w1588;
	wire w1589;
	wire w1590;
	wire w1591;
	wire w1592;
	wire w1593;
	wire w1594;
	wire w1595;
	wire w1596;
	wire w1597;
	wire VPLA1;
	wire w1599;
	wire w1600;
	wire w1601;
	wire w1602;
	wire w1603;
	wire w1604;
	wire w1605;
	wire w1606;
	wire w1607;
	wire w1608;
	wire w1609;
	wire HPLA29;
	wire HPLA31;
	wire w1612;
	wire w1613;
	wire w1614;
	wire w1615;
	wire w1616;
	wire w1617;
	wire w1618;
	wire w1619;
	wire w1620;
	wire w1621;
	wire w1622;
	wire w1623;
	wire HPLA26;
	wire w1625;
	wire HPLA24;
	wire HPLA25;
	wire HPLA23;
	wire w1629;
	wire w1630;
	wire w1631;
	wire w1632;
	wire w1633;
	wire w1634;
	wire w1635;
	wire w1636;
	wire w1637;
	wire w1638;
	wire w1639;
	wire w1640;
	wire w1641;
	wire w1642;
	wire w1643;
	wire w1644;
	wire w1645;
	wire w1646;
	wire w1647;
	wire w1648;
	wire w1649;
	wire w1650;
	wire w1651;
	wire w1652;
	wire w1653;
	wire w1654;
	wire w1655;
	wire w1656;
	wire w1657;
	wire w1658;
	wire w1659;
	wire w1660;
	wire w1661;
	wire w1662;
	wire HPLA30;
	wire w1664;
	wire w1665;
	wire w1666;
	wire w1667;
	wire w1668;
	wire w1669;
	wire w1670;
	wire w1671;
	wire w1672;
	wire w1673;
	wire w1674;
	wire w1675;
	wire w1676;
	wire w1677;
	wire w1678;
	wire w1679;
	wire w1680;
	wire w1681;
	wire w1682;
	wire w1683;
	wire w1684;
	wire w1685;
	wire HPLA3;
	wire HPLA7;
	wire HPLA8;
	wire HPLA6;
	wire w1690;
	wire w1691;
	wire w1692;
	wire w1693;
	wire w1694;
	wire w1695;
	wire w1696;
	wire w1697;
	wire w1698;
	wire w1699;
	wire w1700;
	wire HPLA36;
	wire w1702;
	wire HPLA33;
	wire w1704;
	wire w1705;
	wire w1706;
	wire w1707;
	wire HPLA18;
	wire HPLA17;
	wire w1710;
	wire w1711;
	wire w1712;
	wire w1713;
	wire w1714;
	wire w1715;
	wire w1716;
	wire w1717;
	wire w1718;
	wire w1719;
	wire w1720;
	wire w1721;
	wire w1722;
	wire w1723;
	wire w1724;
	wire w1725;
	wire w1726;
	wire w1727;
	wire w1728;
	wire w1729;
	wire w1730;
	wire w1731;
	wire w1732;
	wire w1733;
	wire w1734;
	wire w1735;
	wire w1736;
	wire HPLA35;
	wire w1738;
	wire w1739;
	wire w1740;
	wire w1741;
	wire w1742;
	wire w1743;
	wire w1744;
	wire w1745;
	wire w1746;
	wire w1747;
	wire w1748;
	wire w1749;
	wire w1750;
	wire w1751;
	wire w1752;
	wire w1753;
	wire w1754;
	wire w1755;
	wire w1756;
	wire VPLA0;
	wire VPLA2;
	wire VPLA3;
	wire w1760;
	wire w1761;
	wire w1762;
	wire w1763;
	wire w1764;
	wire w1765;
	wire w1766;
	wire VPLA7;
	wire VPLA6;
	wire VPLA5;
	wire VPLA4;
	wire w1771;
	wire w1772;
	wire w1773;
	wire w1774;
	wire w1775;
	wire w1776;
	wire w1777;
	wire w1778;
	wire w1779;
	wire w1780;
	wire w1781;
	wire w1782;
	wire w1783;
	wire w1784;
	wire w1785;
	wire w1786;
	wire w1787;
	wire w1788;
	wire w1789;
	wire w1790;
	wire w1791;
	wire w1792;
	wire w1793;
	wire w1794;
	wire HPLA28;
	wire w1796;
	wire HPLA9;
	wire HPLA20;
	wire HPLA19;
	wire HPLA10;
	wire HPLA16;
	wire HPLA27;
	wire w1803;
	wire w1804;
	wire w1805;
	wire w1806;
	wire w1807;
	wire w1808;
	wire w1809;
	wire w1810;
	wire w1811;
	wire w1812;
	wire w1813;
	wire w1814;
	wire w1815;
	wire w1816;
	wire w1817;
	wire w1818;
	wire w1819;
	wire w1820;
	wire w1821;
	wire w1822;
	wire w1823;
	wire w1824;
	wire w1825;
	wire w1826;
	wire w1827;
	wire w1828;
	wire w1829;
	wire w1830;
	wire w1831;
	wire HPLA22;
	wire HPLA4;
	wire HPLA32;
	wire HPLA2;
	wire HPLA5;
	wire HPLA21;
	wire w1838;
	wire HPLA11;
	wire HPLA14;
	wire HPLA15;
	wire w1842;
	wire HPLA1;
	wire HPLA13;
	wire HPLA12;
	wire w1846;
	wire w1847;
	wire w1848;
	wire w1849;
	wire w1850;
	wire w1851;
	wire w1852;
	wire w1853;
	wire w1854;
	wire w1855;
	wire w1856;
	wire w1857;
	wire w1858;
	wire w1859;
	wire w1860;
	wire w1861;
	wire HPLA0;
	wire w1863;
	wire HPLA34;
	wire w1865;
	wire w1866;
	wire w1867;
	wire w1868;
	wire w1869;
	wire w1870;
	wire w1871;
	wire w1872;
	wire w1873;
	wire w1874;
	wire w1875;
	wire w1876;
	wire w1877;
	wire w1878;
	wire w1879;
	wire w1880;
	wire w1881;
	wire w1882;
	wire w1883;
	wire w1884;
	wire w1885;
	wire w1886;
	wire w1887;
	wire w1888;
	wire w1889;
	wire w1890;
	wire w1891;
	wire w1892;
	wire w1893;
	wire w1894;
	wire w1895;
	wire w1896;
	wire w1897;
	wire w1898;
	wire w1899;
	wire w1900;
	wire w1901;
	wire w1902;
	wire w1903;
	wire w1904;
	wire w1905;
	wire w1906;
	wire w1907;
	wire w1908;
	wire w1909;
	wire w1910;
	wire w1911;
	wire w1912;
	wire w1913;
	wire w1914;
	wire w1915;
	wire w1916;
	wire w1917;
	wire w1918;
	wire w1919;
	wire w1920;
	wire w1921;
	wire w1922;
	wire w1923;
	wire w1924;
	wire w1925;
	wire w1926;
	wire w1927;
	wire w1928;
	wire w1929;
	wire w1930;
	wire w1931;
	wire w1932;
	wire w1933;
	wire w1934;
	wire w1935;
	wire w1936;
	wire w1937;
	wire w1938;
	wire w1939;
	wire w1940;
	wire w1941;
	wire w1942;
	wire w1943;
	wire w1944;
	wire w1945;
	wire w1946;
	wire w1947;
	wire w1948;
	wire w1949;
	wire w1950;
	wire w1951;
	wire w1952;
	wire w1953;
	wire w1954;
	wire w1955;
	wire w1956;
	wire w1957;
	wire w1958;
	wire w1959;
	wire w1960;
	wire w1961;
	wire w1962;
	wire w1963;
	wire w1964;
	wire w1965;
	wire w1966;
	wire w1967;
	wire w1968;
	wire w1969;
	wire w1970;
	wire w1971;
	wire w1972;
	wire w1973;
	wire w1974;
	wire w1975;
	wire w1976;
	wire w1977;
	wire w1978;
	wire w1979;
	wire w1980;
	wire w1981;
	wire w1982;
	wire w1983;
	wire w1984;
	wire w1985;
	wire w1986;
	wire w1987;
	wire w1988;
	wire w1989;
	wire w1990;
	wire w1991;
	wire w1992;
	wire w1993;
	wire w1994;
	wire w1995;
	wire w1996;
	wire w1997;
	wire w1998;
	wire w1999;
	wire w2000;
	wire w2001;
	wire w2002;
	wire w2003;
	wire w2004;
	wire w2005;
	wire w2006;
	wire w2007;
	wire w2008;
	wire w2009;
	wire w2010;
	wire w2011;
	wire w2012;
	wire w2013;
	wire w2014;
	wire w2015;
	wire w2016;
	wire w2017;
	wire w2018;
	wire w2019;
	wire w2020;
	wire w2021;
	wire w2022;
	wire w2023;
	wire w2024;
	wire w2025;
	wire w2026;
	wire w2027;
	wire w2028;
	wire w2029;
	wire w2030;
	wire w2031;
	wire w2032;
	wire w2033;
	wire w2034;
	wire w2035;
	wire w2036;
	wire w2037;
	wire w2038;
	wire w2039;
	wire w2040;
	wire w2041;
	wire w2042;
	wire w2043;
	wire w2044;
	wire w2045;
	wire w2046;
	wire w2047;
	wire w2048;
	wire w2049;
	wire w2050;
	wire w2051;
	wire w2052;
	wire w2053;
	wire w2054;
	wire w2055;
	wire w2056;
	wire w2057;
	wire w2058;
	wire w2059;
	wire w2060;
	wire w2061;
	wire w2062;
	wire w2063;
	wire w2064;
	wire w2065;
	wire w2066;
	wire w2067;
	wire w2068;
	wire w2069;
	wire w2070;
	wire w2071;
	wire w2072;
	wire w2073;
	wire w2074;
	wire w2075;
	wire w2076;
	wire w2077;
	wire w2078;
	wire w2079;
	wire w2080;
	wire w2081;
	wire w2082;
	wire w2083;
	wire w2084;
	wire w2085;
	wire w2086;
	wire w2087;
	wire w2088;
	wire w2089;
	wire w2090;
	wire w2091;
	wire w2092;
	wire w2093;
	wire w2094;
	wire w2095;
	wire w2096;
	wire w2097;
	wire w2098;
	wire w2099;
	wire w2100;
	wire w2101;
	wire w2102;
	wire w2103;
	wire w2104;
	wire w2105;
	wire w2106;
	wire w2107;
	wire w2108;
	wire w2109;
	wire w2110;
	wire w2111;
	wire w2112;
	wire w2113;
	wire w2114;
	wire w2115;
	wire w2116;
	wire w2117;
	wire w2118;
	wire w2119;
	wire w2120;
	wire w2121;
	wire w2122;
	wire w2123;
	wire w2124;
	wire PSG_CLK2;
	wire PSG_CLK1;
	wire w2127;
	wire w2128;
	wire w2129;
	wire w2130;
	wire w2131;
	wire w2132;
	wire w2133;
	wire w2134;
	wire PSG_nCLK2;
	wire PSG_nCLK1;
	wire w2137;
	wire w2138;
	wire w2139;
	wire w2140;
	wire w2141;
	wire w2142;
	wire w2143;
	wire w2144;
	wire w2145;
	wire w2146;
	wire w2147;
	wire w2148;
	wire w2149;
	wire w2150;
	wire w2151;
	wire w2152;
	wire w2153;
	wire w2154;
	wire w2155;
	wire w2156;
	wire w2157;
	wire w2158;
	wire w2159;
	wire w2160;
	wire w2161;
	wire w2162;
	wire w2163;
	wire w2164;
	wire w2165;
	wire w2166;
	wire w2167;
	wire w2168;
	wire w2169;
	wire w2170;
	wire w2171;
	wire w2172;
	wire w2173;
	wire w2174;
	wire w2175;
	wire w2176;
	wire w2177;
	wire w2178;
	wire w2179;
	wire w2180;
	wire w2181;
	wire w2182;
	wire w2183;
	wire w2184;
	wire w2185;
	wire w2186;
	wire w2187;
	wire w2188;
	wire w2189;
	wire w2190;
	wire w2191;
	wire w2192;
	wire w2193;
	wire w2194;
	wire w2195;
	wire w2196;
	wire w2197;
	wire w2198;
	wire w2199;
	wire w2200;
	wire w2201;
	wire w2202;
	wire w2203;
	wire w2204;
	wire w2205;
	wire w2206;
	wire w2207;
	wire w2208;
	wire w2209;
	wire w2210;
	wire w2211;
	wire w2212;
	wire w2213;
	wire w2214;
	wire w2215;
	wire w2216;
	wire w2217;
	wire w2218;
	wire w2219;
	wire w2220;
	wire w2221;
	wire w2222;
	wire w2223;
	wire w2224;
	wire w2225;
	wire w2226;
	wire w2227;
	wire w2228;
	wire w2229;
	wire w2230;
	wire w2231;
	wire w2232;
	wire w2233;
	wire w2234;
	wire w2235;
	wire w2236;
	wire w2237;
	wire w2238;
	wire w2239;
	wire w2240;
	wire w2241;
	wire w2242;
	wire w2243;
	wire w2244;
	wire w2245;
	wire w2246;
	wire w2247;
	wire w2248;
	wire w2249;
	wire w2250;
	wire w2251;
	wire w2252;
	wire w2253;
	wire w2254;
	wire w2255;
	wire w2256;
	wire w2257;
	wire w2258;
	wire w2259;
	wire w2260;
	wire w2261;
	wire w2262;
	wire w2263;
	wire w2264;
	wire w2265;
	wire w2266;
	wire w2267;
	wire w2268;
	wire w2269;
	wire w2270;
	wire w2271;
	wire w2272;
	wire w2273;
	wire w2274;
	wire w2275;
	wire w2276;
	wire w2277;
	wire w2278;
	wire w2279;
	wire w2280;
	wire w2281;
	wire w2282;
	wire w2283;
	wire w2284;
	wire w2285;
	wire w2286;
	wire w2287;
	wire w2288;
	wire w2289;
	wire w2290;
	wire w2291;
	wire w2292;
	wire w2293;
	wire w2294;
	wire w2295;
	wire w2296;
	wire w2297;
	wire w2298;
	wire w2299;
	wire w2300;
	wire w2301;
	wire w2302;
	wire w2303;
	wire w2304;
	wire w2305;
	wire w2306;
	wire w2307;
	wire w2308;
	wire w2309;
	wire w2310;
	wire w2311;
	wire w2312;
	wire w2313;
	wire w2314;
	wire w2315;
	wire w2316;
	wire w2317;
	wire w2318;
	wire w2319;
	wire w2320;
	wire w2321;
	wire w2322;
	wire w2323;
	wire w2324;
	wire w2325;
	wire w2326;
	wire w2327;
	wire w2328;
	wire w2329;
	wire w2330;
	wire w2331;
	wire w2332;
	wire w2333;
	wire w2334;
	wire w2335;
	wire w2336;
	wire w2337;
	wire w2338;
	wire w2339;
	wire w2340;
	wire w2341;
	wire w2342;
	wire w2343;
	wire w2344;
	wire w2345;
	wire w2346;
	wire w2347;
	wire w2348;
	wire w2349;
	wire w2350;
	wire w2351;
	wire w2352;
	wire w2353;
	wire w2354;
	wire w2355;
	wire w2356;
	wire w2357;
	wire w2358;
	wire w2359;
	wire w2360;
	wire w2361;
	wire w2362;
	wire w2363;
	wire w2364;
	wire w2365;
	wire w2366;
	wire w2367;
	wire w2368;
	wire w2369;
	wire w2370;
	wire w2371;
	wire w2372;
	wire w2373;
	wire w2374;
	wire w2375;
	wire w2376;
	wire w2377;
	wire w2378;
	wire w2379;
	wire w2380;
	wire w2381;
	wire w2382;
	wire w2383;
	wire w2384;
	wire w2385;
	wire w2386;
	wire w2387;
	wire w2388;
	wire w2389;
	wire w2390;
	wire w2391;
	wire w2392;
	wire w2393;
	wire w2394;
	wire w2395;
	wire w2396;
	wire w2397;
	wire w2398;
	wire w2399;
	wire w2400;
	wire w2401;
	wire w2402;
	wire w2403;
	wire w2404;
	wire w2405;
	wire w2406;
	wire w2407;
	wire w2408;
	wire w2409;
	wire w2410;
	wire w2411;
	wire w2412;
	wire w2413;
	wire w2414;
	wire w2415;
	wire w2416;
	wire w2417;
	wire w2418;
	wire w2419;
	wire w2420;
	wire w2421;
	wire w2422;
	wire w2423;
	wire w2424;
	wire w2425;
	wire w2426;
	wire w2427;
	wire w2428;
	wire w2429;
	wire w2430;
	wire w2431;
	wire w2432;
	wire w2433;
	wire w2434;
	wire w2435;
	wire w2436;
	wire w2437;
	wire w2438;
	wire w2439;
	wire w2440;
	wire w2441;
	wire w2442;
	wire w2443;
	wire w2444;
	wire w2445;
	wire w2446;
	wire w2447;
	wire w2448;
	wire w2449;
	wire w2450;
	wire w2451;
	wire w2452;
	wire w2453;
	wire w2454;
	wire w2455;
	wire w2456;
	wire w2457;
	wire w2458;
	wire w2459;
	wire w2460;
	wire w2461;
	wire w2462;
	wire w2463;
	wire w2464;
	wire w2465;
	wire w2466;
	wire w2467;
	wire w2468;
	wire w2469;
	wire w2470;
	wire w2471;
	wire w2472;
	wire w2473;
	wire w2474;
	wire w2475;
	wire w2476;
	wire w2477;
	wire w2478;
	wire w2479;
	wire w2480;
	wire w2481;
	wire w2482;
	wire w2483;
	wire w2484;
	wire w2485;
	wire w2486;
	wire w2487;
	wire w2488;
	wire w2489;
	wire w2490;
	wire w2491;
	wire w2492;
	wire w2493;
	wire w2494;
	wire w2495;
	wire w2496;
	wire w2497;
	wire w2498;
	wire w2499;
	wire w2500;
	wire w2501;
	wire w2502;
	wire w2503;
	wire w2504;
	wire w2505;
	wire w2506;
	wire w2507;
	wire w2508;
	wire w2509;
	wire w2510;
	wire w2511;
	wire w2512;
	wire w2513;
	wire w2514;
	wire w2515;
	wire w2516;
	wire w2517;
	wire w2518;
	wire w2519;
	wire w2520;
	wire w2521;
	wire w2522;
	wire w2523;
	wire w2524;
	wire w2525;
	wire w2526;
	wire w2527;
	wire w2528;
	wire w2529;
	wire w2530;
	wire w2531;
	wire w2532;
	wire w2533;
	wire w2534;
	wire w2535;
	wire w2536;
	wire w2537;
	wire w2538;
	wire w2539;
	wire w2540;
	wire w2541;
	wire w2542;
	wire w2543;
	wire RES;
	wire w2545;
	wire w2546;
	wire w2547;
	wire w2548;
	wire EDCLK_O;
	wire nYS;
	wire w2551;
	wire w2552;
	wire w2553;
	wire w2554;
	wire w2555;
	wire w2556;
	wire w2557;
	wire w2558;
	wire w2559;
	wire w2560;
	wire w2561;
	wire w2562;
	wire w2563;
	wire w2564;
	wire w2565;
	wire w2566;
	wire w2567;
	wire w2568;
	wire w2569;
	wire w2570;
	wire w2571;
	wire w2572;
	wire w2573;
	wire w2574;
	wire w2575;
	wire w2576;
	wire w2577;
	wire w2578;
	wire w2579;
	wire w2580;
	wire w2581;
	wire w2582;
	wire w2583;
	wire w2584;
	wire w2585;
	wire w2586;
	wire w2587;
	wire w2588;
	wire w2589;
	wire w2590;
	wire w2591;
	wire w2592;
	wire w2593;
	wire w2594;
	wire w2595;
	wire w2596;
	wire w2597;
	wire w2598;
	wire w2599;
	wire w2600;
	wire w2601;
	wire w2602;
	wire w2603;
	wire w2604;
	wire w2605;
	wire w2606;
	wire w2607;
	wire w2608;
	wire w2609;
	wire SPR_PRIO;
	wire w2611;
	wire w2612;
	wire w2613;
	wire w2614;
	wire w2615;
	wire w2616;
	wire w2617;
	wire w2618;
	wire w2619;
	wire w2620;
	wire w2621;
	wire w2622;
	wire w2623;
	wire w2624;
	wire w2625;
	wire w2626;
	wire w2627;
	wire w2628;
	wire w2629;
	wire w2630;
	wire w2631;
	wire w2632;
	wire w2633;
	wire w2634;
	wire w2635;
	wire w2636;
	wire w2637;
	wire w2638;
	wire w2639;
	wire w2640;
	wire w2641;
	wire w2642;
	wire w2643;
	wire w2644;
	wire w2645;
	wire w2646;
	wire w2647;
	wire w2648;
	wire w2649;
	wire w2650;
	wire w2651;
	wire w2652;
	wire w2653;
	wire w2654;
	wire w2655;
	wire w2656;
	wire w2657;
	wire w2658;
	wire w2659;
	wire w2660;
	wire w2661;
	wire w2662;
	wire w2663;
	wire w2664;
	wire w2665;
	wire w2666;
	wire w2667;
	wire w2668;
	wire w2669;
	wire w2670;
	wire w2671;
	wire w2672;
	wire w2673;
	wire w2674;
	wire w2675;
	wire w2676;
	wire w2677;
	wire PLANE_A_PRIO;
	wire PLANE_B_PRIO;
	wire w2680;
	wire w2681;
	wire w2682;
	wire w2683;
	wire w2684;
	wire w2685;
	wire w2686;
	wire w2687;
	wire w2688;
	wire w2689;
	wire w2690;
	wire w2691;
	wire w2692;
	wire w2693;
	wire w2694;
	wire w2695;
	wire w2696;
	wire w2697;
	wire w2698;
	wire w2699;
	wire w2700;
	wire w2701;
	wire w2702;
	wire w2703;
	wire w2704;
	wire w2705;
	wire w2706;
	wire w2707;
	wire w2708;
	wire w2709;
	wire w2710;
	wire w2711;
	wire w2712;
	wire w2713;
	wire w2714;
	wire w2715;
	wire w2716;
	wire w2717;
	wire w2718;
	wire w2719;
	wire w2720;
	wire w2721;
	wire w2722;
	wire w2723;
	wire w2724;
	wire w2725;
	wire w2726;
	wire w2727;
	wire w2728;
	wire w2729;
	wire w2730;
	wire w2731;
	wire w2732;
	wire w2733;
	wire w2734;
	wire w2735;
	wire w2736;
	wire w2737;
	wire w2738;
	wire w2739;
	wire w2740;
	wire w2741;
	wire w2742;
	wire w2743;
	wire w2744;
	wire w2745;
	wire w2746;
	wire w2747;
	wire w2748;
	wire w2749;
	wire w2750;
	wire w2751;
	wire w2752;
	wire w2753;
	wire w2754;
	wire w2755;
	wire w2756;
	wire w2757;
	wire w2758;
	wire w2759;
	wire w2760;
	wire w2761;
	wire w2762;
	wire HIGHLIGHT;
	wire w2764;
	wire w2765;
	wire w2766;
	wire w2767;
	wire w2768;
	wire w2769;
	wire w2770;
	wire w2771;
	wire w2772;
	wire w2773;
	wire w2774;
	wire w2775;
	wire w2776;
	wire w2777;
	wire w2778;
	wire w2779;
	wire w2780;
	wire w2781;
	wire w2782;
	wire w2783;
	wire w2784;
	wire w2785;
	wire SHADOW;
	wire w2787;
	wire w2788;
	wire w2789;
	wire w2790;
	wire w2791;
	wire w2792;
	wire w2793;
	wire w2794;
	wire w2795;
	wire w2796;
	wire w2797;
	wire w2798;
	wire w2799;
	wire w2800;
	wire w2801;
	wire w2802;
	wire w2803;
	wire w2804;
	wire w2805;
	wire w2806;
	wire w2807;
	wire w2808;
	wire w2809;
	wire w2810;
	wire w2811;
	wire w2812;
	wire w2813;
	wire w2814;
	wire w2815;
	wire w2816;
	wire w2817;
	wire w2818;
	wire w2819;
	wire w2820;
	wire w2821;
	wire w2822;
	wire w2823;
	wire w2824;
	wire w2825;
	wire w2826;
	wire w2827;
	wire w2828;
	wire w2829;
	wire w2830;
	wire w2831;
	wire w2832;
	wire w2833;
	wire w2834;
	wire w2835;
	wire w2836;
	wire w2837;
	wire w2838;
	wire w2839;
	wire w2840;
	wire w2841;
	wire w2842;
	wire w2843;
	wire w2844;
	wire w2845;
	wire w2846;
	wire w2847;
	wire w2848;
	wire w2849;
	wire w2850;
	wire w2851;
	wire w2852;
	wire w2853;
	wire w2854;
	wire w2855;
	wire w2856;
	wire w2857;
	wire w2858;
	wire w2859;
	wire w2860;
	wire w2861;
	wire w2862;
	wire w2863;
	wire w2864;
	wire w2865;
	wire w2866;
	wire w2867;
	wire w2868;
	wire w2869;
	wire w2870;
	wire w2871;
	wire w2872;
	wire w2873;
	wire w2874;
	wire w2875;
	wire w2876;
	wire w2877;
	wire w2878;
	wire w2879;
	wire w2880;
	wire w2881;
	wire w2882;
	wire w2883;
	wire w2884;
	wire w2885;
	wire w2886;
	wire w2887;
	wire w2888;
	wire w2889;
	wire w2890;
	wire w2891;
	wire w2892;
	wire w2893;
	wire w2894;
	wire w2895;
	wire w2896;
	wire w2897;
	wire w2898;
	wire w2899;
	wire w2900;
	wire w2901;
	wire w2902;
	wire w2903;
	wire w2904;
	wire w2905;
	wire w2906;
	wire w2907;
	wire w2908;
	wire w2909;
	wire w2910;
	wire w2911;
	wire w2912;
	wire w2913;
	wire w2914;
	wire w2915;
	wire w2916;
	wire w2917;
	wire w2918;
	wire w2919;
	wire w2920;
	wire w2921;
	wire w2922;
	wire w2923;
	wire w2924;
	wire w2925;
	wire w2926;
	wire w2927;
	wire w2928;
	wire w2929;
	wire w2930;
	wire w2931;
	wire w2932;
	wire w2933;
	wire w2934;
	wire w2935;
	wire w2936;
	wire w2937;
	wire w2938;
	wire w2939;
	wire w2940;
	wire w2941;
	wire w2942;
	wire w2943;
	wire w2944;
	wire w2945;
	wire w2946;
	wire w2947;
	wire w2948;
	wire w2949;
	wire w2950;
	wire S[3];
	wire w2952;
	wire w2953;
	wire S[7];
	wire S[2];
	wire w2956;
	wire w2957;
	wire w2958;
	wire w2959;
	wire w2960;
	wire w2961;
	wire S[6];
	wire S[1];
	wire S[5];
	wire S[0];
	wire S[4];
	wire w2967;
	wire w2968;
	wire w2969;
	wire w2970;
	wire w2971;
	wire w2972;
	wire w2973;
	wire w2974;
	wire w2975;
	wire w2976;
	wire w2977;
	wire w2978;
	wire w2979;
	wire w2980;
	wire w2981;
	wire w2982;
	wire w2983;
	wire w2984;
	wire w2985;
	wire w2986;
	wire w2987;
	wire w2988;
	wire w2989;
	wire w2990;
	wire w2991;
	wire w2992;
	wire w2993;
	wire w2994;
	wire w2995;
	wire w2996;
	wire w2997;
	wire w2998;
	wire w2999;
	wire w3000;
	wire w3001;
	wire w3002;
	wire w3003;
	wire w3004;
	wire w3005;
	wire w3006;
	wire w3007;
	wire w3008;
	wire w3009;
	wire w3010;
	wire w3011;
	wire w3012;
	wire w3013;
	wire w3014;
	wire w3015;
	wire w3016;
	wire w3017;
	wire w3018;
	wire w3019;
	wire w3020;
	wire w3021;
	wire w3022;
	wire w3023;
	wire w3024;
	wire w3025;
	wire w3026;
	wire w3027;
	wire w3028;
	wire w3029;
	wire w3030;
	wire w3031;
	wire w3032;
	wire w3033;
	wire w3034;
	wire w3035;
	wire w3036;
	wire w3037;
	wire w3038;
	wire w3039;
	wire w3040;
	wire w3041;
	wire w3042;
	wire w3043;
	wire w3044;
	wire w3045;
	wire w3046;
	wire w3047;
	wire w3048;
	wire w3049;
	wire w3050;
	wire w3051;
	wire w3052;
	wire w3053;
	wire w3054;
	wire w3055;
	wire w3056;
	wire w3057;
	wire w3058;
	wire w3059;
	wire w3060;
	wire w3061;
	wire w3062;
	wire w3063;
	wire w3064;
	wire w3065;
	wire w3066;
	wire w3067;
	wire w3068;
	wire w3069;
	wire w3070;
	wire w3071;
	wire w3072;
	wire w3073;
	wire w3074;
	wire w3075;
	wire w3076;
	wire w3077;
	wire w3078;
	wire w3079;
	wire w3080;
	wire w3081;
	wire w3082;
	wire w3083;
	wire w3084;
	wire w3085;
	wire w3086;
	wire w3087;
	wire w3088;
	wire w3089;
	wire w3090;
	wire w3091;
	wire w3092;
	wire w3093;
	wire w3094;
	wire w3095;
	wire w3096;
	wire w3097;
	wire w3098;
	wire w3099;
	wire w3100;
	wire w3101;
	wire w3102;
	wire w3103;
	wire w3104;
	wire w3105;
	wire w3106;
	wire w3107;
	wire w3108;
	wire w3109;
	wire w3110;
	wire w3111;
	wire w3112;
	wire w3113;
	wire w3114;
	wire w3115;
	wire w3116;
	wire w3117;
	wire w3118;
	wire w3119;
	wire w3120;
	wire w3121;
	wire w3122;
	wire w3123;
	wire w3124;
	wire w3125;
	wire w3126;
	wire w3127;
	wire w3128;
	wire w3129;
	wire w3130;
	wire w3131;
	wire w3132;
	wire w3133;
	wire w3134;
	wire w3135;
	wire w3136;
	wire w3137;
	wire w3138;
	wire w3139;
	wire w3140;
	wire w3141;
	wire w3142;
	wire w3143;
	wire w3144;
	wire w3145;
	wire w3146;
	wire w3147;
	wire w3148;
	wire w3149;
	wire w3150;
	wire w3151;
	wire w3152;
	wire w3153;
	wire w3154;
	wire w3155;
	wire w3156;
	wire w3157;
	wire w3158;
	wire w3159;
	wire w3160;
	wire w3161;
	wire w3162;
	wire w3163;
	wire w3164;
	wire w3165;
	wire w3166;
	wire w3167;
	wire w3168;
	wire w3169;
	wire w3170;
	wire w3171;
	wire w3172;
	wire w3173;
	wire w3174;
	wire w3175;
	wire w3176;
	wire w3177;
	wire w3178;
	wire w3179;
	wire w3180;
	wire w3181;
	wire w3182;
	wire w3183;
	wire w3184;
	wire w3185;
	wire w3186;
	wire w3187;
	wire w3188;
	wire w3189;
	wire w3190;
	wire w3191;
	wire w3192;
	wire w3193;
	wire w3194;
	wire w3195;
	wire w3196;
	wire w3197;
	wire w3198;
	wire w3199;
	wire w3200;
	wire w3201;
	wire w3202;
	wire w3203;
	wire w3204;
	wire w3205;
	wire w3206;
	wire w3207;
	wire w3208;
	wire w3209;
	wire w3210;
	wire w3211;
	wire w3212;
	wire w3213;
	wire w3214;
	wire w3215;
	wire w3216;
	wire w3217;
	wire w3218;
	wire w3219;
	wire w3220;
	wire w3221;
	wire w3222;
	wire w3223;
	wire w3224;
	wire w3225;
	wire w3226;
	wire w3227;
	wire w3228;
	wire w3229;
	wire w3230;
	wire w3231;
	wire w3232;
	wire w3233;
	wire w3234;
	wire w3235;
	wire w3236;
	wire w3237;
	wire w3238;
	wire w3239;
	wire w3240;
	wire w3241;
	wire w3242;
	wire w3243;
	wire w3244;
	wire w3245;
	wire w3246;
	wire w3247;
	wire w3248;
	wire w3249;
	wire w3250;
	wire w3251;
	wire w3252;
	wire w3253;
	wire w3254;
	wire w3255;
	wire w3256;
	wire w3257;
	wire w3258;
	wire w3259;
	wire w3260;
	wire w3261;
	wire w3262;
	wire w3263;
	wire w3264;
	wire w3265;
	wire w3266;
	wire w3267;
	wire w3268;
	wire w3269;
	wire w3270;
	wire w3271;
	wire w3272;
	wire w3273;
	wire w3274;
	wire w3275;
	wire w3276;
	wire w3277;
	wire w3278;
	wire w3279;
	wire w3280;
	wire w3281;
	wire w3282;
	wire w3283;
	wire w3284;
	wire w3285;
	wire w3286;
	wire w3287;
	wire w3288;
	wire w3289;
	wire w3290;
	wire w3291;
	wire w3292;
	wire w3293;
	wire w3294;
	wire w3295;
	wire w3296;
	wire w3297;
	wire w3298;
	wire w3299;
	wire w3300;
	wire w3301;
	wire w3302;
	wire w3303;
	wire w3304;
	wire w3305;
	wire w3306;
	wire w3307;
	wire w3308;
	wire w3309;
	wire w3310;
	wire w3311;
	wire w3312;
	wire w3313;
	wire w3314;
	wire w3315;
	wire w3316;
	wire w3317;
	wire w3318;
	wire w3319;
	wire w3320;
	wire w3321;
	wire w3322;
	wire w3323;
	wire w3324;
	wire w3325;
	wire w3326;
	wire w3327;
	wire w3328;
	wire w3329;
	wire w3330;
	wire w3331;
	wire w3332;
	wire w3333;
	wire w3334;
	wire w3335;
	wire w3336;
	wire w3337;
	wire w3338;
	wire w3339;
	wire w3340;
	wire w3341;
	wire w3342;
	wire w3343;
	wire w3344;
	wire w3345;
	wire w3346;
	wire w3347;
	wire w3348;
	wire w3349;
	wire w3350;
	wire w3351;
	wire w3352;
	wire w3353;
	wire w3354;
	wire w3355;
	wire w3356;
	wire w3357;
	wire w3358;
	wire w3359;
	wire w3360;
	wire w3361;
	wire w3362;
	wire w3363;
	wire w3364;
	wire w3365;
	wire w3366;
	wire w3367;
	wire w3368;
	wire w3369;
	wire w3370;
	wire w3371;
	wire w3372;
	wire w3373;
	wire w3374;
	wire w3375;
	wire w3376;
	wire w3377;
	wire w3378;
	wire w3379;
	wire w3380;
	wire w3381;
	wire w3382;
	wire w3383;
	wire w3384;
	wire w3385;
	wire w3386;
	wire w3387;
	wire w3388;
	wire w3389;
	wire w3390;
	wire w3391;
	wire w3392;
	wire w3393;
	wire w3394;
	wire w3395;
	wire w3396;
	wire w3397;
	wire w3398;
	wire w3399;
	wire w3400;
	wire w3401;
	wire w3402;
	wire w3403;
	wire w3404;
	wire w3405;
	wire w3406;
	wire w3407;
	wire w3408;
	wire w3409;
	wire w3410;
	wire w3411;
	wire w3412;
	wire w3413;
	wire w3414;
	wire w3415;
	wire w3416;
	wire w3417;
	wire w3418;
	wire w3419;
	wire w3420;
	wire w3421;
	wire w3422;
	wire w3423;
	wire w3424;
	wire w3425;
	wire w3426;
	wire w3427;
	wire w3428;
	wire w3429;
	wire w3430;
	wire w3431;
	wire w3432;
	wire w3433;
	wire w3434;
	wire w3435;
	wire w3436;
	wire w3437;
	wire w3438;
	wire w3439;
	wire w3440;
	wire w3441;
	wire w3442;
	wire w3443;
	wire w3444;
	wire w3445;
	wire w3446;
	wire w3447;
	wire w3448;
	wire w3449;
	wire w3450;
	wire w3451;
	wire w3452;
	wire w3453;
	wire w3454;
	wire w3455;
	wire w3456;
	wire w3457;
	wire w3458;
	wire w3459;
	wire w3460;
	wire w3461;
	wire w3462;
	wire w3463;
	wire w3464;
	wire w3465;
	wire w3466;
	wire w3467;
	wire w3468;
	wire w3469;
	wire w3470;
	wire w3471;
	wire w3472;
	wire w3473;
	wire w3474;
	wire w3475;
	wire w3476;
	wire w3477;
	wire w3478;
	wire w3479;
	wire w3480;
	wire w3481;
	wire w3482;
	wire w3483;
	wire w3484;
	wire w3485;
	wire w3486;
	wire w3487;
	wire w3488;
	wire w3489;
	wire w3490;
	wire w3491;
	wire w3492;
	wire w3493;
	wire w3494;
	wire w3495;
	wire w3496;
	wire w3497;
	wire w3498;
	wire w3499;
	wire w3500;
	wire w3501;
	wire w3502;
	wire w3503;
	wire w3504;
	wire w3505;
	wire w3506;
	wire w3507;
	wire w3508;
	wire w3509;
	wire w3510;
	wire w3511;
	wire w3512;
	wire w3513;
	wire w3514;
	wire w3515;
	wire w3516;
	wire w3517;
	wire w3518;
	wire w3519;
	wire w3520;
	wire w3521;
	wire w3522;
	wire w3523;
	wire w3524;
	wire w3525;
	wire w3526;
	wire w3527;
	wire w3528;
	wire w3529;
	wire w3530;
	wire w3531;
	wire w3532;
	wire w3533;
	wire w3534;
	wire w3535;
	wire w3536;
	wire w3537;
	wire w3538;
	wire w3539;
	wire w3540;
	wire w3541;
	wire w3542;
	wire w3543;
	wire w3544;
	wire w3545;
	wire w3546;
	wire w3547;
	wire w3548;
	wire w3549;
	wire w3550;
	wire w3551;
	wire w3552;
	wire w3553;
	wire w3554;
	wire w3555;
	wire w3556;
	wire w3557;
	wire w3558;
	wire w3559;
	wire w3560;
	wire w3561;
	wire w3562;
	wire w3563;
	wire w3564;
	wire w3565;
	wire w3566;
	wire w3567;
	wire w3568;
	wire w3569;
	wire w3570;
	wire w3571;
	wire w3572;
	wire w3573;
	wire w3574;
	wire w3575;
	wire w3576;
	wire w3577;
	wire w3578;
	wire w3579;
	wire w3580;
	wire w3581;
	wire w3582;
	wire w3583;
	wire w3584;
	wire w3585;
	wire w3586;
	wire w3587;
	wire w3588;
	wire w3589;
	wire w3590;
	wire w3591;
	wire w3592;
	wire w3593;
	wire w3594;
	wire w3595;
	wire w3596;
	wire w3597;
	wire w3598;
	wire w3599;
	wire w3600;
	wire w3601;
	wire w3602;
	wire w3603;
	wire w3604;
	wire w3605;
	wire w3606;
	wire w3607;
	wire w3608;
	wire w3609;
	wire w3610;
	wire w3611;
	wire w3612;
	wire w3613;
	wire w3614;
	wire w3615;
	wire w3616;
	wire w3617;
	wire w3618;
	wire w3619;
	wire w3620;
	wire w3621;
	wire w3622;
	wire w3623;
	wire w3624;
	wire w3625;
	wire w3626;
	wire w3627;
	wire w3628;
	wire w3629;
	wire w3630;
	wire w3631;
	wire w3632;
	wire w3633;
	wire w3634;
	wire w3635;
	wire w3636;
	wire w3637;
	wire w3638;
	wire w3639;
	wire w3640;
	wire w3641;
	wire w3642;
	wire w3643;
	wire w3644;
	wire w3645;
	wire w3646;
	wire w3647;
	wire w3648;
	wire w3649;
	wire w3650;
	wire w3651;
	wire w3652;
	wire w3653;
	wire w3654;
	wire w3655;
	wire w3656;
	wire w3657;
	wire w3658;
	wire w3659;
	wire w3660;
	wire w3661;
	wire w3662;
	wire w3663;
	wire w3664;
	wire w3665;
	wire w3666;
	wire w3667;
	wire w3668;
	wire w3669;
	wire w3670;
	wire w3671;
	wire w3672;
	wire w3673;
	wire w3674;
	wire w3675;
	wire w3676;
	wire w3677;
	wire w3678;
	wire w3679;
	wire w3680;
	wire w3681;
	wire w3682;
	wire w3683;
	wire w3684;
	wire w3685;
	wire w3686;
	wire w3687;
	wire w3688;
	wire w3689;
	wire w3690;
	wire w3691;
	wire w3692;
	wire w3693;
	wire w3694;
	wire w3695;
	wire w3696;
	wire w3697;
	wire w3698;
	wire w3699;
	wire w3700;
	wire w3701;
	wire w3702;
	wire w3703;
	wire w3704;
	wire w3705;
	wire w3706;
	wire w3707;
	wire w3708;
	wire w3709;
	wire w3710;
	wire w3711;
	wire w3712;
	wire w3713;
	wire w3714;
	wire w3715;
	wire w3716;
	wire w3717;
	wire w3718;
	wire w3719;
	wire w3720;
	wire w3721;
	wire w3722;
	wire w3723;
	wire w3724;
	wire w3725;
	wire w3726;
	wire w3727;
	wire w3728;
	wire w3729;
	wire w3730;
	wire w3731;
	wire w3732;
	wire w3733;
	wire w3734;
	wire w3735;
	wire w3736;
	wire w3737;
	wire w3738;
	wire w3739;
	wire w3740;
	wire w3741;
	wire w3742;
	wire w3743;
	wire w3744;
	wire w3745;
	wire w3746;
	wire w3747;
	wire w3748;
	wire w3749;
	wire w3750;
	wire w3751;
	wire w3752;
	wire w3753;
	wire w3754;
	wire w3755;
	wire w3756;
	wire w3757;
	wire w3758;
	wire w3759;
	wire w3760;
	wire w3761;
	wire w3762;
	wire w3763;
	wire w3764;
	wire w3765;
	wire w3766;
	wire w3767;
	wire w3768;
	wire w3769;
	wire w3770;
	wire w3771;
	wire w3772;
	wire w3773;
	wire w3774;
	wire w3775;
	wire w3776;
	wire w3777;
	wire w3778;
	wire w3779;
	wire w3780;
	wire w3781;
	wire w3782;
	wire w3783;
	wire w3784;
	wire w3785;
	wire con0;
	wire w3787;
	wire w3788;
	wire w3789;
	wire w3790;
	wire w3791;
	wire w3792;
	wire w3793;
	wire w3794;
	wire w3795;
	wire w3796;
	wire w3797;
	wire w3798;
	wire w3799;
	wire w3800;
	wire w3801;
	wire w3802;
	wire w3803;
	wire w3804;
	wire w3805;
	wire w3806;
	wire w3807;
	wire w3808;
	wire w3809;
	wire w3810;
	wire w3811;
	wire w3812;
	wire w3813;
	wire w3814;
	wire w3815;
	wire w3816;
	wire w3817;
	wire w3818;
	wire w3819;
	wire w3820;
	wire w3821;
	wire w3822;
	wire w3823;
	wire w3824;
	wire w3825;
	wire w3826;
	wire w3827;
	wire w3828;
	wire w3829;
	wire w3830;
	wire w3831;
	wire w3832;
	wire w3833;
	wire w3834;
	wire w3835;
	wire w3836;
	wire w3837;
	wire w3838;
	wire w3839;
	wire w3840;
	wire w3841;
	wire w3842;
	wire w3843;
	wire w3844;
	wire w3845;
	wire w3846;
	wire w3847;
	wire w3848;
	wire w3849;
	wire w3850;
	wire w3851;
	wire w3852;
	wire w3853;
	wire w3854;
	wire w3855;
	wire w3856;
	wire w3857;
	wire w3858;
	wire w3859;
	wire w3860;
	wire w3861;
	wire w3862;
	wire w3863;
	wire w3864;
	wire w3865;
	wire w3866;
	wire w3867;
	wire w3868;
	wire w3869;
	wire w3870;
	wire w3871;
	wire w3872;
	wire w3873;
	wire w3874;
	wire w3875;
	wire w3876;
	wire w3877;
	wire w3878;
	wire w3879;
	wire w3880;
	wire w3881;
	wire w3882;
	wire w3883;
	wire w3884;
	wire w3885;
	wire w3886;
	wire w3887;
	wire w3888;
	wire w3889;
	wire w3890;
	wire w3891;
	wire w3892;
	wire w3893;
	wire w3894;
	wire w3895;
	wire w3896;
	wire w3897;
	wire w3898;
	wire w3899;
	wire w3900;
	wire w3901;
	wire w3902;
	wire w3903;
	wire w3904;
	wire w3905;
	wire w3906;
	wire w3907;
	wire w3908;
	wire w3909;
	wire w3910;
	wire w3911;
	wire w3912;
	wire w3913;
	wire w3914;
	wire w3915;
	wire w3916;
	wire w3917;
	wire w3918;
	wire w3919;
	wire w3920;
	wire w3921;
	wire w3922;
	wire w3923;
	wire w3924;
	wire w3925;
	wire w3926;
	wire w3927;
	wire w3928;
	wire w3929;
	wire w3930;
	wire w3931;
	wire w3932;
	wire w3933;
	wire w3934;
	wire w3935;
	wire w3936;
	wire w3937;
	wire w3938;
	wire w3939;
	wire w3940;
	wire w3941;
	wire w3942;
	wire w3943;
	wire w3944;
	wire w3945;
	wire w3946;
	wire w3947;
	wire w3948;
	wire w3949;
	wire w3950;
	wire w3951;
	wire w3952;
	wire w3953;
	wire w3954;
	wire w3955;
	wire w3956;
	wire w3957;
	wire w3958;
	wire w3959;
	wire w3960;
	wire w3961;
	wire w3962;
	wire w3963;
	wire w3964;
	wire w3965;
	wire w3966;
	wire w3967;
	wire w3968;
	wire w3969;
	wire w3970;
	wire w3971;
	wire w3972;
	wire w3973;
	wire w3974;
	wire w3975;
	wire w3976;
	wire w3977;
	wire w3978;
	wire w3979;
	wire w3980;
	wire w3981;
	wire w3982;
	wire w3983;
	wire w3984;
	wire w3985;
	wire w3986;
	wire w3987;
	wire w3988;
	wire w3989;
	wire w3990;
	wire w3991;
	wire w3992;
	wire w3993;
	wire w3994;
	wire w3995;
	wire w3996;
	wire w3997;
	wire w3998;
	wire w3999;
	wire w4000;
	wire w4001;
	wire w4002;
	wire w4003;
	wire w4004;
	wire w4005;
	wire w4006;
	wire w4007;
	wire w4008;
	wire w4009;
	wire w4010;
	wire w4011;
	wire w4012;
	wire w4013;
	wire w4014;
	wire w4015;
	wire w4016;
	wire w4017;
	wire w4018;
	wire w4019;
	wire w4020;
	wire w4021;
	wire w4022;
	wire w4023;
	wire w4024;
	wire w4025;
	wire w4026;
	wire w4027;
	wire w4028;
	wire w4029;
	wire w4030;
	wire w4031;
	wire w4032;
	wire w4033;
	wire w4034;
	wire w4035;
	wire w4036;
	wire w4037;
	wire w4038;
	wire w4039;
	wire w4040;
	wire w4041;
	wire w4042;
	wire w4043;
	wire w4044;
	wire w4045;
	wire w4046;
	wire w4047;
	wire w4048;
	wire w4049;
	wire w4050;
	wire w4051;
	wire w4052;
	wire w4053;
	wire w4054;
	wire w4055;
	wire w4056;
	wire w4057;
	wire w4058;
	wire w4059;
	wire w4060;
	wire w4061;
	wire w4062;
	wire w4063;
	wire w4064;
	wire w4065;
	wire w4066;
	wire w4067;
	wire w4068;
	wire w4069;
	wire w4070;
	wire w4071;
	wire w4072;
	wire w4073;
	wire w4074;
	wire w4075;
	wire w4076;
	wire w4077;
	wire w4078;
	wire w4079;
	wire w4080;
	wire w4081;
	wire w4082;
	wire w4083;
	wire w4084;
	wire w4085;
	wire w4086;
	wire w4087;
	wire w4088;
	wire w4089;
	wire w4090;
	wire w4091;
	wire w4092;
	wire w4093;
	wire w4094;
	wire w4095;
	wire w4096;
	wire w4097;
	wire w4098;
	wire w4099;
	wire w4100;
	wire w4101;
	wire w4102;
	wire w4103;
	wire w4104;
	wire w4105;
	wire w4106;
	wire w4107;
	wire w4108;
	wire w4109;
	wire w4110;
	wire w4111;
	wire w4112;
	wire w4113;
	wire w4114;
	wire w4115;
	wire w4116;
	wire w4117;
	wire w4118;
	wire w4119;
	wire w4120;
	wire w4121;
	wire w4122;
	wire w4123;
	wire w4124;
	wire w4125;
	wire w4126;
	wire w4127;
	wire w4128;
	wire w4129;
	wire w4130;
	wire w4131;
	wire w4132;
	wire w4133;
	wire w4134;
	wire w4135;
	wire w4136;
	wire w4137;
	wire w4138;
	wire w4139;
	wire w4140;
	wire w4141;
	wire w4142;
	wire w4143;
	wire w4144;
	wire w4145;
	wire w4146;
	wire w4147;
	wire w4148;
	wire w4149;
	wire w4150;
	wire w4151;
	wire w4152;
	wire w4153;
	wire w4154;
	wire w4155;
	wire w4156;
	wire w4157;
	wire w4158;
	wire w4159;
	wire w4160;
	wire w4161;
	wire w4162;
	wire w4163;
	wire w4164;
	wire w4165;
	wire w4166;
	wire w4167;
	wire w4168;
	wire w4169;
	wire w4170;
	wire w4171;
	wire w4172;
	wire w4173;
	wire w4174;
	wire w4175;
	wire w4176;
	wire w4177;
	wire w4178;
	wire w4179;
	wire w4180;
	wire w4181;
	wire w4182;
	wire w4183;
	wire w4184;
	wire w4185;
	wire w4186;
	wire w4187;
	wire w4188;
	wire w4189;
	wire w4190;
	wire w4191;
	wire w4192;
	wire w4193;
	wire w4194;
	wire w4195;
	wire w4196;
	wire w4197;
	wire w4198;
	wire w4199;
	wire w4200;
	wire w4201;
	wire w4202;
	wire w4203;
	wire w4204;
	wire w4205;
	wire w4206;
	wire w4207;
	wire w4208;
	wire w4209;
	wire w4210;
	wire w4211;
	wire w4212;
	wire w4213;
	wire w4214;
	wire w4215;
	wire w4216;
	wire w4217;
	wire w4218;
	wire w4219;
	wire w4220;
	wire w4221;
	wire w4222;
	wire w4223;
	wire w4224;
	wire w4225;
	wire w4226;
	wire w4227;
	wire w4228;
	wire w4229;
	wire w4230;
	wire w4231;
	wire w4232;
	wire w4233;
	wire w4234;
	wire w4235;
	wire w4236;
	wire w4237;
	wire w4238;
	wire w4239;
	wire w4240;
	wire w4241;
	wire w4242;
	wire w4243;
	wire w4244;
	wire w4245;
	wire w4246;
	wire w4247;
	wire w4248;
	wire w4249;
	wire w4250;
	wire w4251;
	wire w4252;
	wire w4253;
	wire w4254;
	wire w4255;
	wire w4256;
	wire w4257;
	wire w4258;
	wire w4259;
	wire w4260;
	wire w4261;
	wire w4262;
	wire w4263;
	wire w4264;
	wire w4265;
	wire w4266;
	wire w4267;
	wire w4268;
	wire w4269;
	wire w4270;
	wire w4271;
	wire w4272;
	wire w4273;
	wire w4274;
	wire w4275;
	wire w4276;
	wire w4277;
	wire w4278;
	wire w4279;
	wire w4280;
	wire w4281;
	wire w4282;
	wire w4283;
	wire w4284;
	wire w4285;
	wire w4286;
	wire w4287;
	wire w4288;
	wire w4289;
	wire w4290;
	wire w4291;
	wire w4292;
	wire w4293;
	wire w4294;
	wire w4295;
	wire w4296;
	wire w4297;
	wire w4298;
	wire w4299;
	wire w4300;
	wire w4301;
	wire w4302;
	wire w4303;
	wire w4304;
	wire w4305;
	wire w4306;
	wire w4307;
	wire w4308;
	wire w4309;
	wire w4310;
	wire M68K_CPU_CLOCK;
	wire w4312;
	wire w4313;
	wire w4314;
	wire w4315;
	wire w4316;
	wire w4317;
	wire w4318;
	wire w4319;
	wire w4320;
	wire w4321;
	wire w4322;
	wire w4323;
	wire w4324;
	wire w4325;
	wire w4326;
	wire w4327;
	wire w4328;
	wire w4329;
	wire w4330;
	wire w4331;
	wire w4332;
	wire w4333;
	wire w4334;
	wire w4335;
	wire w4336;
	wire w4337;
	wire w4338;
	wire w4339;
	wire w4340;
	wire w4341;
	wire w4342;
	wire w4343;
	wire w4344;
	wire w4345;
	wire w4346;
	wire w4347;
	wire w4348;
	wire w4349;
	wire w4350;
	wire w4351;
	wire w4352;
	wire w4353;
	wire nRAS1;
	wire nCAS1;
	wire nWE1;
	wire nWE0;
	wire nOE1;
	wire AD_RD_DIR;
	wire w4360;
	wire w4361;
	wire w4362;
	wire w4363;
	wire w4364;
	wire w4365;
	wire w4366;
	wire w4367;
	wire w4368;
	wire w4369;
	wire w4370;
	wire w4371;
	wire w4372;
	wire w4373;
	wire w4374;
	wire w4375;
	wire w4376;
	wire w4377;
	wire w4378;
	wire w4379;
	wire w4380;
	wire w4381;
	wire w4382;
	wire w4383;
	wire w4384;
	wire w4385;
	wire w4386;
	wire w4387;
	wire w4388;
	wire w4389;
	wire w4390;
	wire w4391;
	wire w4392;
	wire w4393;
	wire w4394;
	wire w4395;
	wire w4396;
	wire w4397;
	wire w4398;
	wire w4399;
	wire w4400;
	wire w4401;
	wire w4402;
	wire w4403;
	wire w4404;
	wire w4405;
	wire w4406;
	wire w4407;
	wire w4408;
	wire w4409;
	wire w4410;
	wire w4411;
	wire w4412;
	wire w4413;
	wire w4414;
	wire w4415;
	wire w4416;
	wire w4417;
	wire w4418;
	wire w4419;
	wire w4420;
	wire w4421;
	wire w4422;
	wire w4423;
	wire w4424;
	wire w4425;
	wire w4426;
	wire w4427;
	wire w4428;
	wire w4429;
	wire w4430;
	wire w4431;
	wire w4432;
	wire w4433;
	wire w4434;
	wire w4435;
	wire w4436;
	wire w4437;
	wire w4438;
	wire w4439;
	wire w4440;
	wire w4441;
	wire w4442;
	wire w4443;
	wire w4444;
	wire w4445;
	wire w4446;
	wire w4447;
	wire w4448;
	wire w4449;
	wire w4450;
	wire w4451;
	wire w4452;
	wire w4453;
	wire w4454;
	wire w4455;
	wire w4456;
	wire w4457;
	wire w4458;
	wire w4459;
	wire w4460;
	wire w4461;
	wire w4462;
	wire w4463;
	wire w4464;
	wire w4465;
	wire w4466;
	wire w4467;
	wire w4468;
	wire w4469;
	wire w4470;
	wire w4471;
	wire w4472;
	wire w4473;
	wire w4474;
	wire w4475;
	wire w4476;
	wire w4477;
	wire w4478;
	wire w4479;
	wire w4480;
	wire w4481;
	wire w4482;
	wire w4483;
	wire w4484;
	wire w4485;
	wire w4486;
	wire w4487;
	wire w4488;
	wire w4489;
	wire w4490;
	wire w4491;
	wire w4492;
	wire w4493;
	wire w4494;
	wire w4495;
	wire w4496;
	wire w4497;
	wire w4498;
	wire w4499;
	wire w4500;
	wire w4501;
	wire w4502;
	wire w4503;
	wire w4504;
	wire w4505;
	wire w4506;
	wire w4507;
	wire w4508;
	wire w4509;
	wire w4510;
	wire w4511;
	wire w4512;
	wire w4513;
	wire w4514;
	wire w4515;
	wire w4516;
	wire w4517;
	wire w4518;
	wire w4519;
	wire w4520;
	wire w4521;
	wire w4522;
	wire w4523;
	wire w4524;
	wire w4525;
	wire w4526;
	wire w4527;
	wire w4528;
	wire w4529;
	wire w4530;
	wire w4531;
	wire w4532;
	wire w4533;
	wire w4534;
	wire w4535;
	wire w4536;
	wire w4537;
	wire w4538;
	wire w4539;
	wire w4540;
	wire w4541;
	wire w4542;
	wire w4543;
	wire w4544;
	wire w4545;
	wire w4546;
	wire w4547;
	wire w4548;
	wire w4549;
	wire w4550;
	wire w4551;
	wire w4552;
	wire w4553;
	wire w4554;
	wire w4555;
	wire w4556;
	wire w4557;
	wire w4558;
	wire w4559;
	wire w4560;
	wire w4561;
	wire w4562;
	wire w4563;
	wire w4564;
	wire w4565;
	wire w4566;
	wire w4567;
	wire w4568;
	wire w4569;
	wire w4570;
	wire w4571;
	wire w4572;
	wire w4573;
	wire w4574;
	wire w4575;
	wire w4576;
	wire w4577;
	wire w4578;
	wire w4579;
	wire w4580;
	wire w4581;
	wire w4582;
	wire w4583;
	wire w4584;
	wire w4585;
	wire w4586;
	wire w4587;
	wire w4588;
	wire w4589;
	wire w4590;
	wire w4591;
	wire w4592;
	wire w4593;
	wire w4594;
	wire w4595;
	wire w4596;
	wire w4597;
	wire w4598;
	wire w4599;
	wire w4600;
	wire w4601;
	wire w4602;
	wire w4603;
	wire w4604;
	wire w4605;
	wire w4606;
	wire w4607;
	wire w4608;
	wire w4609;
	wire w4610;
	wire w4611;
	wire w4612;
	wire w4613;
	wire w4614;
	wire w4615;
	wire w4616;
	wire w4617;
	wire w4618;
	wire w4619;
	wire w4620;
	wire w4621;
	wire w4622;
	wire w4623;
	wire w4624;
	wire w4625;
	wire w4626;
	wire w4627;
	wire w4628;
	wire w4629;
	wire w4630;
	wire w4631;
	wire w4632;
	wire w4633;
	wire w4634;
	wire w4635;
	wire w4636;
	wire w4637;
	wire w4638;
	wire w4639;
	wire w4640;
	wire w4641;
	wire w4642;
	wire w4643;
	wire w4644;
	wire w4645;
	wire w4646;
	wire w4647;
	wire w4648;
	wire w4649;
	wire w4650;
	wire w4651;
	wire w4652;
	wire w4653;
	wire w4654;
	wire w4655;
	wire w4656;
	wire w4657;
	wire w4658;
	wire w4659;
	wire w4660;
	wire w4661;
	wire w4662;
	wire w4663;
	wire w4664;
	wire w4665;
	wire w4666;
	wire w4667;
	wire w4668;
	wire w4669;
	wire w4670;
	wire w4671;
	wire w4672;
	wire w4673;
	wire w4674;
	wire w4675;
	wire w4676;
	wire w4677;
	wire w4678;
	wire w4679;
	wire w4680;
	wire w4681;
	wire w4682;
	wire w4683;
	wire w4684;
	wire w4685;
	wire w4686;
	wire w4687;
	wire w4688;
	wire w4689;
	wire w4690;
	wire w4691;
	wire w4692;
	wire w4693;
	wire w4694;
	wire w4695;
	wire w4696;
	wire w4697;
	wire w4698;
	wire w4699;
	wire w4700;
	wire w4701;
	wire w4702;
	wire w4703;
	wire w4704;
	wire w4705;
	wire w4706;
	wire w4707;
	wire w4708;
	wire w4709;
	wire w4710;
	wire w4711;
	wire w4712;
	wire w4713;
	wire w4714;
	wire w4715;
	wire w4716;
	wire w4717;
	wire w4718;
	wire w4719;
	wire w4720;
	wire w4721;
	wire w4722;
	wire w4723;
	wire w4724;
	wire w4725;
	wire w4726;
	wire w4727;
	wire w4728;
	wire w4729;
	wire w4730;
	wire w4731;
	wire w4732;
	wire w4733;
	wire w4734;
	wire w4735;
	wire w4736;
	wire w4737;
	wire w4738;
	wire w4739;
	wire w4740;
	wire w4741;
	wire w4742;
	wire w4743;
	wire w4744;
	wire w4745;
	wire w4746;
	wire w4747;
	wire w4748;
	wire w4749;
	wire w4750;
	wire w4751;
	wire w4752;
	wire w4753;
	wire w4754;
	wire w4755;
	wire w4756;
	wire w4757;
	wire w4758;
	wire w4759;
	wire w4760;
	wire w4761;
	wire w4762;
	wire w4763;
	wire w4764;
	wire w4765;
	wire w4766;
	wire w4767;
	wire w4768;
	wire w4769;
	wire w4770;
	wire w4771;
	wire w4772;
	wire w4773;
	wire w4774;
	wire w4775;
	wire w4776;
	wire w4777;
	wire w4778;
	wire w4779;
	wire w4780;
	wire w4781;
	wire w4782;
	wire w4783;
	wire w4784;
	wire w4785;
	wire w4786;
	wire w4787;
	wire w4788;
	wire w4789;
	wire w4790;
	wire w4791;
	wire w4792;
	wire w4793;
	wire w4794;
	wire w4795;
	wire w4796;
	wire w4797;
	wire w4798;
	wire w4799;
	wire w4800;
	wire w4801;
	wire w4802;
	wire w4803;
	wire w4804;
	wire w4805;
	wire w4806;
	wire w4807;
	wire w4808;
	wire w4809;
	wire w4810;
	wire w4811;
	wire w4812;
	wire w4813;
	wire w4814;
	wire w4815;
	wire w4816;
	wire w4817;
	wire w4818;
	wire w4819;
	wire w4820;
	wire w4821;
	wire w4822;
	wire w4823;
	wire w4824;
	wire w4825;
	wire w4826;
	wire w4827;
	wire w4828;
	wire w4829;
	wire w4830;
	wire w4831;
	wire w4832;
	wire w4833;
	wire w4834;
	wire w4835;
	wire w4836;
	wire w4837;
	wire w4838;
	wire w4839;
	wire w4840;
	wire w4841;
	wire w4842;
	wire w4843;
	wire w4844;
	wire w4845;
	wire w4846;
	wire w4847;
	wire w4848;
	wire w4849;
	wire w4850;
	wire w4851;
	wire w4852;
	wire w4853;
	wire w4854;
	wire w4855;
	wire w4856;
	wire w4857;
	wire w4858;
	wire w4859;
	wire w4860;
	wire w4861;
	wire w4862;
	wire w4863;
	wire w4864;
	wire w4865;
	wire w4866;
	wire w4867;
	wire w4868;
	wire w4869;
	wire w4870;
	wire w4871;
	wire w4872;
	wire w4873;
	wire w4874;
	wire w4875;
	wire w4876;
	wire w4877;
	wire w4878;
	wire w4879;
	wire w4880;
	wire w4881;
	wire w4882;
	wire w4883;
	wire w4884;
	wire w4885;
	wire w4886;
	wire w4887;
	wire w4888;
	wire w4889;
	wire w4890;
	wire w4891;
	wire w4892;
	wire w4893;
	wire w4894;
	wire w4895;
	wire w4896;
	wire w4897;
	wire w4898;
	wire w4899;
	wire w4900;
	wire w4901;
	wire w4902;
	wire w4903;
	wire w4904;
	wire w4905;
	wire w4906;
	wire w4907;
	wire w4908;
	wire w4909;
	wire w4910;
	wire w4911;
	wire w4912;
	wire w4913;
	wire w4914;
	wire w4915;
	wire w4916;
	wire w4917;
	wire w4918;
	wire w4919;
	wire w4920;
	wire w4921;
	wire w4922;
	wire w4923;
	wire w4924;
	wire w4925;
	wire w4926;
	wire w4927;
	wire w4928;
	wire w4929;
	wire w4930;
	wire w4931;
	wire w4932;
	wire w4933;
	wire w4934;
	wire w4935;
	wire w4936;
	wire w4937;
	wire w4938;
	wire w4939;
	wire w4940;
	wire w4941;
	wire w4942;
	wire w4943;
	wire w4944;
	wire w4945;
	wire w4946;
	wire w4947;
	wire w4948;
	wire w4949;
	wire w4950;
	wire w4951;
	wire w4952;
	wire w4953;
	wire w4954;
	wire w4955;
	wire w4956;
	wire w4957;
	wire w4958;
	wire w4959;
	wire w4960;
	wire w4961;
	wire w4962;
	wire w4963;
	wire w4964;
	wire w4965;
	wire w4966;
	wire w4967;
	wire w4968;
	wire w4969;
	wire w4970;
	wire w4971;
	wire w4972;
	wire w4973;
	wire w4974;
	wire w4975;
	wire w4976;
	wire w4977;
	wire w4978;
	wire w4979;
	wire w4980;
	wire w4981;
	wire w4982;
	wire w4983;
	wire w4984;
	wire w4985;
	wire w4986;
	wire w4987;
	wire w4988;
	wire w4989;
	wire w4990;
	wire w4991;
	wire w4992;
	wire w4993;
	wire w4994;
	wire w4995;
	wire w4996;
	wire w4997;
	wire w4998;
	wire w4999;
	wire w5000;
	wire w5001;
	wire w5002;
	wire w5003;
	wire w5004;
	wire w5005;
	wire w5006;
	wire w5007;
	wire w5008;
	wire w5009;
	wire w5010;
	wire w5011;
	wire w5012;
	wire w5013;
	wire w5014;
	wire w5015;
	wire w5016;
	wire w5017;
	wire w5018;
	wire w5019;
	wire w5020;
	wire w5021;
	wire w5022;
	wire w5023;
	wire w5024;
	wire w5025;
	wire w5026;
	wire w5027;
	wire w5028;
	wire w5029;
	wire w5030;
	wire w5031;
	wire w5032;
	wire w5033;
	wire w5034;
	wire w5035;
	wire w5036;
	wire w5037;
	wire w5038;
	wire w5039;
	wire w5040;
	wire w5041;
	wire w5042;
	wire w5043;
	wire w5044;
	wire w5045;
	wire w5046;
	wire w5047;
	wire w5048;
	wire w5049;
	wire w5050;
	wire w5051;
	wire w5052;
	wire w5053;
	wire w5054;
	wire w5055;
	wire w5056;
	wire w5057;
	wire w5058;
	wire w5059;
	wire w5060;
	wire w5061;
	wire w5062;
	wire w5063;
	wire w5064;
	wire w5065;
	wire w5066;
	wire w5067;
	wire w5068;
	wire w5069;
	wire w5070;
	wire w5071;
	wire w5072;
	wire w5073;
	wire w5074;
	wire w5075;
	wire w5076;
	wire w5077;
	wire w5078;
	wire w5079;
	wire w5080;
	wire w5081;
	wire w5082;
	wire w5083;
	wire w5084;
	wire w5085;
	wire w5086;
	wire w5087;
	wire w5088;
	wire w5089;
	wire w5090;
	wire w5091;
	wire w5092;
	wire w5093;
	wire w5094;
	wire w5095;
	wire w5096;
	wire w5097;
	wire w5098;
	wire w5099;
	wire w5100;
	wire w5101;
	wire w5102;
	wire w5103;
	wire w5104;
	wire w5105;
	wire w5106;
	wire w5107;
	wire w5108;
	wire w5109;
	wire w5110;
	wire w5111;
	wire w5112;
	wire w5113;
	wire w5114;
	wire w5115;
	wire w5116;
	wire w5117;
	wire w5118;
	wire w5119;
	wire w5120;
	wire w5121;
	wire w5122;
	wire w5123;
	wire w5124;
	wire w5125;
	wire w5126;
	wire w5127;
	wire w5128;
	wire w5129;
	wire w5130;
	wire w5131;
	wire w5132;
	wire w5133;
	wire w5134;
	wire w5135;
	wire w5136;
	wire w5137;
	wire w5138;
	wire w5139;
	wire w5140;
	wire w5141;
	wire w5142;
	wire w5143;
	wire w5144;
	wire w5145;
	wire w5146;
	wire w5147;
	wire w5148;
	wire w5149;
	wire w5150;
	wire w5151;
	wire w5152;
	wire w5153;
	wire w5154;
	wire w5155;
	wire w5156;
	wire w5157;
	wire w5158;
	wire w5159;
	wire w5160;
	wire w5161;
	wire w5162;
	wire w5163;
	wire w5164;
	wire w5165;
	wire w5166;
	wire w5167;
	wire w5168;
	wire w5169;
	wire w5170;
	wire w5171;
	wire w5172;
	wire w5173;
	wire w5174;
	wire w5175;
	wire w5176;
	wire w5177;
	wire w5178;
	wire w5179;
	wire w5180;
	wire w5181;
	wire w5182;
	wire w5183;
	wire w5184;
	wire w5185;
	wire w5186;
	wire w5187;
	wire w5188;
	wire w5189;
	wire w5190;
	wire w5191;
	wire w5192;
	wire w5193;
	wire w5194;
	wire w5195;
	wire w5196;
	wire w5197;
	wire w5198;
	wire w5199;
	wire w5200;
	wire w5201;
	wire w5202;
	wire w5203;
	wire w5204;
	wire w5205;
	wire w5206;
	wire w5207;
	wire w5208;
	wire w5209;
	wire w5210;
	wire w5211;
	wire w5212;
	wire w5213;
	wire w5214;
	wire w5215;
	wire w5216;
	wire w5217;
	wire w5218;
	wire w5219;
	wire w5220;
	wire w5221;
	wire w5222;
	wire w5223;
	wire w5224;
	wire w5225;
	wire w5226;
	wire w5227;
	wire w5228;
	wire w5229;
	wire w5230;
	wire w5231;
	wire w5232;
	wire w5233;
	wire w5234;
	wire w5235;
	wire w5236;
	wire w5237;
	wire w5238;
	wire w5239;
	wire w5240;
	wire w5241;
	wire w5242;
	wire w5243;
	wire w5244;
	wire w5245;
	wire w5246;
	wire w5247;
	wire w5248;
	wire w5249;
	wire w5250;
	wire w5251;
	wire w5252;
	wire w5253;
	wire w5254;
	wire w5255;
	wire w5256;
	wire w5257;
	wire w5258;
	wire w5259;
	wire w5260;
	wire w5261;
	wire w5262;
	wire w5263;
	wire w5264;
	wire w5265;
	wire w5266;
	wire w5267;
	wire w5268;
	wire w5269;
	wire w5270;
	wire w5271;
	wire w5272;
	wire w5273;
	wire w5274;
	wire w5275;
	wire w5276;
	wire w5277;
	wire w5278;
	wire w5279;
	wire w5280;
	wire w5281;
	wire w5282;
	wire w5283;
	wire w5284;
	wire w5285;
	wire w5286;
	wire w5287;
	wire w5288;
	wire w5289;
	wire w5290;
	wire w5291;
	wire w5292;
	wire w5293;
	wire w5294;
	wire w5295;
	wire w5296;
	wire w5297;
	wire w5298;
	wire w5299;
	wire w5300;
	wire w5301;
	wire w5302;
	wire w5303;
	wire w5304;
	wire w5305;
	wire w5306;
	wire w5307;
	wire w5308;
	wire w5309;
	wire w5310;
	wire w5311;
	wire w5312;
	wire w5313;
	wire w5314;
	wire w5315;
	wire w5316;
	wire w5317;
	wire w5318;
	wire w5319;
	wire w5320;
	wire w5321;
	wire w5322;
	wire w5323;
	wire w5324;
	wire w5325;
	wire w5326;
	wire w5327;
	wire w5328;
	wire w5329;
	wire w5330;
	wire w5331;
	wire w5332;
	wire w5333;
	wire w5334;
	wire w5335;
	wire w5336;
	wire w5337;
	wire w5338;
	wire w5339;
	wire w5340;
	wire w5341;
	wire w5342;
	wire w5343;
	wire w5344;
	wire w5345;
	wire w5346;
	wire w5347;
	wire w5348;
	wire w5349;
	wire w5350;
	wire w5351;
	wire w5352;
	wire w5353;
	wire w5354;
	wire w5355;
	wire w5356;
	wire w5357;
	wire w5358;
	wire w5359;
	wire w5360;
	wire w5361;
	wire w5362;
	wire w5363;
	wire w5364;
	wire w5365;
	wire w5366;
	wire w5367;
	wire w5368;
	wire w5369;
	wire w5370;
	wire w5371;
	wire w5372;
	wire w5373;
	wire w5374;
	wire w5375;
	wire w5376;
	wire w5377;
	wire w5378;
	wire w5379;
	wire w5380;
	wire w5381;
	wire w5382;
	wire w5383;
	wire w5384;
	wire w5385;
	wire w5386;
	wire w5387;
	wire w5388;
	wire w5389;
	wire w5390;
	wire w5391;
	wire w5392;
	wire w5393;
	wire w5394;
	wire w5395;
	wire w5396;
	wire w5397;
	wire w5398;
	wire w5399;
	wire w5400;
	wire w5401;
	wire w5402;
	wire w5403;
	wire w5404;
	wire w5405;
	wire w5406;
	wire w5407;
	wire w5408;
	wire w5409;
	wire w5410;
	wire w5411;
	wire w5412;
	wire w5413;
	wire w5414;
	wire w5415;
	wire w5416;
	wire w5417;
	wire w5418;
	wire w5419;
	wire w5420;
	wire w5421;
	wire w5422;
	wire w5423;
	wire w5424;
	wire w5425;
	wire w5426;
	wire w5427;
	wire w5428;
	wire w5429;
	wire w5430;
	wire w5431;
	wire w5432;
	wire w5433;
	wire w5434;
	wire w5435;
	wire w5436;
	wire w5437;
	wire w5438;
	wire w5439;
	wire w5440;
	wire w5441;
	wire w5442;
	wire w5443;
	wire w5444;
	wire w5445;
	wire w5446;
	wire w5447;
	wire w5448;
	wire w5449;
	wire w5450;
	wire w5451;
	wire w5452;
	wire w5453;
	wire w5454;
	wire w5455;
	wire w5456;
	wire w5457;
	wire w5458;
	wire w5459;
	wire w5460;
	wire w5461;
	wire w5462;
	wire w5463;
	wire w5464;
	wire w5465;
	wire w5466;
	wire w5467;
	wire w5468;
	wire w5469;
	wire w5470;
	wire w5471;
	wire w5472;
	wire w5473;
	wire w5474;
	wire w5475;
	wire w5476;
	wire w5477;
	wire w5478;
	wire w5479;
	wire w5480;
	wire w5481;
	wire w5482;
	wire w5483;
	wire w5484;
	wire w5485;
	wire w5486;
	wire w5487;
	wire w5488;
	wire w5489;
	wire w5490;
	wire w5491;
	wire w5492;
	wire w5493;
	wire w5494;
	wire w5495;
	wire w5496;
	wire w5497;
	wire w5498;
	wire w5499;
	wire w5500;
	wire w5501;
	wire w5502;
	wire w5503;
	wire w5504;
	wire w5505;
	wire w5506;
	wire w5507;
	wire w5508;
	wire w5509;
	wire w5510;
	wire w5511;
	wire w5512;
	wire w5513;
	wire w5514;
	wire w5515;
	wire w5516;
	wire w5517;
	wire w5518;
	wire w5519;
	wire w5520;
	wire w5521;
	wire w5522;
	wire w5523;
	wire w5524;
	wire w5525;
	wire w5526;
	wire w5527;
	wire w5528;
	wire w5529;
	wire w5530;
	wire w5531;
	wire w5532;
	wire w5533;
	wire w5534;
	wire w5535;
	wire w5536;
	wire w5537;
	wire w5538;
	wire w5539;
	wire w5540;
	wire w5541;
	wire w5542;
	wire w5543;
	wire w5544;
	wire w5545;
	wire w5546;
	wire w5547;
	wire w5548;
	wire w5549;
	wire w5550;
	wire w5551;
	wire w5552;
	wire w5553;
	wire w5554;
	wire w5555;
	wire w5556;
	wire w5557;
	wire w5558;
	wire w5559;
	wire w5560;
	wire w5561;
	wire w5562;
	wire w5563;
	wire w5564;
	wire w5565;
	wire w5566;
	wire w5567;
	wire w5568;
	wire w5569;
	wire w5570;
	wire w5571;
	wire w5572;
	wire w5573;
	wire w5574;
	wire w5575;
	wire w5576;
	wire w5577;
	wire w5578;
	wire w5579;
	wire w5580;
	wire w5581;
	wire w5582;
	wire w5583;
	wire w5584;
	wire w5585;
	wire w5586;
	wire w5587;
	wire w5588;
	wire w5589;
	wire w5590;
	wire w5591;
	wire w5592;
	wire w5593;
	wire w5594;
	wire w5595;
	wire w5596;
	wire w5597;
	wire w5598;
	wire w5599;
	wire w5600;
	wire w5601;
	wire w5602;
	wire w5603;
	wire w5604;
	wire w5605;
	wire w5606;
	wire w5607;
	wire w5608;
	wire w5609;
	wire w5610;
	wire w5611;
	wire w5612;
	wire w5613;
	wire w5614;
	wire w5615;
	wire w5616;
	wire w5617;
	wire w5618;
	wire w5619;
	wire w5620;
	wire w5621;
	wire w5622;
	wire w5623;
	wire w5624;
	wire w5625;
	wire w5626;
	wire w5627;
	wire w5628;
	wire w5629;
	wire w5630;
	wire w5631;
	wire w5632;
	wire w5633;
	wire w5634;
	wire w5635;
	wire w5636;
	wire w5637;
	wire w5638;
	wire w5639;
	wire w5640;
	wire w5641;
	wire w5642;
	wire w5643;
	wire w5644;
	wire w5645;
	wire w5646;
	wire w5647;
	wire w5648;
	wire w5649;
	wire w5650;
	wire w5651;
	wire w5652;
	wire w5653;
	wire w5654;
	wire w5655;
	wire w5656;
	wire w5657;
	wire w5658;
	wire w5659;
	wire w5660;
	wire w5661;
	wire w5662;
	wire w5663;
	wire w5664;
	wire w5665;
	wire w5666;
	wire w5667;
	wire w5668;
	wire w5669;
	wire w5670;
	wire w5671;
	wire w5672;
	wire w5673;
	wire w5674;
	wire w5675;
	wire w5676;
	wire w5677;
	wire w5678;
	wire w5679;
	wire w5680;
	wire w5681;
	wire w5682;
	wire w5683;
	wire w5684;
	wire w5685;
	wire w5686;
	wire w5687;
	wire w5688;
	wire w5689;
	wire w5690;
	wire w5691;
	wire w5692;
	wire w5693;
	wire w5694;
	wire w5695;
	wire w5696;
	wire w5697;
	wire w5698;
	wire w5699;
	wire w5700;
	wire w5701;
	wire w5702;
	wire w5703;
	wire w5704;
	wire w5705;
	wire w5706;
	wire w5707;
	wire w5708;
	wire w5709;
	wire w5710;
	wire w5711;
	wire w5712;
	wire w5713;
	wire w5714;
	wire w5715;
	wire w5716;
	wire w5717;
	wire w5718;
	wire w5719;
	wire w5720;
	wire w5721;
	wire w5722;
	wire w5723;
	wire w5724;
	wire w5725;
	wire w5726;
	wire w5727;
	wire w5728;
	wire w5729;
	wire w5730;
	wire w5731;
	wire w5732;
	wire w5733;
	wire w5734;
	wire w5735;
	wire w5736;
	wire w5737;
	wire w5738;
	wire w5739;
	wire w5740;
	wire w5741;
	wire w5742;
	wire w5743;
	wire w5744;
	wire w5745;
	wire w5746;
	wire w5747;
	wire w5748;
	wire w5749;
	wire w5750;
	wire w5751;
	wire w5752;
	wire w5753;
	wire w5754;
	wire w5755;
	wire w5756;
	wire w5757;
	wire w5758;
	wire w5759;
	wire w5760;
	wire w5761;
	wire w5762;
	wire w5763;
	wire w5764;
	wire w5765;
	wire w5766;
	wire w5767;
	wire w5768;
	wire w5769;
	wire w5770;
	wire w5771;
	wire w5772;
	wire w5773;
	wire w5774;
	wire w5775;
	wire w5776;
	wire w5777;
	wire w5778;
	wire w5779;
	wire w5780;
	wire w5781;
	wire w5782;
	wire w5783;
	wire w5784;
	wire w5785;
	wire w5786;
	wire w5787;
	wire w5788;
	wire w5789;
	wire w5790;
	wire w5791;
	wire w5792;
	wire w5793;
	wire w5794;
	wire w5795;
	wire w5796;
	wire w5797;
	wire w5798;
	wire w5799;
	wire w5800;
	wire w5801;
	wire w5802;
	wire w5803;
	wire w5804;
	wire w5805;
	wire w5806;
	wire w5807;
	wire w5808;
	wire w5809;
	wire w5810;
	wire w5811;
	wire w5812;
	wire w5813;
	wire w5814;
	wire w5815;
	wire w5816;
	wire w5817;
	wire w5818;
	wire w5819;
	wire w5820;
	wire w5821;
	wire w5822;
	wire w5823;
	wire w5824;
	wire w5825;
	wire w5826;
	wire w5827;
	wire w5828;
	wire w5829;
	wire w5830;
	wire w5831;
	wire w5832;
	wire w5833;
	wire w5834;
	wire w5835;
	wire w5836;
	wire w5837;
	wire w5838;
	wire w5839;
	wire w5840;
	wire w5841;
	wire w5842;
	wire w5843;
	wire w5844;
	wire w5845;
	wire w5846;
	wire w5847;
	wire w5848;
	wire w5849;
	wire w5850;
	wire w5851;
	wire w5852;
	wire w5853;
	wire w5854;
	wire w5855;
	wire w5856;
	wire w5857;
	wire w5858;
	wire w5859;
	wire w5860;
	wire w5861;
	wire w5862;
	wire w5863;
	wire w5864;
	wire w5865;
	wire w5866;
	wire w5867;
	wire w5868;
	wire w5869;
	wire w5870;
	wire w5871;
	wire w5872;
	wire w5873;
	wire w5874;
	wire w5875;
	wire w5876;
	wire w5877;
	wire w5878;
	wire w5879;
	wire w5880;
	wire w5881;
	wire w5882;
	wire w5883;
	wire w5884;
	wire w5885;
	wire w5886;
	wire w5887;
	wire w5888;
	wire w5889;
	wire w5890;
	wire w5891;
	wire w5892;
	wire w5893;
	wire w5894;
	wire w5895;
	wire w5896;
	wire w5897;
	wire w5898;
	wire w5899;
	wire w5900;
	wire w5901;
	wire w5902;
	wire w5903;
	wire w5904;
	wire w5905;
	wire w5906;
	wire w5907;
	wire w5908;
	wire w5909;
	wire w5910;
	wire w5911;
	wire w5912;
	wire w5913;
	wire w5914;
	wire w5915;
	wire w5916;
	wire w5917;
	wire w5918;
	wire w5919;
	wire w5920;
	wire w5921;
	wire w5922;
	wire w5923;
	wire w5924;
	wire w5925;
	wire w5926;
	wire w5927;
	wire w5928;
	wire w5929;
	wire w5930;
	wire w5931;
	wire w5932;
	wire w5933;
	wire w5934;
	wire w5935;
	wire w5936;
	wire w5937;
	wire w5938;
	wire w5939;
	wire w5940;
	wire w5941;
	wire w5942;
	wire w5943;
	wire w5944;
	wire w5945;
	wire w5946;
	wire w5947;
	wire w5948;
	wire w5949;
	wire w5950;
	wire w5951;
	wire w5952;
	wire w5953;
	wire w5954;
	wire w5955;
	wire w5956;
	wire w5957;
	wire w5958;
	wire w5959;
	wire w5960;
	wire w5961;
	wire w5962;
	wire w5963;
	wire w5964;
	wire w5965;
	wire w5966;
	wire w5967;
	wire w5968;
	wire w5969;
	wire w5970;
	wire w5971;
	wire w5972;
	wire w5973;
	wire w5974;
	wire w5975;
	wire w5976;
	wire w5977;
	wire w5978;
	wire w5979;
	wire w5980;
	wire w5981;
	wire w5982;
	wire w5983;
	wire w5984;
	wire w5985;
	wire w5986;
	wire w5987;
	wire w5988;
	wire w5989;
	wire w5990;
	wire w5991;
	wire w5992;
	wire w5993;
	wire w5994;
	wire w5995;
	wire w5996;
	wire w5997;
	wire w5998;
	wire w5999;
	wire w6000;
	wire w6001;
	wire w6002;
	wire w6003;
	wire w6004;
	wire w6005;
	wire w6006;
	wire w6007;
	wire w6008;
	wire w6009;
	wire w6010;
	wire w6011;
	wire w6012;
	wire w6013;
	wire w6014;
	wire w6015;
	wire w6016;
	wire w6017;
	wire w6018;
	wire w6019;
	wire w6020;
	wire w6021;
	wire w6022;
	wire w6023;
	wire w6024;
	wire w6025;
	wire w6026;
	wire w6027;
	wire w6028;
	wire w6029;
	wire w6030;
	wire w6031;
	wire w6032;
	wire w6033;
	wire w6034;
	wire w6035;
	wire w6036;
	wire w6037;
	wire w6038;
	wire w6039;
	wire w6040;
	wire w6041;
	wire w6042;
	wire w6043;
	wire w6044;
	wire w6045;
	wire w6046;
	wire w6047;
	wire w6048;
	wire w6049;
	wire w6050;
	wire w6051;
	wire w6052;
	wire w6053;
	wire w6054;
	wire w6055;
	wire w6056;
	wire w6057;
	wire w6058;
	wire w6059;
	wire w6060;
	wire w6061;
	wire w6062;
	wire w6063;
	wire w6064;
	wire w6065;
	wire w6066;
	wire w6067;
	wire w6068;
	wire w6069;
	wire w6070;
	wire w6071;
	wire w6072;
	wire w6073;
	wire w6074;
	wire w6075;
	wire w6076;
	wire w6077;
	wire w6078;
	wire w6079;
	wire w6080;
	wire w6081;
	wire w6082;
	wire w6083;
	wire w6084;
	wire w6085;
	wire w6086;
	wire w6087;
	wire w6088;
	wire w6089;
	wire w6090;
	wire w6091;
	wire w6092;
	wire w6093;
	wire w6094;
	wire w6095;
	wire w6096;
	wire w6097;
	wire w6098;
	wire w6099;
	wire w6100;
	wire w6101;
	wire w6102;
	wire w6103;
	wire w6104;
	wire w6105;
	wire w6106;
	wire w6107;
	wire w6108;
	wire w6109;
	wire w6110;
	wire w6111;
	wire w6112;
	wire w6113;
	wire w6114;
	wire w6115;
	wire w6116;
	wire w6117;
	wire w6118;
	wire w6119;
	wire w6120;
	wire w6121;
	wire w6122;
	wire w6123;
	wire w6124;
	wire w6125;
	wire w6126;
	wire w6127;
	wire w6128;
	wire w6129;
	wire w6130;
	wire w6131;
	wire w6132;
	wire w6133;
	wire w6134;
	wire w6135;
	wire w6136;
	wire w6137;
	wire w6138;
	wire w6139;
	wire w6140;
	wire w6141;
	wire w6142;
	wire w6143;
	wire w6144;
	wire w6145;
	wire w6146;
	wire w6147;
	wire w6148;
	wire w6149;
	wire w6150;
	wire w6151;
	wire w6152;
	wire w6153;
	wire w6154;
	wire w6155;
	wire w6156;
	wire w6157;
	wire w6158;
	wire w6159;
	wire w6160;
	wire w6161;
	wire w6162;
	wire w6163;
	wire w6164;
	wire w6165;
	wire w6166;
	wire w6167;
	wire w6168;
	wire w6169;
	wire w6170;
	wire w6171;
	wire w6172;
	wire w6173;
	wire w6174;
	wire w6175;
	wire w6176;
	wire w6177;
	wire w6178;
	wire w6179;
	wire w6180;
	wire w6181;
	wire w6182;
	wire w6183;
	wire w6184;
	wire w6185;
	wire w6186;
	wire w6187;
	wire w6188;
	wire w6189;
	wire w6190;
	wire w6191;
	wire w6192;
	wire w6193;
	wire w6194;
	wire w6195;
	wire w6196;
	wire w6197;
	wire w6198;
	wire w6199;
	wire w6200;
	wire w6201;
	wire w6202;
	wire w6203;
	wire w6204;
	wire w6205;
	wire w6206;
	wire w6207;
	wire w6208;
	wire w6209;
	wire w6210;
	wire w6211;
	wire w6212;
	wire w6213;
	wire w6214;
	wire w6215;
	wire w6216;
	wire w6217;
	wire w6218;
	wire w6219;
	wire w6220;
	wire w6221;
	wire w6222;
	wire w6223;
	wire w6224;
	wire w6225;
	wire w6226;
	wire w6227;
	wire w6228;
	wire w6229;
	wire w6230;
	wire w6231;
	wire w6232;
	wire w6233;
	wire w6234;
	wire w6235;
	wire w6236;
	wire w6237;
	wire w6238;
	wire w6239;
	wire w6240;
	wire w6241;
	wire w6242;
	wire w6243;
	wire w6244;
	wire w6245;
	wire w6246;
	wire w6247;
	wire w6248;
	wire w6249;
	wire w6250;
	wire w6251;
	wire w6252;
	wire w6253;
	wire w6254;
	wire w6255;
	wire w6256;
	wire w6257;
	wire w6258;
	wire w6259;
	wire w6260;
	wire w6261;
	wire w6262;
	wire w6263;
	wire w6264;
	wire w6265;
	wire w6266;
	wire w6267;
	wire w6268;
	wire w6269;
	wire w6270;
	wire w6271;
	wire w6272;
	wire w6273;
	wire w6274;
	wire w6275;
	wire w6276;
	wire w6277;
	wire w6278;
	wire w6279;
	wire w6280;
	wire w6281;
	wire w6282;
	wire w6283;
	wire w6284;
	wire w6285;
	wire w6286;
	wire w6287;
	wire w6288;
	wire w6289;
	wire w6290;
	wire w6291;
	wire w6292;
	wire w6293;
	wire w6294;
	wire w6295;
	wire w6296;
	wire w6297;
	wire w6298;
	wire w6299;
	wire w6300;
	wire w6301;
	wire w6302;
	wire w6303;
	wire w6304;
	wire w6305;
	wire w6306;
	wire w6307;
	wire w6308;
	wire w6309;
	wire w6310;
	wire w6311;
	wire w6312;
	wire w6313;
	wire w6314;
	wire w6315;
	wire w6316;
	wire w6317;
	wire w6318;
	wire w6319;
	wire w6320;
	wire w6321;
	wire w6322;
	wire w6323;
	wire w6324;
	wire w6325;
	wire w6326;
	wire w6327;
	wire w6328;
	wire w6329;
	wire w6330;
	wire w6331;
	wire w6332;
	wire w6333;
	wire w6334;
	wire w6335;
	wire w6336;
	wire w6337;
	wire w6338;
	wire w6339;
	wire w6340;
	wire w6341;
	wire w6342;
	wire w6343;
	wire w6344;
	wire w6345;
	wire w6346;
	wire w6347;
	wire w6348;
	wire w6349;
	wire w6350;
	wire w6351;
	wire w6352;
	wire w6353;
	wire w6354;
	wire w6355;
	wire w6356;
	wire w6357;
	wire w6358;
	wire w6359;
	wire w6360;
	wire w6361;
	wire w6362;
	wire w6363;
	wire w6364;
	wire w6365;
	wire w6366;
	wire w6367;
	wire w6368;
	wire w6369;
	wire w6370;
	wire w6371;
	wire w6372;
	wire w6373;
	wire w6374;
	wire w6375;
	wire w6376;
	wire w6377;
	wire w6378;
	wire w6379;
	wire w6380;
	wire w6381;
	wire w6382;
	wire w6383;
	wire w6384;
	wire w6385;
	wire w6386;
	wire w6387;
	wire w6388;
	wire w6389;
	wire w6390;
	wire w6391;
	wire w6392;
	wire w6393;
	wire w6394;
	wire w6395;
	wire w6396;
	wire w6397;
	wire w6398;
	wire w6399;
	wire w6400;
	wire w6401;
	wire w6402;
	wire w6403;
	wire w6404;
	wire w6405;
	wire w6406;
	wire w6407;
	wire w6408;
	wire w6409;
	wire w6410;
	wire w6411;
	wire w6412;
	wire w6413;
	wire w6414;
	wire w6415;
	wire w6416;
	wire w6417;
	wire w6418;
	wire w6419;
	wire w6420;
	wire w6421;
	wire w6422;
	wire w6423;
	wire w6424;
	wire w6425;
	wire w6426;
	wire w6427;
	wire w6428;
	wire w6429;
	wire w6430;
	wire w6431;
	wire w6432;
	wire w6433;
	wire w6434;
	wire w6435;
	wire w6436;
	wire w6437;
	wire w6438;
	wire w6439;
	wire w6440;
	wire w6441;
	wire w6442;
	wire w6443;
	wire w6444;
	wire w6445;
	wire w6446;
	wire w6447;
	wire w6448;
	wire w6449;
	wire w6450;
	wire w6451;
	wire w6452;
	wire w6453;
	wire w6454;
	wire w6455;
	wire w6456;
	wire w6457;
	wire w6458;
	wire w6459;
	wire w6460;
	wire w6461;
	wire w6462;
	wire w6463;
	wire w6464;
	wire w6465;
	wire w6466;
	wire w6467;
	wire w6468;
	wire w6469;
	wire w6470;
	wire w6471;
	wire w6472;
	wire w6473;
	wire w6474;
	wire w6475;
	wire w6476;
	wire w6477;
	wire w6478;
	wire w6479;
	wire w6480;
	wire w6481;
	wire w6482;
	wire w6483;
	wire w6484;
	wire w6485;
	wire w6486;
	wire w6487;
	wire w6488;
	wire w6489;
	wire w6490;
	wire w6491;
	wire w6492;
	wire w6493;
	wire w6494;
	wire w6495;
	wire w6496;
	wire w6497;
	wire w6498;
	wire w6499;
	wire w6500;
	wire w6501;
	wire w6502;
	wire w6503;
	wire w6504;
	wire w6505;
	wire w6506;
	wire w6507;
	wire w6508;
	wire w6509;
	wire w6510;
	wire w6511;
	wire w6512;
	wire w6513;
	wire w6514;
	wire w6515;
	wire w6516;
	wire w6517;
	wire w6518;
	wire w6519;
	wire w6520;
	wire w6521;
	wire w6522;
	wire w6523;
	wire w6524;
	wire w6525;
	wire w6526;
	wire w6527;
	wire w6528;
	wire w6529;
	wire w6530;
	wire w6531;
	wire w6532;
	wire w6533;
	wire w6534;
	wire w6535;
	wire w6536;
	wire w6537;
	wire w6538;
	wire w6539;
	wire w6540;
	wire w6541;
	wire w6542;
	wire w6543;
	wire w6544;
	wire w6545;
	wire w6546;
	wire w6547;
	wire w6548;
	wire w6549;
	wire w6550;
	wire w6551;
	wire w6552;
	wire w6553;
	wire w6554;
	wire w6555;
	wire w6556;
	wire w6557;
	wire w6558;
	wire w6559;
	wire w6560;
	wire w6561;
	wire w6562;
	wire w6563;
	wire w6564;
	wire w6565;
	wire w6566;
	wire w6567;
	wire w6568;
	wire w6569;
	wire w6570;
	wire w6571;
	wire w6572;
	wire w6573;
	wire w6574;
	wire w6575;
	wire w6576;
	wire w6577;
	wire w6578;
	wire w6579;
	wire w6580;
	wire w6581;
	wire w6582;
	wire w6583;
	wire w6584;
	wire w6585;
	wire w6586;
	wire w6587;
	wire w6588;
	wire w6589;
	wire w6590;
	wire w6591;
	wire w6592;
	wire w6593;
	wire w6594;
	wire w6595;
	wire w6596;
	wire w6597;
	wire w6598;
	wire w6599;
	wire w6600;
	wire w6601;
	wire w6602;
	wire w6603;
	wire w6604;
	wire w6605;
	wire w6606;
	wire w6607;
	wire w6608;
	wire w6609;
	wire w6610;
	wire w6611;
	wire w6612;
	wire w6613;
	wire w6614;
	wire w6615;
	wire w6616;
	wire w6617;
	wire w6618;
	wire w6619;
	wire w6620;

	assign CH0_EN = w1942;
	assign CH0VOL[0] = w1945;
	assign CH0VOL[1] = w1946;
	assign CH1_EN = w1943;
	assign CH1VOL[0] = w2005;
	assign CH1VOL[1] = w2006;
	assign CH2_EN = w1940;
	assign CH2VOL[0] = w2025;
	assign CH2VOL[1] = w2024;
	assign CH3_EN = w1941;
	assign CH3VOL[0] = w2047;
	assign CH3VOL[1] = w2046;
	assign PSGDAC0[0] = w1947;
	assign PSGDAC0[1] = w1948;
	assign PSGDAC0[2] = w1949;
	assign PSGDAC0[3] = w1950;
	assign PSGDAC0[4] = w1951;
	assign PSGDAC0[5] = w1952;
	assign PSGDAC0[6] = w1953;
	assign PSGDAC0[7] = w1954;
	assign PSGDAC1[0] = w2007;
	assign PSGDAC1[1] = w2008;
	assign PSGDAC1[2] = w2009;
	assign PSGDAC1[3] = w2010;
	assign PSGDAC1[4] = w2011;
	assign PSGDAC1[5] = w2012;
	assign PSGDAC1[6] = w2013;
	assign PSGDAC1[7] = w2014;
	assign PSGDAC2[0] = w2036;
	assign PSGDAC2[1] = w2037;
	assign PSGDAC2[2] = w2038;
	assign PSGDAC2[3] = w2039;
	assign PSGDAC2[4] = w2040;
	assign PSGDAC2[5] = w2041;
	assign PSGDAC2[6] = w2042;
	assign PSGDAC2[7] = w2043;
	assign PSGDAC3[0] = w2045;
	assign PSGDAC3[1] = w2044;
	assign PSGDAC3[2] = w2052;
	assign PSGDAC3[3] = w2051;
	assign PSGDAC3[4] = w2050;
	assign PSGDAC3[5] = w2049;
	assign PSGDAC3[6] = w2048;
	assign PSGDAC3[7] = w2053;
	assign w1166 = CAi[22];
	assign CAo[22] = w1317;
	assign CA[19] = CA[19];
	assign DTACK_OUT = w1021;
	assign Z80_INT = w1022;
	assign RA[7] = w1072;
	assign RA[6] = w1084;
	assign RA[5] = w1073;
	assign RA[4] = w1074;
	assign RA[2] = w1076;
	assign RA[1] = w1083;
	assign RA[0] = w1077;
	assign nRAS0 = w1294;
	assign RA[3] = w1075;
	assign nCAS0 = w1363;
	assign nOE0 = w1354;
	assign nLWR = w1355;
	assign nUWR = w1270;
	assign w1342 = DTACK_IN;
	assign w967 = RnW;
	assign w1337 = nLDS;
	assign w1328 = nUDS;
	assign w1215 = nAS;
	assign w1326 = nM1;
	assign w1327 = nWR;
	assign w1324 = nRD;
	assign w1325 = nIORQ;
	assign nILP2 = w1330;
	assign nILP1 = w1329;
	assign w1197 = nINTAK;
	assign w1323 = nMREQ;
	assign w1198 = nBG;
	assign BGACK_OUT = w1213;
	assign w1341 = BGACK_IN;
	assign nBR = w1383;
	assign VSYNC = w1642;
	assign nCSYNC = w1928;
	assign w1636 = nCSYNC_IN;
	assign nHSYNC = w1699;
	assign w1898 = nHSYNC_IN;
	assign DB[15] = DB[15];
	assign DB[14] = DB[14];
	assign DB[13] = DB[13];
	assign DB[12] = DB[12];
	assign DB[11] = DB[11];
	assign DB[10] = DB[10];
	assign DB[9] = DB[9];
	assign DB[8] = DB[8];
	assign DB[7] = DB[7];
	assign DB[6] = DB[6];
	assign DB[5] = DB[5];
	assign DB[4] = DB[4];
	assign DB[3] = DB[3];
	assign DB[2] = DB[2];
	assign DB[1] = DB[1];
	assign DB[0] = DB[0];
	assign CA[0] = CA[0];
	assign CA[1] = CA[1];
	assign CA[2] = CA[2];
	assign CA[3] = CA[3];
	assign CA[4] = CA[4];
	assign CA[5] = CA[5];
	assign CA[6] = CA[6];
	assign CA[7] = CA[7];
	assign CA[8] = CA[8];
	assign CA[9] = CA[9];
	assign CA[10] = CA[10];
	assign CA[11] = CA[11];
	assign CA[12] = CA[12];
	assign CA[13] = CA[13];
	assign CA[14] = CA[14];
	assign CA[15] = CA[15];
	assign CA[17] = CA[17];
	assign CA[18] = CA[18];
	assign CA[20] = CA[20];
	assign CA[21] = CA[21];
	assign R_DAC[0] = w2849;
	assign R_DAC[1] = w2814;
	assign R_DAC[2] = w2848;
	assign R_DAC[3] = w2813;
	assign R_DAC[4] = w2847;
	assign R_DAC[5] = w2846;
	assign R_DAC[6] = w2845;
	assign R_DAC[7] = w2844;
	assign R_DAC[8] = w2810;
	assign G_DAC[0] = w2842;
	assign G_DAC[1] = w2841;
	assign G_DAC[2] = w2804;
	assign G_DAC[3] = w2803;
	assign G_DAC[4] = w2802;
	assign G_DAC[5] = w2801;
	assign G_DAC[6] = w2800;
	assign G_DAC[7] = w2799;
	assign G_DAC[8] = w2798;
	assign R_DAC[9] = w2811;
	assign R_DAC[10] = w2808;
	assign R_DAC[11] = w2812;
	assign R_DAC[12] = w2807;
	assign R_DAC[13] = w2809;
	assign R_DAC[14] = w2806;
	assign R_DAC[15] = w2805;
	assign R_DAC[16] = w2843;
	assign B_DAC[0] = w2790;
	assign B_DAC[1] = w2840;
	assign B_DAC[2] = w2836;
	assign B_DAC[3] = w2837;
	assign B_DAC[4] = w2838;
	assign B_DAC[5] = w2835;
	assign B_DAC[6] = w2839;
	assign B_DAC[7] = w2895;
	assign B_DAC[8] = w2791;
	assign G_DAC[9] = w2792;
	assign G_DAC[10] = w2797;
	assign G_DAC[11] = w2796;
	assign G_DAC[12] = w2893;
	assign G_DAC[13] = w2795;
	assign G_DAC[14] = w2794;
	assign G_DAC[15] = w2793;
	assign G_DAC[16] = w2894;
	assign B_DAC[9] = w2788;
	assign B_DAC[10] = w2789;
	assign B_DAC[11] = w2834;
	assign B_DAC[12] = w2833;
	assign B_DAC[13] = w2832;
	assign B_DAC[14] = w2831;
	assign B_DAC[15] = w2829;
	assign B_DAC[16] = w2830;
	assign nOE1 = nOE1;
	assign nWE0 = nWE0;
	assign nWE1 = nWE1;
	assign nCAS1 = nCAS1;
	assign nRAS1 = nRAS1;
	assign AD_RD_DIR = AD_RD_DIR;
	assign nYS = nYS;
	assign nSC = w2513;
	assign nSE0_1 = w2408;
	assign ADo[7] = w2491;
	assign ADo[6] = w2603;
	assign ADo[5] = w2592;
	assign ADo[4] = w2605;
	assign ADo[3] = w2597;
	assign ADo[2] = w2595;
	assign ADo[1] = w2604;
	assign ADo[0] = w2593;
	assign RDo[6] = w2551;
	assign RDo[5] = w2570;
	assign RDo[4] = w2556;
	assign RDo[3] = w2555;
	assign RDo[2] = w2571;
	assign RDo[1] = w2594;
	assign RDo[0] = w2415;
	assign w2454 = RDi[6];
	assign w2371 = RDi[7];
	assign w2383 = RDi[4];
	assign w2582 = RDi[5];
	assign w2448 = RDi[2];
	assign w2456 = RDi[3];
	assign w2572 = RDi[0];
	assign w2490 = RDi[1];
	assign w2455 = ADi[6];
	assign w2554 = ADi[7];
	assign w2401 = ADi[4];
	assign w2609 = ADi[5];
	assign w2443 = ADi[2];
	assign w2447 = ADi[3];
	assign w2416 = ADi[0];
	assign w2435 = ADi[1];
	assign RDo[7] = w2553;
	assign w5099 = SD[7];
	assign w5100 = SD[6];
	assign w6422 = SD[5];
	assign w6424 = SD[4];
	assign w5101 = SD[3];
	assign w5098 = SD[2];
	assign w6423 = SD[1];
	assign w5097 = SD[0];
	assign CLK1 = M68K_CPU_CLOCK;
	assign CLK0 = w1357;
	assign w4332 = EDCLKi;
	assign EDCLKo = EDCLK_O;
	assign w4310 = MCLK;
	assign SUB_CLK = w4299;
	assign w4350 = nRES_PAD;
	assign w1384 = M68kCLKi;
	assign EDCLKd = w1440;
	assign CA_PAD_DIR = w2368;
	assign DB_PAD_DIR = w2369;
	assign SEL0_M3 = SEL0_M3;
	assign w6428 = nPAL;
	assign w428 = nHL;
	assign SPA_Bo = w2723;
	assign w2700 = SPA_Bi;

	// Instances

	vdp_slatch g1 (.nQ(w351), .D(VPOS[7]), .C(w1511), .nC(w1512) );
	vdp_slatch g2 (.nQ(w1474), .D(HPOS[8]), .C(w372), .nC(w373) );
	vdp_slatch g3 (.nQ(w356), .D(w298), .C(w1413), .nC(w374) );
	vdp_slatch g4 (.D(w299), .C(w1509), .nC(w1510), .nQ(w6530) );
	vdp_slatch g5 (.nQ(w357), .D(w358), .C(w1507), .nC(w1508) );
	vdp_slatch g6 (.nQ(w301), .D(w302), .C(w1505), .nC(w1506) );
	vdp_slatch g7 (.nQ(w359), .D(w358), .C(w375), .nC(w376) );
	vdp_slatch g8 (.nQ(w362), .D(w302), .C(w377), .nC(w378) );
	vdp_slatch g9 (.nQ(w360), .D(w358), .C(w417), .nC(w1410) );
	vdp_slatch g10 (.nQ(w363), .D(w302), .C(w1409), .nC(w383) );
	vdp_slatch g11 (.nQ(w361), .D(w358), .C(w381), .nC(w380) );
	vdp_slatch g12 (.nQ(w304), .D(w302), .C(w379), .nC(w1408) );
	vdp_slatch g13 (.Q(w302), .D(DB[7]), .C(w365), .nC(w364) );
	vdp_slatch g14 (.Q(w358), .D(w899), .C(w368), .nC(w367) );
	vdp_sr_bit g15 (.D(w305), .C2(HCLK2), .C1(HCLK1), .Q(FIFOo[7]), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g16 (.A(1'b1), .nZ(DB[7]), .nE(w1407) );
	vdp_notif0 g17 (.A(w304), .nZ(w305), .nE(w1944) );
	vdp_notif0 g18 (.A(w361), .nZ(w355), .nE(w382) );
	vdp_notif0 g19 (.A(w303), .nZ(AD_DATA[7]), .nE(w1553) );
	vdp_notif0 g20 (.A(w363), .nZ(w305), .nE(w1504) );
	vdp_notif0 g21 (.A(w360), .nZ(w355), .nE(w1552) );
	vdp_notif0 g22 (.A(w1480), .nZ(AD_DATA[7]), .nE(w392) );
	vdp_notif0 g23 (.A(w362), .nZ(w305), .nE(w391) );
	vdp_notif0 g24 (.A(w359), .nZ(w355), .nE(w1411) );
	vdp_notif0 g25 (.A(w1479), .nZ(AD_DATA[7]), .nE(w406) );
	vdp_notif0 g26 (.A(w301), .nZ(w305), .nE(w384) );
	vdp_notif0 g27 (.A(w300), .nZ(AD_DATA[7]), .nE(w404) );
	vdp_notif0 g28 (.A(w356), .nZ(DB[7]), .nE(w1550) );
	vdp_notif0 g29 (.nZ(DB[15]), .nE(w385), .A(w6530) );
	vdp_notif0 g30 (.A(w357), .nZ(w355), .nE(w1551) );
	vdp_notif0 g31 (.A(w351), .nZ(DB[15]), .nE(w1549) );
	vdp_notif0 g32 (.A(w420), .nZ(DB[7]), .nE(w386) );
	vdp_aon22 g33 (.Z(w420), .A1(w1474), .A2(w1513), .B1(w390), .B2(w351) );
	vdp_aon22 g34 (.A2(w388), .B1(w389), .B2(AD_DATA[7]), .A1(w355), .Z(w298) );
	vdp_aon22 g35 (.A2(w6436), .B1(w6437), .B2(w355), .A1(AD_DATA[7]), .Z(w299) );
	vdp_aon22 g36 (.Z(w300), .A2(w387), .B1(w1514), .B2(w301), .A1(w357) );
	vdp_aon22 g37 (.Z(w1479), .A2(w411), .B1(w410), .B2(w359), .A1(w362) );
	vdp_aon22 g38 (.Z(w1480), .A2(w418), .B1(w419), .B2(w360), .A1(w363) );
	vdp_aon22 g39 (.Z(w303), .A2(w6432), .B1(w6433), .B2(w304), .A1(w361) );
	vdp_aon22 g40 (.Z(w899), .A1(DB[15]), .A2(w366), .B1(w370), .B2(DB[7]) );
	vdp_slatch g41 (.nQ(w220), .D(VPOS[6]), .C(w1511), .nC(w1512) );
	vdp_slatch g42 (.nQ(w223), .D(HPOS[7]), .C(w372), .nC(w373) );
	vdp_slatch g43 (.nQ(w225), .D(w261), .C(w1413), .nC(w374) );
	vdp_slatch g44 (.nQ(w263), .D(w1379), .C(w1509), .nC(w1510) );
	vdp_slatch g45 (.nQ(w226), .D(w227), .C(w1507), .nC(w1508) );
	vdp_slatch g46 (.nQ(w265), .D(w266), .C(w1505), .nC(w1506) );
	vdp_slatch g47 (.nQ(w228), .D(w227), .C(w375), .nC(w376) );
	vdp_slatch g48 (.nQ(w230), .D(w266), .C(w377), .nC(w378) );
	vdp_slatch g49 (.nQ(w231), .D(w227), .C(w417), .nC(w1410) );
	vdp_slatch g50 (.nQ(w233), .D(w266), .C(w1409), .nC(w383) );
	vdp_slatch g51 (.nQ(w234), .D(w227), .C(w381), .nC(w380) );
	vdp_slatch g52 (.nQ(w268), .D(w266), .C(w379), .nC(w1408) );
	vdp_slatch g53 (.Q(w266), .D(DB[6]), .C(w365), .nC(w364) );
	vdp_slatch g54 (.Q(w227), .D(w269), .C(w368), .nC(w367) );
	vdp_sr_bit g55 (.D(w262), .Q(FIFOo[6]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g56 (.A(1'b1), .nZ(DB[6]), .nE(w1407) );
	vdp_notif0 g57 (.A(w268), .nZ(w262), .nE(w1944) );
	vdp_notif0 g58 (.A(w234), .nZ(RD_DATA[6]), .nE(w382) );
	vdp_notif0 g59 (.A(w267), .nZ(AD_DATA[6]), .nE(w1553) );
	vdp_notif0 g60 (.A(w233), .nZ(w262), .nE(w1504) );
	vdp_notif0 g61 (.A(w231), .nZ(RD_DATA[6]), .nE(w1552) );
	vdp_notif0 g62 (.A(w232), .nZ(AD_DATA[6]), .nE(w392) );
	vdp_notif0 g63 (.A(w230), .nZ(w262), .nE(w391) );
	vdp_notif0 g64 (.A(w228), .nZ(RD_DATA[6]), .nE(w1411) );
	vdp_notif0 g65 (.A(w229), .nZ(AD_DATA[6]), .nE(w406) );
	vdp_notif0 g66 (.A(w265), .nZ(w262), .nE(w384) );
	vdp_notif0 g67 (.A(w264), .nZ(AD_DATA[6]), .nE(w404) );
	vdp_notif0 g68 (.A(w225), .nZ(DB[6]), .nE(w1550) );
	vdp_notif0 g69 (.A(w263), .nZ(DB[14]), .nE(w385) );
	vdp_notif0 g70 (.A(w226), .nZ(RD_DATA[6]), .nE(w1551) );
	vdp_notif0 g71 (.A(w220), .nZ(DB[14]), .nE(w1549) );
	vdp_notif0 g72 (.A(w224), .nZ(DB[6]), .nE(w386) );
	vdp_aon22 g73 (.A2(w1513), .B1(w390), .B2(w220), .A1(w223), .Z(w224) );
	vdp_aon22 g74 (.Z(w261), .A2(w388), .B1(w389), .B2(AD_DATA[6]), .A1(RD_DATA[6]) );
	vdp_aon22 g75 (.Z(w1379), .A2(w6436), .B1(w6437), .B2(RD_DATA[6]), .A1(AD_DATA[6]) );
	vdp_aon22 g76 (.Z(w264), .A2(w387), .B1(w1514), .B2(w265), .A1(w226) );
	vdp_aon22 g77 (.Z(w229), .A2(w411), .B1(w410), .B2(w230), .A1(w228) );
	vdp_aon22 g78 (.Z(w232), .A2(w418), .B1(w419), .B2(w233), .A1(w231) );
	vdp_aon22 g79 (.Z(w267), .A2(w6432), .B1(w6433), .B2(w268), .A1(w234) );
	vdp_aon22 g80 (.Z(w269), .A1(DB[14]), .A2(w366), .B1(w370), .B2(DB[6]) );
	vdp_slatch g81 (.nQ(w335), .D(VPOS[5]), .C(w1511), .nC(w1512) );
	vdp_slatch g82 (.nQ(w1475), .D(HPOS[6]), .C(w372), .nC(w373) );
	vdp_slatch g83 (.nQ(w340), .D(w289), .C(w1413), .nC(w374) );
	vdp_slatch g84 (.D(w290), .C(w1509), .nC(w1510), .nQ(w6531) );
	vdp_slatch g85 (.nQ(w341), .D(w347), .C(w1507), .nC(w1508) );
	vdp_slatch g86 (.nQ(w292), .D(w293), .C(w1505), .nC(w1506) );
	vdp_slatch g87 (.nQ(w343), .D(w347), .C(w375), .nC(w376) );
	vdp_slatch g88 (.nQ(w342), .D(w293), .C(w377), .nC(w378) );
	vdp_slatch g89 (.nQ(w345), .D(w347), .C(w417), .nC(w1410) );
	vdp_slatch g90 (.nQ(w348), .D(w293), .C(w1409), .nC(w383) );
	vdp_slatch g91 (.nQ(w349), .D(w347), .C(w381), .nC(w380) );
	vdp_slatch g92 (.nQ(w295), .D(w293), .C(w379), .nC(w1408) );
	vdp_slatch g93 (.Q(w293), .D(DB[5]), .C(w365), .nC(w364) );
	vdp_slatch g94 (.Q(w347), .D(w296), .C(w368), .nC(w367) );
	vdp_sr_bit g95 (.D(w297), .Q(FIFOo[5]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g96 (.A(1'b1), .nZ(DB[5]), .nE(w1407) );
	vdp_notif0 g97 (.A(w295), .nZ(w297), .nE(w1944) );
	vdp_notif0 g98 (.A(w349), .nZ(RD_DATA[5]), .nE(w382) );
	vdp_notif0 g99 (.A(w294), .nZ(AD_DATA[5]), .nE(w1553) );
	vdp_notif0 g100 (.A(w348), .nZ(w297), .nE(w1504) );
	vdp_notif0 g101 (.A(w345), .nZ(RD_DATA[5]), .nE(w1552) );
	vdp_notif0 g102 (.A(w346), .nZ(AD_DATA[5]), .nE(w392) );
	vdp_notif0 g103 (.A(w342), .nZ(w297), .nE(w391) );
	vdp_notif0 g104 (.A(w343), .nZ(RD_DATA[5]), .nE(w1411) );
	vdp_notif0 g105 (.A(w344), .nZ(AD_DATA[5]), .nE(w406) );
	vdp_notif0 g106 (.A(w292), .nZ(w297), .nE(w384) );
	vdp_notif0 g107 (.A(w291), .nZ(AD_DATA[5]), .nE(w404) );
	vdp_notif0 g108 (.A(w340), .nZ(DB[5]), .nE(w1550) );
	vdp_notif0 g109 (.nZ(DB[13]), .nE(w385), .A(w6531) );
	vdp_notif0 g110 (.A(w341), .nZ(RD_DATA[5]), .nE(w1551) );
	vdp_notif0 g111 (.A(w335), .nZ(DB[13]), .nE(w1549) );
	vdp_notif0 g112 (.A(w339), .nZ(DB[5]), .nE(w386) );
	vdp_aon22 g113 (.Z(w339), .A1(w1475), .A2(w1513), .B1(w390), .B2(w335) );
	vdp_aon22 g114 (.A2(w388), .B1(w389), .B2(AD_DATA[5]), .A1(RD_DATA[5]), .Z(w289) );
	vdp_aon22 g115 (.A2(w6436), .B1(w6437), .B2(RD_DATA[5]), .A1(AD_DATA[5]), .Z(w290) );
	vdp_aon22 g116 (.Z(w291), .A2(w387), .B1(w1514), .B2(w292), .A1(w341) );
	vdp_aon22 g117 (.Z(w344), .A2(w411), .B1(w410), .B2(w343), .A1(w342) );
	vdp_aon22 g118 (.Z(w346), .A2(w418), .B1(w419), .B2(w345), .A1(w348) );
	vdp_aon22 g119 (.Z(w294), .A2(w6432), .B1(w6433), .B2(w295), .A1(w349) );
	vdp_aon22 g120 (.Z(w296), .A1(DB[13]), .A2(w366), .B1(w370), .B2(DB[5]) );
	vdp_slatch g121 (.nQ(w205), .D(VPOS[4]), .C(w1511), .nC(w1512) );
	vdp_slatch g122 (.nQ(w208), .D(HPOS[5]), .C(w372), .nC(w373) );
	vdp_slatch g123 (.nQ(w1515), .D(w253), .C(w1413), .nC(w374) );
	vdp_slatch g124 (.D(w1478), .C(w1509), .nC(w1510), .nQ(w6532) );
	vdp_slatch g125 (.nQ(w210), .D(w211), .C(w1507), .nC(w1508) );
	vdp_slatch g126 (.nQ(w256), .D(w257), .C(w1505), .nC(w1506) );
	vdp_slatch g127 (.nQ(w212), .D(w211), .C(w375), .nC(w376) );
	vdp_slatch g128 (.nQ(w214), .D(w257), .C(w377), .nC(w378) );
	vdp_slatch g129 (.nQ(w215), .D(w211), .C(w417), .nC(w1410) );
	vdp_slatch g130 (.nQ(w217), .D(w257), .C(w1409), .nC(w383) );
	vdp_slatch g131 (.nQ(w218), .D(w211), .C(w381), .nC(w380) );
	vdp_slatch g132 (.nQ(w259), .D(w257), .C(w379), .nC(w1408) );
	vdp_slatch g133 (.Q(w257), .D(DB[4]), .C(w365), .nC(w364) );
	vdp_slatch g134 (.Q(w211), .D(w260), .C(w368), .nC(w367) );
	vdp_sr_bit g135 (.D(w254), .Q(FIFOo[4]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g136 (.A(1'b1), .nZ(DB[4]), .nE(w1407) );
	vdp_notif0 g137 (.A(w259), .nZ(w254), .nE(w1944) );
	vdp_notif0 g138 (.A(w218), .nZ(RD_DATA[4]), .nE(w382) );
	vdp_notif0 g139 (.A(w258), .nZ(AD_DATA[4]), .nE(w1553) );
	vdp_notif0 g140 (.A(w217), .nZ(w254), .nE(w1504) );
	vdp_notif0 g141 (.A(w215), .nZ(RD_DATA[4]), .nE(w1552) );
	vdp_notif0 g142 (.A(w216), .nZ(AD_DATA[4]), .nE(w392) );
	vdp_notif0 g143 (.A(w214), .nZ(w254), .nE(w391) );
	vdp_notif0 g144 (.A(w212), .nZ(RD_DATA[4]), .nE(w1411) );
	vdp_notif0 g145 (.A(w213), .nZ(AD_DATA[4]), .nE(w406) );
	vdp_notif0 g146 (.A(w256), .nZ(w254), .nE(w384) );
	vdp_notif0 g147 (.A(w255), .nZ(AD_DATA[4]), .nE(w404) );
	vdp_notif0 g148 (.A(w1515), .nZ(DB[4]), .nE(w1550) );
	vdp_notif0 g149 (.nZ(DB[12]), .nE(w385), .A(w6532) );
	vdp_notif0 g150 (.A(w210), .nZ(RD_DATA[4]), .nE(w1551) );
	vdp_notif0 g151 (.A(w205), .nZ(DB[12]), .nE(w1549) );
	vdp_notif0 g152 (.A(w209), .nZ(DB[4]), .nE(w386) );
	vdp_aon22 g153 (.A2(w1513), .B1(w390), .B2(w205), .A1(w208), .Z(w209) );
	vdp_aon22 g154 (.Z(w253), .A2(w388), .B1(w389), .B2(AD_DATA[4]), .A1(RD_DATA[4]) );
	vdp_aon22 g155 (.Z(w1478), .A2(w6436), .B1(w6437), .B2(RD_DATA[4]), .A1(AD_DATA[4]) );
	vdp_aon22 g156 (.Z(w255), .A2(w387), .B1(w1514), .B2(w256), .A1(w210) );
	vdp_aon22 g157 (.Z(w213), .A2(w411), .B1(w410), .B2(w214), .A1(w212) );
	vdp_aon22 g158 (.Z(w216), .A2(w418), .B1(w419), .B2(w217), .A1(w215) );
	vdp_aon22 g159 (.Z(w258), .A2(w6432), .B1(w6433), .B2(w259), .A1(w218) );
	vdp_aon22 g160 (.Z(w260), .A1(DB[12]), .A2(w366), .B1(w370), .B2(DB[4]) );
	vdp_slatch g161 (.nQ(w319), .D(VPOS[3]), .C(w1511), .nC(w1512) );
	vdp_slatch g162 (.nQ(w1476), .D(HPOS[4]), .C(w372), .nC(w373) );
	vdp_slatch g163 (.nQ(w324), .D(w280), .C(w1413), .nC(w374) );
	vdp_slatch g164 (.D(w281), .C(w1509), .nC(w1510), .nQ(w6533) );
	vdp_slatch g165 (.nQ(w325), .D(w328), .C(w1507), .nC(w1508) );
	vdp_slatch g166 (.nQ(w283), .D(w284), .C(w1505), .nC(w1506) );
	vdp_slatch g167 (.nQ(w326), .D(w328), .C(w375), .nC(w376) );
	vdp_slatch g168 (.nQ(w327), .D(w284), .C(w377), .nC(w378) );
	vdp_slatch g169 (.nQ(w330), .D(w328), .C(w417), .nC(w1410) );
	vdp_slatch g170 (.nQ(w332), .D(w284), .C(w1409), .nC(w383) );
	vdp_slatch g171 (.nQ(w333), .D(w328), .C(w381), .nC(w380) );
	vdp_slatch g172 (.nQ(w286), .D(w284), .C(w379), .nC(w1408) );
	vdp_slatch g173 (.Q(w284), .D(DB[3]), .C(w365), .nC(w364) );
	vdp_slatch g174 (.Q(w328), .D(w287), .C(w368), .nC(w367) );
	vdp_sr_bit g175 (.D(w288), .Q(FIFOo[3]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g176 (.A(1'b1), .nZ(DB[3]), .nE(w1407) );
	vdp_notif0 g177 (.A(w286), .nZ(w288), .nE(w1944) );
	vdp_notif0 g178 (.A(w333), .nZ(w321), .nE(w382) );
	vdp_notif0 g179 (.A(w285), .nZ(AD_DATA[3]), .nE(w1553) );
	vdp_notif0 g180 (.A(w332), .nZ(w288), .nE(w1504) );
	vdp_notif0 g181 (.A(w330), .nZ(w321), .nE(w1552) );
	vdp_notif0 g182 (.A(w331), .nZ(AD_DATA[3]), .nE(w392) );
	vdp_notif0 g183 (.A(w327), .nZ(w288), .nE(w391) );
	vdp_notif0 g184 (.A(w326), .nZ(w321), .nE(w1411) );
	vdp_notif0 g185 (.A(w329), .nZ(AD_DATA[3]), .nE(w406) );
	vdp_notif0 g186 (.A(w283), .nZ(w288), .nE(w384) );
	vdp_notif0 g187 (.A(w282), .nZ(AD_DATA[3]), .nE(w404) );
	vdp_notif0 g188 (.A(w324), .nZ(DB[3]), .nE(w1550) );
	vdp_notif0 g189 (.nZ(DB[11]), .nE(w385), .A(w6533) );
	vdp_notif0 g190 (.A(w325), .nZ(w321), .nE(w1551) );
	vdp_notif0 g191 (.A(w319), .nZ(DB[11]), .nE(w1549) );
	vdp_notif0 g192 (.A(w323), .nZ(DB[3]), .nE(w386) );
	vdp_aon22 g193 (.Z(w323), .A1(w1476), .A2(w1513), .B1(w390), .B2(w319) );
	vdp_aon22 g194 (.A2(w388), .B1(w389), .B2(AD_DATA[3]), .A1(w321), .Z(w280) );
	vdp_aon22 g195 (.A2(w6436), .B1(w6437), .B2(w321), .A1(AD_DATA[3]), .Z(w281) );
	vdp_aon22 g196 (.Z(w282), .A2(w387), .B1(w1514), .B2(w283), .A1(w325) );
	vdp_aon22 g197 (.Z(w329), .A2(w411), .B1(w410), .B2(w326), .A1(w327) );
	vdp_aon22 g198 (.Z(w331), .A2(w418), .B1(w419), .B2(w330), .A1(w332) );
	vdp_aon22 g199 (.Z(w285), .A2(w6432), .B1(w6433), .B2(w286), .A1(w333) );
	vdp_aon22 g200 (.Z(w287), .A1(DB[11]), .A2(w366), .B1(w370), .B2(DB[3]) );
	vdp_slatch g201 (.nQ(w191), .D(VPOS[2]), .C(w1511), .nC(w1512) );
	vdp_slatch g202 (.nQ(w1516), .D(HPOS[3]), .C(w372), .nC(w373) );
	vdp_slatch g203 (.nQ(w193), .D(w244), .C(w1413), .nC(w374) );
	vdp_slatch g204 (.D(w1414), .C(w1509), .nC(w1510), .nQ(w6534) );
	vdp_slatch g205 (.nQ(w194), .D(w197), .C(w1507), .nC(w1508) );
	vdp_slatch g206 (.nQ(w247), .D(w248), .C(w1505), .nC(w1506) );
	vdp_slatch g207 (.nQ(w195), .D(w197), .C(w375), .nC(w376) );
	vdp_slatch g208 (.nQ(w198), .D(w248), .C(w377), .nC(w378) );
	vdp_slatch g209 (.nQ(w199), .D(w197), .C(w417), .nC(w1410) );
	vdp_slatch g210 (.nQ(w201), .D(w248), .C(w1409), .nC(w383) );
	vdp_slatch g211 (.nQ(w202), .D(w197), .C(w381), .nC(w380) );
	vdp_slatch g212 (.nQ(w250), .D(w248), .C(w379), .nC(w1408) );
	vdp_slatch g213 (.Q(w248), .D(DB[2]), .C(w365), .nC(w364) );
	vdp_slatch g214 (.Q(w197), .D(w251), .C(w368), .nC(w367) );
	vdp_sr_bit g215 (.D(w245), .Q(FIFOo[2]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g216 (.A(w203), .nZ(DB[2]), .nE(w1407) );
	vdp_notif0 g217 (.A(w250), .nZ(w245), .nE(w1944) );
	vdp_notif0 g218 (.A(w202), .nZ(RD_DATA[2]), .nE(w382) );
	vdp_notif0 g219 (.A(w249), .nZ(AD_DATA[2]), .nE(w1553) );
	vdp_notif0 g220 (.A(w201), .nZ(w245), .nE(w1504) );
	vdp_notif0 g221 (.A(w199), .nZ(RD_DATA[2]), .nE(w1552) );
	vdp_notif0 g222 (.A(w200), .nZ(AD_DATA[2]), .nE(w392) );
	vdp_notif0 g223 (.A(w198), .nZ(w245), .nE(w391) );
	vdp_notif0 g224 (.A(w195), .nZ(RD_DATA[2]), .nE(w1411) );
	vdp_notif0 g225 (.A(w196), .nZ(AD_DATA[2]), .nE(w406) );
	vdp_notif0 g226 (.A(w247), .nZ(w245), .nE(w384) );
	vdp_notif0 g227 (.A(w246), .nZ(AD_DATA[2]), .nE(w404) );
	vdp_notif0 g228 (.A(w193), .nZ(DB[2]), .nE(w1550) );
	vdp_notif0 g229 (.nZ(DB[10]), .nE(w385), .A(w6534) );
	vdp_notif0 g230 (.A(w194), .nZ(RD_DATA[2]), .nE(w1551) );
	vdp_notif0 g231 (.A(w191), .nZ(DB[10]), .nE(w1549) );
	vdp_notif0 g232 (.A(w192), .nZ(DB[2]), .nE(w386) );
	vdp_aon22 g233 (.A2(w1513), .B1(w390), .B2(w191), .A1(w1516), .Z(w192) );
	vdp_aon22 g234 (.Z(w244), .A2(w388), .B1(w389), .B2(AD_DATA[2]), .A1(RD_DATA[2]) );
	vdp_aon22 g235 (.Z(w1414), .A2(w6436), .B1(w6437), .B2(RD_DATA[2]), .A1(AD_DATA[2]) );
	vdp_aon22 g236 (.Z(w246), .A2(w387), .B1(w1514), .B2(w247), .A1(w194) );
	vdp_aon22 g237 (.Z(w196), .A2(w411), .B1(w410), .B2(w198), .A1(w195) );
	vdp_aon22 g238 (.Z(w200), .A2(w418), .B1(w419), .B2(w201), .A1(w199) );
	vdp_aon22 g239 (.Z(w249), .A2(w6432), .B1(w6433), .B2(w250), .A1(w202) );
	vdp_aon22 g240 (.Z(w251), .A1(DB[10]), .A2(w366), .B1(w370), .B2(DB[2]) );
	vdp_slatch g241 (.nQ(w306), .D(VPOS[1]), .C(w1511), .nC(w1512) );
	vdp_slatch g242 (.nQ(w1477), .D(HPOS[2]), .C(w372), .nC(w373) );
	vdp_slatch g243 (.nQ(w309), .D(w270), .C(w1413), .nC(w374) );
	vdp_slatch g244 (.D(w271), .C(w1509), .nC(w1510), .nQ(w6535) );
	vdp_slatch g245 (.nQ(w310), .D(w313), .C(w1507), .nC(w1508) );
	vdp_slatch g246 (.nQ(w273), .D(w274), .C(w1505), .nC(w1506) );
	vdp_slatch g247 (.nQ(w312), .D(w313), .C(w375), .nC(w376) );
	vdp_slatch g248 (.nQ(w311), .D(w274), .C(w377), .nC(w378) );
	vdp_slatch g249 (.nQ(w315), .D(w313), .C(w417), .nC(w1410) );
	vdp_slatch g250 (.nQ(w317), .D(w274), .C(w1409), .nC(w383) );
	vdp_slatch g251 (.nQ(w318), .D(w313), .C(w381), .nC(w380) );
	vdp_slatch g252 (.nQ(w276), .D(w274), .C(w379), .nC(w1408) );
	vdp_slatch g253 (.Q(w274), .D(DB[1]), .C(w365), .nC(w364) );
	vdp_slatch g254 (.Q(w313), .D(w278), .C(w368), .nC(w367) );
	vdp_sr_bit g255 (.D(w279), .Q(FIFOo[1]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g256 (.A(w1554), .nZ(DB[1]), .nE(w1407) );
	vdp_notif0 g257 (.A(w276), .nZ(w279), .nE(w1944) );
	vdp_notif0 g258 (.A(w318), .nZ(RD_DATA[1]), .nE(w382) );
	vdp_notif0 g259 (.A(w275), .nZ(AD_DATA[1]), .nE(w1553) );
	vdp_notif0 g260 (.A(w317), .nZ(w279), .nE(w1504) );
	vdp_notif0 g261 (.A(w315), .nZ(RD_DATA[1]), .nE(w1552) );
	vdp_notif0 g262 (.A(w316), .nZ(AD_DATA[1]), .nE(w392) );
	vdp_notif0 g263 (.A(w311), .nZ(w279), .nE(w391) );
	vdp_notif0 g264 (.A(w312), .nZ(RD_DATA[1]), .nE(w1411) );
	vdp_notif0 g265 (.A(w314), .nZ(AD_DATA[1]), .nE(w406) );
	vdp_notif0 g266 (.A(w273), .nZ(w279), .nE(w384) );
	vdp_notif0 g267 (.A(w272), .nZ(AD_DATA[1]), .nE(w404) );
	vdp_notif0 g268 (.A(w309), .nZ(DB[1]), .nE(w1550) );
	vdp_notif0 g269 (.nZ(DB[9]), .nE(w385), .A(w6535) );
	vdp_notif0 g270 (.A(w310), .nZ(RD_DATA[1]), .nE(w1551) );
	vdp_notif0 g271 (.A(w306), .nZ(DB[9]), .nE(w1549) );
	vdp_notif0 g272 (.A(w1412), .nZ(DB[1]), .nE(w386) );
	vdp_aon22 g273 (.Z(w1412), .A1(w1477), .A2(w1513), .B1(w390), .B2(w306) );
	vdp_aon22 g274 (.A2(w388), .B1(w389), .B2(AD_DATA[1]), .A1(RD_DATA[1]), .Z(w270) );
	vdp_aon22 g275 (.A2(w6436), .B1(w6437), .B2(RD_DATA[1]), .A1(AD_DATA[1]), .Z(w271) );
	vdp_aon22 g276 (.Z(w272), .A2(w387), .B1(w1514), .B2(w273), .A1(w310) );
	vdp_aon22 g277 (.Z(w314), .A2(w411), .B1(w410), .B2(w312), .A1(w311) );
	vdp_aon22 g278 (.Z(w316), .A2(w418), .B1(w419), .B2(w315), .A1(w317) );
	vdp_aon22 g279 (.Z(w275), .A2(w6432), .B1(w6433), .B2(w276), .A1(w318) );
	vdp_aon22 g280 (.Z(w278), .A1(DB[9]), .A2(w366), .B1(w370), .B2(DB[1]) );
	vdp_slatch g281 (.nQ(w176), .D(VPOS_80), .C(w1511), .nC(w1512) );
	vdp_slatch g282 (.D(HPOS[1]), .nQ(w1406), .C(w372), .nC(w373) );
	vdp_slatch g283 (.nQ(w178), .D(w236), .C(w1413), .nC(w374) );
	vdp_slatch g284 (.D(w1381), .C(w1509), .nC(w1510), .nQ(w6536) );
	vdp_slatch g285 (.nQ(w179), .D(w183), .C(w1507), .nC(w1508) );
	vdp_slatch g286 (.nQ(w239), .D(w240), .C(w1505), .nC(w1506) );
	vdp_slatch g287 (.nQ(w180), .D(w183), .C(w375), .nC(w376) );
	vdp_slatch g288 (.nQ(w182), .D(w240), .C(w377), .nC(w378) );
	vdp_slatch g289 (.nQ(w184), .D(w183), .C(w417), .nC(w1410) );
	vdp_slatch g290 (.nQ(w186), .D(w240), .C(w1409), .nC(w383) );
	vdp_slatch g291 (.nQ(w187), .D(w183), .C(w381), .nC(w380) );
	vdp_slatch g292 (.nQ(w242), .D(w240), .C(w379), .nC(w1408) );
	vdp_slatch g293 (.Q(w240), .D(DB[0]), .C(w365), .nC(w364) );
	vdp_slatch g294 (.D(w243), .Q(w183), .C(w368), .nC(w367) );
	vdp_sr_bit g295 (.D(w237), .C2(HCLK2), .C1(HCLK1), .Q(FIFOo[0]), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g296 (.A(1'b1), .nZ(DB[0]), .nE(w1407) );
	vdp_notif0 g297 (.A(w242), .nZ(w237), .nE(w1944) );
	vdp_notif0 g298 (.A(w187), .nZ(RD_DATA[0]), .nE(w382) );
	vdp_notif0 g299 (.A(w241), .nZ(AD_DATA[0]), .nE(w1553) );
	vdp_notif0 g300 (.A(w186), .nZ(w237), .nE(w1504) );
	vdp_notif0 g301 (.A(w184), .nZ(RD_DATA[0]), .nE(w1552) );
	vdp_notif0 g302 (.A(w185), .nZ(AD_DATA[0]), .nE(w392) );
	vdp_notif0 g303 (.A(w182), .nZ(w237), .nE(w391) );
	vdp_notif0 g304 (.A(w180), .nZ(RD_DATA[0]), .nE(w1411) );
	vdp_notif0 g305 (.A(w181), .nZ(AD_DATA[0]), .nE(w406) );
	vdp_notif0 g306 (.A(w239), .nZ(w237), .nE(w384) );
	vdp_notif0 g307 (.A(w238), .nZ(AD_DATA[0]), .nE(w404) );
	vdp_notif0 g308 (.A(w178), .nZ(DB[0]), .nE(w1550) );
	vdp_notif0 g309 (.nZ(DB[8]), .nE(w385), .A(w6536) );
	vdp_notif0 g310 (.A(w179), .nZ(RD_DATA[0]), .nE(w1551) );
	vdp_notif0 g311 (.A(w176), .nZ(DB[8]), .nE(w1549) );
	vdp_notif0 g312 (.A(w177), .nZ(DB[0]), .nE(w386) );
	vdp_aon22 g313 (.A2(w1513), .B1(w390), .B2(w176), .A1(w1406), .Z(w177) );
	vdp_aon22 g314 (.Z(w236), .A2(w388), .B1(w389), .B2(AD_DATA[0]), .A1(RD_DATA[0]) );
	vdp_aon22 g315 (.Z(w1381), .A2(w6436), .B1(w6437), .B2(RD_DATA[0]), .A1(AD_DATA[0]) );
	vdp_aon22 g316 (.Z(w238), .A2(w387), .B1(w1514), .B2(w239), .A1(w179) );
	vdp_aon22 g317 (.Z(w181), .A2(w411), .B1(w410), .B2(w182), .A1(w180) );
	vdp_aon22 g318 (.Z(w185), .A2(w418), .B1(w419), .B2(w186), .A1(w184) );
	vdp_aon22 g319 (.Z(w241), .A2(w6432), .B1(w6433), .B2(w242), .A1(w187) );
	vdp_aon22 g320 (.Z(w243), .A1(DB[8]), .A2(w366), .B1(w370), .B2(DB[0]) );
	vdp_not g321 (.A(w277), .nZ(w1554) );
	vdp_not g322 (.A(w252), .nZ(w203) );
	vdp_not g323 (.A(w394), .nZ(w1549) );
	vdp_not g324 (.A(w398), .nZ(w386) );
	vdp_not g325 (.A(w403), .nZ(w1550) );
	vdp_not g326 (.A(w403), .nZ(w385) );
	vdp_sr_bit g327 (.D(w402), .C2(HCLK2), .C1(HCLK1), .Q(w914), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g328 (.D(w447), .Q(w416), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g329 (.D(w416), .Q(w414), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g330 (.D(w414), .Q(w408), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g331 (.D(w412), .Q(w453), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g332 (.D(w453), .Q(w409), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g333 (.D(w454), .Q(w402), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g334 (.D(w405), .Q(w399), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g335 (.A(w436), .nZ(w1551) );
	vdp_not g336 (.A(w436), .nZ(w404) );
	vdp_not g337 (.A(w436), .nZ(w384) );
	vdp_not g338 (.A(w438), .nZ(w1411) );
	vdp_not g339 (.A(w438), .nZ(w406) );
	vdp_not g340 (.A(w438), .nZ(w391) );
	vdp_not g341 (.A(w450), .nZ(w1552) );
	vdp_not g342 (.A(w450), .nZ(w392) );
	vdp_not g343 (.A(w450), .nZ(w1504) );
	vdp_not g344 (.A(w439), .nZ(w382) );
	vdp_not g345 (.A(w439), .nZ(w1553) );
	vdp_not g346 (.A(w439), .nZ(w1944) );
	vdp_not g347 (.A(w987), .nZ(w1407) );
	vdp_not g348 (.A(w414), .nZ(w393) );
	vdp_not g349 (.A(SEL0_M3), .nZ(w396) );
	vdp_comp_str g350 (.A(w429), .Z(w1511), .nZ(w1512) );
	vdp_comp_str g351 (.A(w430), .Z(w372), .nZ(w373) );
	vdp_comp_str g352 (.A(w400), .Z(w1413), .nZ(w374) );
	vdp_comp_str g353 (.A(w401), .Z(w1509), .nZ(w1510) );
	vdp_comp_str g354 (.A(w455), .Z(w1507), .nZ(w1508) );
	vdp_comp_str g355 (.A(w455), .Z(w1505), .nZ(w1506) );
	vdp_comp_str g356 (.A(w452), .Z(w375), .nZ(w376) );
	vdp_comp_str g357 (.A(w452), .Z(w377), .nZ(w378) );
	vdp_comp_str g358 (.A(w495), .Z(w417), .nZ(w1410) );
	vdp_comp_str g359 (.A(w495), .Z(w1409), .nZ(w383) );
	vdp_comp_str g360 (.A(w446), .Z(w381), .nZ(w380) );
	vdp_comp_str g361 (.A(w446), .Z(w379), .nZ(w1408) );
	vdp_comp_str g362 (.A(w456), .Z(w365), .nZ(w364) );
	vdp_comp_str g363 (.A(w456), .Z(w368), .nZ(w367) );
	vdp_comp_we g364 (.A(SEL0_M3), .Z(w366), .nZ(w370) );
	vdp_comp_we g365 (.A(w435), .Z(w6432), .nZ(w6433) );
	vdp_comp_we g366 (.A(w435), .Z(w418), .nZ(w419) );
	vdp_comp_we g367 (.A(w435), .Z(w411), .nZ(w410) );
	vdp_comp_we g368 (.A(w435), .Z(w387), .nZ(w1514) );
	vdp_comp_we g369 (.A(w440), .Z(w6436), .nZ(w6437) );
	vdp_comp_we g370 (.A(w397), .Z(w388), .nZ(w389) );
	vdp_comp_we g371 (.A(w433), .Z(w1513), .nZ(w390) );
	vdp_and g372 (.Z(w400), .B(HCLK1), .A(w399) );
	vdp_and g373 (.Z(w401), .B(HCLK1), .A(w402) );
	vdp_and g374 (.Z(w405), .B(w409), .A(w407) );
	vdp_and g375 (.Z(w454), .B(w409), .A(w413) );
	vdp_nand g376 (.Z(w413), .B(w440), .A(w393) );
	vdp_nand g377 (.Z(w407), .B(w440), .A(w414) );
	vdp_and3 g378 (.Z(w440), .B(w426), .A(SEL0_M3), .C(w427) );
	vdp_and3 g379 (.Z(w397), .B(w396), .A(w408), .C(VRAM128k) );
	vdp_not g380 (.A(VRAM128k), .nZ(w427) );
	vdp_sr_bit g381 (.D(w424), .C2(HCLK2), .C1(HCLK1), .Q(w423), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g382 (.D(w1390), .Q(w460), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g383 (.D(w1469), .C2(HCLK2), .C1(HCLK1), .Q(w486), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g384 (.A(w487), .nZ(w415) );
	vdp_fa g385 (.SUM(w448), .A(w486), .B(1'b0), .CI(w488) );
	vdp_not g386 (.A(w424), .nZ(w422) );
	vdp_not g387 (.A(M5), .nZ(w459) );
	vdp_not g388 (.A(w432), .nZ(w430) );
	vdp_not g389 (.A(w442), .nZ(w443) );
	vdp_not g390 (.A(w493), .nZ(w445) );
	vdp_not g391 (.A(w486), .nZ(w444) );
	vdp_slatch g392 (.Q(w480), .D(w484), .C(w466), .nC(w421) );
	vdp_slatch g393 (.Q(w1457), .D(w484), .C(w478), .nC(w451) );
	vdp_slatch g394 (.Q(w481), .D(w484), .C(w464), .nC(w437) );
	vdp_slatch g395 (.Q(w482), .D(w484), .C(w462), .nC(w434) );
	vdp_slatch g396 (.Q(w483), .D(w457), .C(w466), .nC(w421) );
	vdp_slatch g397 (.Q(w485), .D(w457), .C(w478), .nC(w451) );
	vdp_slatch g398 (.Q(w1456), .D(w457), .E(w464), .nE(w437) );
	vdp_slatch g399 (.Q(w479), .D(w457), .C(w462), .nC(w434) );
	vdp_slatch g400 (.Q(w471), .D(w458), .C(w466), .nC(w421) );
	vdp_slatch g401 (.Q(w465), .D(w458), .C(w478), .nC(w451) );
	vdp_slatch g402 (.Q(w469), .D(w458), .C(w464), .nC(w437) );
	vdp_slatch g403 (.Q(w472), .D(w458), .C(w462), .nC(w434) );
	vdp_comp_dff g404 (.D(w428), .C2(HCLK2), .C1(HCLK1), .Q(w424), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and g405 (.Z(w1390), .B(w422), .A(w423) );
	vdp_or g406 (.Z(w429), .B(w459), .A(w430) );
	vdp_or g407 (.Z(w433), .B(CA[0]), .A(SEL0_M3) );
	vdp_and3 g408 (.Z(w436), .B(w487), .A(w444), .C(w493) );
	vdp_and3 g409 (.Z(w438), .B(w487), .A(w445), .C(w486) );
	vdp_and3 g410 (.Z(w439), .B(w444), .A(w445), .C(w487) );
	vdp_xor g411 (.Z(w441), .B(w491), .A(w490) );
	vdp_aon22 g412 (.Z(w435), .A1(w443), .A2(w491), .B1(w508), .B2(w442) );
	vdp_and3 g413 (.Z(w450), .B(w486), .A(w493), .C(w487) );
	vdp_comp_str g414 (.A(w495), .Z(w466), .nZ(w421) );
	vdp_comp_str g415 (.A(w446), .Z(w462), .nZ(w434) );
	vdp_comp_str g416 (.A(w455), .Z(w464), .nZ(w437) );
	vdp_comp_str g417 (.A(w452), .Z(w478), .nZ(w451) );
	vdp_nand g418 (.Z(w442), .B(w492), .A(w441) );
	vdp_and g419 (.Z(w1469), .B(w489), .A(w448) );
	vdp_aoi21 g420 (.Z(w432), .B(w431), .A1(HCLK1), .A2(w460) );
	vdp_nor g421 (.Z(w431), .B(M3), .A(w459) );
	vdp_nor g422 (.Z(w426), .B(w457), .A(w458) );
	vdp_not g423 (.A(w474), .nZ(w534) );
	vdp_not g424 (.A(w473), .nZ(w538) );
	vdp_nor g425 (.Z(w596), .A(w519), .B(w474) );
	vdp_or g426 (.A(w1389), .Z(w475), .B(w476) );
	vdp_comp_we g427 (.A(w571), .nZ(w467), .Z(w513) );
	vdp_aon22 g428 (.Z(w473), .A1(w513), .A2(w458), .B1(w467), .B2(w477) );
	vdp_aon22 g429 (.Z(w537), .A1(w513), .A2(w498), .B1(w467), .B2(w475) );
	vdp_aon22 g430 (.Z(w528), .A1(w513), .A2(w524), .B1(w467), .B2(w490) );
	vdp_aon22 g431 (.Z(w474), .A1(w513), .A2(w457), .B1(w467), .B2(w520) );
	vdp_aon22 g432 (.Z(w533), .A1(w513), .A2(w518), .B1(w467), .B2(w491) );
	vdp_aon22 g433 (.Z(w519), .A1(w513), .A2(w484), .B1(w467), .B2(w512) );
	vdp_and g434 (.Z(w532), .A(w511), .B(w510) );
	vdp_and g435 (.Z(w470), .A(w511), .B(w493) );
	vdp_and g436 (.Z(w1458), .A(w486), .B(w510) );
	vdp_and g437 (.Z(w468), .A(w486), .B(w493) );
	vdp_and g438 (.Z(w1391), .A(w489), .B(w506) );
	vdp_fa g439 (.SUM(w506), .A(w493), .B(w494), .CO(w488), .CI(w507) );
	vdp_sr_bit g440 (.D(w1391), .C2(HCLK2), .C1(HCLK1), .Q(w493), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g441 (.A(w509), .nZ(w1393) );
	vdp_not g442 (.A(w499), .nZ(w502) );
	vdp_and g443 (.Z(w494), .A(w567), .B(w1393) );
	vdp_and3 g444 (.Z(w452), .B(w500), .A(w499), .C(w503) );
	vdp_and3 g445 (.Z(w495), .B(w500), .A(w499), .C(w501) );
	vdp_xor g446 (.Z(w505), .A(w486), .B(w499) );
	vdp_not g447 (.A(w493), .nZ(w510) );
	vdp_not g448 (.A(w486), .nZ(w511) );
	vdp_not g449 (.A(w492), .nZ(w1392) );
	vdp_and5 g450 (.Z(w36), .A(w535), .B(w528), .C(w539), .D(w538), .E(w474) );
	vdp_and5 g451 (.Z(w35), .A(w535), .B(w533), .C(w539), .D(w538), .E(w474) );
	vdp_aon2222 g452 (.C2(w529), .B2(w527), .A2(w526), .C1(w1458), .B1(w470), .A1(w532), .Z(w476), .D2(w530), .D1(w468) );
	vdp_aon2222 g453 (.C2(w465), .B2(w469), .A2(w472), .C1(w1458), .B1(w470), .A1(w532), .Z(w477), .D2(w471), .D1(w468) );
	vdp_aon2222 g454 (.C2(w1404), .B2(w523), .A2(w1405), .C1(w1458), .B1(w470), .A1(w532), .Z(w490), .D2(w521), .D1(w468) );
	vdp_aon2222 g455 (.C2(w485), .B2(w1456), .A2(w479), .C1(w1458), .B1(w470), .A1(w532), .Z(w520), .D2(w483), .D1(w468) );
	vdp_aon2222 g456 (.C2(w1459), .B2(w517), .A2(w514), .C1(w1458), .B1(w470), .A1(w532), .Z(w491), .D2(w531), .D1(w468) );
	vdp_aon2222 g457 (.C2(w1457), .B2(w481), .A2(w482), .C1(w1458), .B1(w470), .A1(w532), .Z(w512), .D2(w480), .D1(w468) );
	vdp_nor g458 (.Z(w509), .A(w1392), .B(w441) );
	vdp_or g459 (.Z(w456), .B(w496), .A(w941) );
	vdp_cnt_bit g460 (.R(SYSRES), .Q(w499), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2), .CI(w497) );
	vdp_cnt_bit g461 (.R(SYSRES), .Q(w501), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2), .CI(w560), .CO(w497) );
	vdp_not g462 (.A(w501), .nZ(w503) );
	vdp_not g463 (.A(w1394), .nZ(w500) );
	vdp_and3 g464 (.Z(w446), .B(w500), .A(w502), .C(w503) );
	vdp_and3 g465 (.Z(w455), .B(w500), .A(w502), .C(w501) );
	vdp_xor g466 (.Z(w504), .A(w493), .B(w501) );
	vdp_fa g467 (.SUM(w1518), .A(w568), .B(w508), .CO(w507), .CI(1'b0) );
	vdp_and g468 (.Z(w568), .A(w509), .B(w567) );
	vdp_and g469 (.Z(w1403), .A(w489), .B(w1518) );
	vdp_sr_bit g470 (.D(w1403), .C2(HCLK2), .C1(HCLK1), .Q(w508), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g471 (.A(w1401), .nZ(w553) );
	vdp_comp_str g472 (.A(w446), .Z(w547), .nZ(w525) );
	vdp_comp_str g473 (.A(w455), .Z(w555), .nZ(w515) );
	vdp_comp_str g474 (.A(w452), .Z(w554), .nZ(w522) );
	vdp_comp_str g475 (.A(w495), .Z(w556), .nZ(w516) );
	vdp_slatch g476 (.Q(w531), .D(w518), .C(w556), .nC(w516) );
	vdp_slatch g477 (.Q(w1459), .D(w518), .C(w554), .nC(w522) );
	vdp_slatch g478 (.Q(w517), .D(w518), .C(w555), .nC(w515) );
	vdp_slatch g479 (.Q(w514), .D(w518), .C(w547), .nC(w525) );
	vdp_slatch g480 (.Q(w521), .D(w524), .C(w556), .nC(w516) );
	vdp_slatch g481 (.Q(w1404), .D(w524), .C(w554), .nC(w522) );
	vdp_slatch g482 (.Q(w523), .D(w524), .C(w555), .nC(w515) );
	vdp_slatch g483 (.Q(w1405), .D(w524), .C(w547), .nC(w525) );
	vdp_slatch g484 (.Q(w530), .D(w498), .C(w556), .nC(w516) );
	vdp_slatch g485 (.Q(w529), .D(w498), .C(w554), .nC(w522) );
	vdp_slatch g486 (.Q(w527), .D(w498), .C(w555), .nC(w515) );
	vdp_slatch g487 (.Q(w526), .D(w498), .C(w547), .nC(w525) );
	vdp_and5 g488 (.Z(w173), .A(w535), .B(w528), .C(w538), .D(w519), .E(w534) );
	vdp_and5 g489 (.Z(w172), .A(w535), .B(w533), .C(w538), .D(w519), .E(w534) );
	vdp_not g490 (.A(M5), .nZ(w1389) );
	vdp_not g491 (.A(w519), .nZ(w539) );
	vdp_not g492 (.A(w536), .nZ(w535) );
	vdp_oai21 g493 (.A1(w571), .Z(w536), .A2(w567), .B(w537) );
	vdp_and3 g494 (.Z(w558), .B(w567), .A(w492), .C(w508) );
	vdp_nor g495 (.Z(w1402), .A(w557), .B(w508) );
	vdp_nor g496 (.Z(w565), .A(w505), .B(w504) );
	vdp_aoi21 g497 (.A1(DCLK1), .Z(w1394), .A2(w496), .B(w559) );
	vdp_comb1 g498 (.Z(w1401), .A1(w567), .B(w569), .A2(w1402), .C(HCLK1) );
	vdp_not g499 (.A(w545), .nZ(w33) );
	vdp_not g500 (.A(w1461), .nZ(w540) );
	vdp_not g501 (.A(VRAM128k), .nZ(w543) );
	vdp_not g502 (.A(w542), .nZ(w121) );
	vdp_not g503 (.A(w1462), .nZ(w122) );
	vdp_not g504 (.A(w1463), .nZ(w541) );
	vdp_not g505 (.A(VRAMA[0]), .nZ(w1464) );
	vdp_not g506 (.A(w549), .nZ(w548) );
	vdp_not g507 (.A(w486), .nZ(w593) );
	vdp_not g508 (.A(w493), .nZ(w595) );
	vdp_not g509 (.A(w570), .nZ(w592) );
	vdp_not g510 (.A(SEL0_M3), .nZ(w591) );
	vdp_not g511 (.A(VRAM128k), .nZ(w1468) );
	vdp_not g512 (.A(w508), .nZ(w587) );
	vdp_not g513 (.A(SYSRES), .nZ(w489) );
	vdp_not g514 (.A(FIFO_EMPTY), .nZ(w1396) );
	vdp_not g515 (.A(w32), .nZ(w1395) );
	vdp_not g516 (.A(w566), .nZ(w583) );
	vdp_not g517 (.A(w559), .nZ(w563) );
	vdp_not g518 (.A(w563), .nZ(w564) );
	vdp_sr_bit g519 (.D(w1397), .C2(HCLK2), .C1(HCLK1), .Q(w567), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g520 (.D(w1400), .Q(w571), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_slatch g521 (.Q(w447), .D(VRAMA[0]), .C(w583), .nC(w566) );
	vdp_and g522 (.A(w30), .Z(w1397), .B(w1396) );
	vdp_and g523 (.A(w1395), .Z(w487), .B(w3) );
	vdp_and g524 (.A(w3), .Z(w566), .B(HCLK1) );
	vdp_and g525 (.A(FIFO_EMPTY), .Z(w32), .B(w573) );
	vdp_and g526 (.A(w574), .Z(w34), .B(FIFO_EMPTY) );
	vdp_and g527 (.A(w574), .B(w558) );
	vdp_or g528 (.A(w562), .Z(w560), .B(w496) );
	vdp_or g529 (.A(w564), .Z(w913), .B(1'b0) );
	vdp_or g530 (.A(SYSRES), .Z(w585), .B(w578) );
	vdp_and g531 (.A(w567), .Z(w1398), .B(DMA_BUSY) );
	vdp_and g532 (.A(w596), .Z(w492), .B(w1467) );
	vdp_and g533 (.A(w1468), .Z(w1467), .B(SEL0_M3) );
	vdp_or g534 (.A(w558), .Z(w590), .B(w557) );
	vdp_or g535 (.A(DMA_BUSY), .Z(w1465), .B(w552) );
	vdp_or g536 (.A(DMA_BUSY), .Z(w1466), .B(w551) );
	vdp_and g537 (.A(M5), .Z(w570), .B(REG_BUS[0]) );
	vdp_or g538 (.A(w528), .Z(w544), .B(w543) );
	vdp_and g539 (.A(w533), .Z(w1460), .B(VRAM128k) );
	vdp_aon22 g540 (.Z(w518), .A2(w1465), .B1(w591), .B2(w570), .A1(SEL0_M3) );
	vdp_aon22 g541 (.Z(w524), .A2(w1466), .B1(w592), .B2(w591), .A1(SEL0_M3) );
	vdp_and3 g542 (.A(w30), .Z(w1400), .B(w34), .C(w1399) );
	vdp_rs_ff g543 (.Q(w1399), .R(w585), .S(w1398) );
	vdp_oai21 g544 (.A1(VRAMA[0]), .Z(w549), .A2(VRAM128k), .B(w577) );
	vdp_oai21 g545 (.A1(VRAM128k), .Z(w1463), .A2(w1464), .B(w577) );
	vdp_aoi21 g546 (.A1(w533), .Z(w1462), .A2(w546), .B(w548) );
	vdp_aoi21 g547 (.A1(w528), .Z(w542), .A2(w546), .B(w541) );
	vdp_aoi21 g548 (.A1(w546), .Z(w1461), .A2(w544), .B(w577) );
	vdp_aoi21 g549 (.A1(w546), .Z(w545), .A2(w1460), .B(w577) );
	vdp_and4 g550 (.A(w535), .Z(w546), .B(w539), .C(w534), .D(w538) );
	vdp_not g551 (.A(w621), .nZ(w1388) );
	vdp_not g552 (.A(w633), .nZ(w632) );
	vdp_and3 g553 (.A(w587), .Z(w588), .B(w623), .C(w632) );
	vdp_and3 g554 (.A(w595), .Z(w610), .B(w597), .C(w593) );
	vdp_and3 g555 (.A(w493), .Z(w614), .B(w597), .C(w593) );
	vdp_and3 g556 (.A(w595), .Z(w603), .B(w597), .C(w486) );
	vdp_and3 g557 (.A(w493), .Z(w607), .B(w597), .C(w486) );
	vdp_or g558 (.A(w589), .Z(w620), .B(w622) );
	vdp_or g559 (.A(w589), .Z(w626), .B(w630) );
	vdp_or g560 (.A(w654), .Z(w576), .B(w629) );
	vdp_and3 g561 (.Z(w574), .B(DMA_BUSY), .A(w653), .C(w628) );
	vdp_or3 g562 (.Z(w580), .B(w571), .A(w577), .C(w627) );
	vdp_and g563 (.A(w581), .Z(w496), .B(w582) );
	vdp_and g564 (.A(w567), .Z(w597), .B(w587) );
	vdp_bufif0 g565 (.A(w579), .Z(VRAMA[8]), .nE(w634) );
	vdp_aoi221 g566 (.Z(w621), .A2(w588), .B1(FIFO_EMPTY), .B2(w565), .A1(w565), .C(SYSRES) );
	vdp_aon33 g567 (.Z(FIFO_FULL), .A2(w565), .B1(w1498), .B2(w565), .A1(w631), .A3(w1498), .B3(w584) );
	vdp_not g568 (.A(w590), .nZ(w1416) );
	vdp_comp_str g569 (.A(w553), .Z(w1417), .nZ(w617) );
	vdp_not g570 (.A(w614), .nZ(w616) );
	vdp_comp_str g571 (.A(w455), .Z(w1419), .nZ(w1418) );
	vdp_not g572 (.A(w590), .nZ(w823) );
	vdp_comp_str g573 (.A(w553), .Z(w618), .nZ(w619) );
	vdp_not g574 (.A(w569), .nZ(w634) );
	vdp_not g575 (.A(w614), .nZ(w1499) );
	vdp_comp_str g576 (.A(w455), .Z(w1420), .nZ(w615) );
	vdp_not g577 (.A(w610), .nZ(w609) );
	vdp_comp_str g578 (.A(w446), .Z(w1421), .nZ(w1503) );
	vdp_not g579 (.A(w610), .nZ(w611) );
	vdp_comp_str g580 (.A(w495), .Z(w1422), .nZ(w608) );
	vdp_comp_str g581 (.A(w446), .Z(w612), .nZ(w613) );
	vdp_not g582 (.A(w603), .nZ(w600) );
	vdp_comp_str g583 (.A(w452), .Z(w601), .nZ(w602) );
	vdp_not g584 (.A(w603), .nZ(w822) );
	vdp_comp_str g585 (.A(w452), .Z(w1501), .nZ(w1502) );
	vdp_not g586 (.A(w607), .nZ(w604) );
	vdp_comp_str g587 (.A(w495), .Z(w605), .nZ(w606) );
	vdp_not g588 (.A(w607), .nZ(w1500) );
	vdp_sr_bit g589 (.D(w1388), .Q(FIFO_EMPTY), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g590 (.D(w623), .Q(w633), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g591 (.D(w567), .Q(w623), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g592 (.D(FIFO_FULL), .Q(w631), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g593 (.D(w560), .Q(w584), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_not g594 (.A(SYSRES), .nZ(w1498) );
	vdp_not g595 (.A(w1470), .nZ(w627) );
	vdp_sr_bit g596 (.D(w581), .Q(w582), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g597 (.D(w572), .C2(HCLK2), .C1(HCLK1), .Q(w578), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_dlatch_inv g598 (.D(w581), .C(HCLK2), .Q(w1470), .nC(nHCLK2) );
	vdp_slatch g599 (.D(w644), .C(w601), .nC(w602), .nQ(w6452) );
	vdp_slatch g600 (.D(REG_BUS[7]), .C(w1501), .nC(w1502), .nQ(w6453) );
	vdp_slatch g601 (.D(w644), .C(w605), .nC(w606), .nQ(w6472) );
	vdp_slatch g602 (.D(REG_BUS[7]), .C(w1422), .nC(w608), .nQ(w6470) );
	vdp_slatch g603 (.D(w644), .C(w1421), .nC(w1503), .nQ(w6486) );
	vdp_slatch g604 (.D(REG_BUS[7]), .C(w612), .nC(w613), .nQ(w6488) );
	vdp_slatch g605 (.D(w644), .C(w1420), .nC(w615), .nQ(w6506) );
	vdp_slatch g606 (.D(REG_BUS[7]), .C(w1419), .nC(w1418), .nQ(w6504) );
	vdp_slatch g607 (.D(VRAMA[9]), .C(w1417), .nC(w617), .nQ(w6520) );
	vdp_slatch g608 (.D(VRAMA[7]), .C(w618), .nC(w619), .nQ(w6521) );
	vdp_notif0 g609 (.nZ(VRAMA[7]), .nE(w823), .A(w6521) );
	vdp_notif0 g610 (.nZ(VRAMA[9]), .nE(w1416), .A(w6520) );
	vdp_notif0 g611 (.nZ(VRAMA[7]), .nE(w616), .A(w6504) );
	vdp_notif0 g612 (.nZ(VRAMA[9]), .nE(w1499), .A(w6506) );
	vdp_notif0 g613 (.nZ(VRAMA[7]), .nE(w611), .A(w6488) );
	vdp_notif0 g614 (.nZ(VRAMA[9]), .nE(w604), .A(w6472) );
	vdp_notif0 g615 (.nZ(VRAMA[7]), .nE(w1500), .A(w6470) );
	vdp_notif0 g616 (.nZ(VRAMA[9]), .nE(w609), .A(w6486) );
	vdp_notif0 g617 (.nZ(VRAMA[9]), .nE(w600), .A(w6452) );
	vdp_notif0 g618 (.nZ(VRAMA[7]), .nE(w822), .A(w6453) );
	vdp_bufif0 g619 (.A(w644), .Z(VRAMA[9]), .nE(w634) );
	vdp_bufif0 g620 (.A(REG_BUS[7]), .Z(VRAMA[7]), .nE(w634) );
	vdp_bufif0 g621 (.A(w637), .Z(VRAMA[8]), .nE(w1452) );
	vdp_bufif0 g622 (.A(w637), .Z(CA[8]), .nE(w825) );
	vdp_bufif0 g623 (.A(w636), .Z(VRAMA[7]), .nE(w1450) );
	vdp_bufif0 g624 (.A(w636), .Z(CA[7]), .nE(w824) );
	vdp_slatch g625 (.Q(w653), .D(REG_BUS[7]), .nQ(w651), .C(w1544), .nC(w1545) );
	vdp_not g626 (.A(REG_BUS[0]), .nZ(w649) );
	vdp_not g627 (.A(REG_BUS[7]), .nZ(w655) );
	vdp_and3 g628 (.Z(w654), .B(w628), .A(w651), .C(DMA_BUSY) );
	vdp_nand g629 (.A(w647), .Z(w675), .B(w648) );
	vdp_cnt_bit_load g630 (.D(REG_BUS[0]), .nL(w1547), .L(w1556), .R(1'b0), .Q(w637), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w620), .CO(w641) );
	vdp_cnt_bit_load g631 (.D(REG_BUS[7]), .nL(w1387), .L(w782), .R(1'b0), .Q(w636), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w639), .CO(w622) );
	vdp_cnt_bit_load g632 (.D(w649), .nL(w1546), .L(w791), .R(1'b0), .Q(w647), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w626), .CO(w646) );
	vdp_cnt_bit_load g633 (.D(w655), .nL(w772), .L(w773), .R(1'b0), .Q(w650), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w652), .CO(w630) );
	vdp_slatch g634 (.D(w663), .C(w601), .nC(w602), .nQ(w6451) );
	vdp_slatch g635 (.D(REG_BUS[6]), .C(w1501), .nC(w1502), .nQ(w6454) );
	vdp_slatch g636 (.D(w663), .C(w605), .nC(w606), .nQ(w6471) );
	vdp_slatch g637 (.D(REG_BUS[6]), .C(w1422), .nC(w608), .nQ(w6469) );
	vdp_slatch g638 (.D(w663), .C(w1421), .nC(w1503), .nQ(w6485) );
	vdp_slatch g639 (.D(REG_BUS[6]), .C(w612), .nC(w613), .nQ(w6487) );
	vdp_slatch g640 (.D(w663), .C(w1420), .nC(w615), .nQ(w6505) );
	vdp_slatch g641 (.D(REG_BUS[6]), .C(w1419), .nC(w1418), .nQ(w6503) );
	vdp_slatch g642 (.D(VRAMA[10]), .C(w1417), .nC(w617), .nQ(w6519) );
	vdp_slatch g643 (.D(VRAMA[6]), .C(w618), .nC(w619), .nQ(w6522) );
	vdp_notif0 g644 (.nZ(VRAMA[6]), .nE(w823), .A(w6522) );
	vdp_notif0 g645 (.nZ(VRAMA[10]), .nE(w1416), .A(w6519) );
	vdp_notif0 g646 (.nZ(VRAMA[6]), .nE(w616), .A(w6503) );
	vdp_notif0 g647 (.nZ(VRAMA[10]), .nE(w1499), .A(w6505) );
	vdp_notif0 g648 (.nZ(VRAMA[6]), .nE(w611), .A(w6487) );
	vdp_notif0 g649 (.nZ(VRAMA[10]), .nE(w604), .A(w6471) );
	vdp_notif0 g650 (.nZ(VRAMA[6]), .nE(w1500), .A(w6469) );
	vdp_notif0 g651 (.nZ(VRAMA[10]), .nE(w609), .A(w6485) );
	vdp_notif0 g652 (.nZ(VRAMA[10]), .nE(w600), .A(w6451) );
	vdp_notif0 g653 (.nZ(VRAMA[6]), .nE(w822), .A(w6454) );
	vdp_bufif0 g654 (.A(w663), .Z(VRAMA[10]), .nE(w634) );
	vdp_bufif0 g655 (.A(REG_BUS[6]), .Z(VRAMA[6]), .nE(w1453) );
	vdp_bufif0 g656 (.A(w635), .Z(VRAMA[9]), .nE(w1452) );
	vdp_bufif0 g657 (.A(w635), .Z(CA[9]), .nE(w825) );
	vdp_bufif0 g658 (.A(w657), .Z(VRAMA[6]), .nE(w1450) );
	vdp_bufif0 g659 (.A(w657), .Z(CA[6]), .nE(w824) );
	vdp_slatch g660 (.Q(w670), .D(REG_BUS[6]), .nQ(w628), .C(w1544), .nC(w1545) );
	vdp_not g661 (.A(REG_BUS[1]), .nZ(w666) );
	vdp_not g662 (.A(REG_BUS[6]), .nZ(w668) );
	vdp_and3 g663 (.Z(w629), .B(DMA_BUSY), .A(w670), .C(w651) );
	vdp_cnt_bit_load g664 (.D(REG_BUS[1]), .nL(w1547), .L(w1556), .R(1'b0), .Q(w635), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w641), .CO(w659) );
	vdp_cnt_bit_load g665 (.D(REG_BUS[6]), .nL(w1387), .L(w782), .R(1'b0), .Q(w657), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w658), .CO(w639) );
	vdp_cnt_bit_load g666 (.D(w666), .nL(w1546), .L(w791), .R(1'b0), .Q(w648), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w646), .CO(w665) );
	vdp_cnt_bit_load g667 (.D(w668), .nL(w772), .L(w773), .R(1'b0), .Q(w667), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w671), .CO(w652) );
	vdp_nand3 g668 (.Z(w674), .B(w667), .A(w673), .C(w650) );
	vdp_slatch g669 (.D(w686), .C(w601), .nC(w602), .nQ(w6450) );
	vdp_slatch g670 (.D(REG_BUS[5]), .C(w1501), .nC(w1502), .nQ(w6455) );
	vdp_slatch g671 (.D(w686), .C(w605), .nC(w606), .nQ(w6473) );
	vdp_slatch g672 (.D(REG_BUS[5]), .C(w1422), .nC(w608), .nQ(w6468) );
	vdp_slatch g673 (.D(w686), .C(w1421), .nC(w1503), .nQ(w6484) );
	vdp_slatch g674 (.D(w686), .C(w1420), .nC(w615), .nQ(w6507) );
	vdp_slatch g675 (.D(REG_BUS[5]), .C(w1419), .nC(w1418), .nQ(w6502) );
	vdp_slatch g676 (.D(VRAMA[11]), .C(w1417), .nC(w617), .nQ(w6518) );
	vdp_slatch g677 (.D(VRAMA[5]), .C(w618), .nC(w619), .nQ(w6523) );
	vdp_notif0 g678 (.nZ(VRAMA[5]), .nE(w823), .A(w6523) );
	vdp_notif0 g679 (.nZ(VRAMA[11]), .nE(w1416), .A(w6518) );
	vdp_notif0 g680 (.nZ(VRAMA[5]), .nE(w616), .A(w6502) );
	vdp_notif0 g681 (.nZ(VRAMA[11]), .nE(w1499), .A(w6507) );
	vdp_notif0 g682 (.nZ(VRAMA[5]), .nE(w611), .A(w6489) );
	vdp_notif0 g683 (.nZ(VRAMA[11]), .nE(w604), .A(w6473) );
	vdp_notif0 g684 (.nZ(VRAMA[5]), .nE(w1500), .A(w6468) );
	vdp_notif0 g685 (.nZ(VRAMA[11]), .nE(w609), .A(w6484) );
	vdp_notif0 g686 (.nZ(VRAMA[11]), .nE(w600), .A(w6450) );
	vdp_notif0 g687 (.nZ(VRAMA[5]), .nE(w822), .A(w6455) );
	vdp_bufif0 g688 (.A(w686), .Z(VRAMA[11]), .nE(w634) );
	vdp_bufif0 g689 (.A(REG_BUS[5]), .Z(VRAMA[5]), .nE(w1453) );
	vdp_bufif0 g690 (.A(w656), .Z(VRAMA[10]), .nE(w1452) );
	vdp_bufif0 g691 (.A(w656), .Z(CA[10]), .nE(w825) );
	vdp_bufif0 g692 (.A(w688), .Z(VRAMA[5]), .nE(w1450) );
	vdp_bufif0 g693 (.A(w688), .Z(CA[5]), .nE(w824) );
	vdp_slatch g694 (.Q(CA[18]), .D(REG_BUS[2]), .C(w1544), .nC(w1545) );
	vdp_not g695 (.A(REG_BUS[2]), .nZ(w681) );
	vdp_not g696 (.A(REG_BUS[5]), .nZ(w680) );
	vdp_and3 g697 (.Z(w573), .B(DMA_BUSY), .A(w670), .C(w653) );
	vdp_cnt_bit_load g698 (.D(REG_BUS[2]), .nL(w1547), .L(w1556), .R(1'b0), .Q(w656), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w659), .CO(w691) );
	vdp_cnt_bit_load g699 (.D(REG_BUS[5]), .nL(w1387), .L(w782), .R(1'b0), .Q(w688), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w687), .CO(w658) );
	vdp_cnt_bit_load g700 (.D(w681), .nL(w1546), .L(w791), .R(1'b0), .Q(w672), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w665), .CO(w682) );
	vdp_cnt_bit_load g701 (.D(w680), .nL(w772), .L(w773), .R(1'b0), .Q(w673), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w677), .CO(w671) );
	vdp_nand3 g702 (.Z(w685), .B(w683), .A(w684), .C(w672) );
	vdp_slatch g703 (.D(w699), .C(w601), .nC(w602), .nQ(w6449) );
	vdp_slatch g704 (.D(REG_BUS[4]), .C(w1501), .nC(w1502), .nQ(w6456) );
	vdp_slatch g705 (.D(w699), .C(w605), .nC(w606), .nQ(w6474) );
	vdp_slatch g706 (.D(REG_BUS[4]), .C(w1422), .nC(w608), .nQ(w6467) );
	vdp_slatch g707 (.D(w699), .C(w1421), .nC(w1503), .nQ(w6483) );
	vdp_slatch g708 (.D(w699), .C(w1420), .nC(w615), .nQ(w6508) );
	vdp_slatch g709 (.D(REG_BUS[4]), .C(w1419), .nC(w1418), .nQ(w6501) );
	vdp_slatch g710 (.D(VRAMA[12]), .C(w1417), .nC(w617), .nQ(w6517) );
	vdp_slatch g711 (.D(VRAMA[4]), .C(w618), .nC(w619), .nQ(w6524) );
	vdp_notif0 g712 (.nZ(VRAMA[4]), .nE(w823), .A(w6524) );
	vdp_notif0 g713 (.nZ(VRAMA[12]), .nE(w1416), .A(w6517) );
	vdp_notif0 g714 (.nZ(VRAMA[4]), .nE(w616), .A(w6501) );
	vdp_notif0 g715 (.nZ(VRAMA[12]), .nE(w1499), .A(w6508) );
	vdp_notif0 g716 (.nZ(VRAMA[4]), .nE(w611), .A(w6490) );
	vdp_notif0 g717 (.nZ(VRAMA[12]), .nE(w604), .A(w6474) );
	vdp_notif0 g718 (.nZ(VRAMA[4]), .nE(w1500), .A(w6467) );
	vdp_notif0 g719 (.nZ(VRAMA[12]), .nE(w609), .A(w6483) );
	vdp_notif0 g720 (.nZ(VRAMA[12]), .nE(w600), .A(w6449) );
	vdp_notif0 g721 (.nZ(VRAMA[4]), .nE(w822), .A(w6456) );
	vdp_bufif0 g722 (.A(w699), .Z(VRAMA[12]), .nE(w634) );
	vdp_bufif0 g723 (.A(REG_BUS[4]), .Z(VRAMA[4]), .nE(w1453) );
	vdp_bufif0 g724 (.A(w690), .Z(VRAMA[11]), .nE(w1452) );
	vdp_bufif0 g725 (.A(w690), .Z(CA[11]), .nE(w825) );
	vdp_bufif0 g726 (.A(w700), .Z(VRAMA[4]), .nE(w1450) );
	vdp_bufif0 g727 (.A(w700), .Z(CA[4]), .nE(w824) );
	vdp_slatch g728 (.Q(CA[19]), .D(REG_BUS[3]), .C(w1544), .nC(w1545) );
	vdp_not g729 (.A(REG_BUS[3]), .nZ(w701) );
	vdp_not g730 (.A(REG_BUS[4]), .nZ(w703) );
	vdp_and g731 (.Z(w572), .B(w679), .A(w711) );
	vdp_cnt_bit_load g732 (.D(REG_BUS[3]), .nL(w1547), .L(w1556), .R(1'b0), .Q(w690), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w691), .CO(w695) );
	vdp_cnt_bit_load g733 (.D(REG_BUS[4]), .nL(w1387), .L(w782), .R(1'b0), .Q(w700), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w705), .CO(w687) );
	vdp_cnt_bit_load g734 (.D(w701), .nL(w1546), .L(w791), .R(1'b0), .Q(w683), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w682), .CO(w706) );
	vdp_cnt_bit_load g735 (.D(w703), .nL(w772), .L(w773), .R(1'b0), .Q(w709), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w710), .CO(w677) );
	vdp_nor3 g736 (.Z(w679), .B(w685), .A(w708), .C(w675) );
	vdp_slatch g737 (.D(w716), .C(w601), .nC(w602), .nQ(w6448) );
	vdp_slatch g738 (.D(REG_BUS[3]), .C(w1501), .nC(w1502), .nQ(w6457) );
	vdp_slatch g739 (.D(w716), .C(w605), .nC(w606), .nQ(w6475) );
	vdp_slatch g740 (.D(REG_BUS[3]), .C(w1422), .nC(w608), .nQ(w6466) );
	vdp_slatch g741 (.D(w716), .C(w1421), .nC(w1503), .nQ(w6482) );
	vdp_slatch g742 (.D(REG_BUS[3]), .C(w612), .nC(w613), .nQ(w6492) );
	vdp_slatch g743 (.D(w716), .C(w1420), .nC(w615), .nQ(w6510) );
	vdp_slatch g744 (.D(REG_BUS[3]), .C(w1419), .nC(w1418), .nQ(w6500) );
	vdp_slatch g745 (.D(VRAMA[13]), .C(w1417), .nC(w617), .nQ(w6516) );
	vdp_slatch g746 (.D(VRAMA[3]), .C(w618), .nC(w619), .nQ(w6525) );
	vdp_notif0 g747 (.nZ(VRAMA[3]), .nE(w823), .A(w6525) );
	vdp_notif0 g748 (.nZ(VRAMA[13]), .nE(w1416), .A(w6516) );
	vdp_notif0 g749 (.nZ(VRAMA[3]), .nE(w616), .A(w6500) );
	vdp_notif0 g750 (.nZ(VRAMA[13]), .nE(w1499), .A(w6510) );
	vdp_notif0 g751 (.nZ(VRAMA[3]), .nE(w611), .A(w6492) );
	vdp_notif0 g752 (.nZ(VRAMA[13]), .nE(w604), .A(w6475) );
	vdp_notif0 g753 (.nZ(VRAMA[3]), .nE(w1500), .A(w6466) );
	vdp_notif0 g754 (.nZ(VRAMA[13]), .nE(w609), .A(w6482) );
	vdp_notif0 g755 (.nZ(VRAMA[13]), .nE(w600), .A(w6448) );
	vdp_notif0 g756 (.nZ(VRAMA[3]), .nE(w822), .A(w6457) );
	vdp_bufif0 g757 (.A(w716), .Z(VRAMA[13]), .nE(w634) );
	vdp_bufif0 g758 (.A(REG_BUS[3]), .Z(VRAMA[3]), .nE(w1453) );
	vdp_bufif0 g759 (.A(w694), .Z(VRAMA[12]), .nE(w1452) );
	vdp_bufif0 g760 (.A(w694), .Z(CA[12]), .nE(w825) );
	vdp_bufif0 g761 (.A(w724), .Z(VRAMA[3]), .nE(w1450) );
	vdp_bufif0 g762 (.A(w724), .Z(CA[3]), .nE(w824) );
	vdp_slatch g763 (.Q(w730), .D(REG_BUS[4]), .C(w1544), .nC(w1545) );
	vdp_not g764 (.A(REG_BUS[4]), .nZ(w718) );
	vdp_not g765 (.A(REG_BUS[3]), .nZ(w719) );
	vdp_cnt_bit_load g766 (.D(REG_BUS[4]), .nL(w1547), .L(w1556), .R(1'b0), .Q(w694), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w695), .CO(w715) );
	vdp_cnt_bit_load g767 (.D(REG_BUS[3]), .nL(w1387), .L(w782), .R(1'b0), .Q(w724), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w713), .CO(w705) );
	vdp_cnt_bit_load g768 (.D(w718), .nL(w1546), .L(w791), .R(1'b0), .Q(w684), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w706), .CO(w723) );
	vdp_cnt_bit_load g769 (.D(w719), .nL(w772), .L(w773), .R(1'b0), .Q(w728), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w720), .CO(w710) );
	vdp_nor3 g770 (.Z(w711), .B(w729), .A(w727), .C(w674) );
	vdp_bufif0 g771 (.A(w730), .Z(CA[20]), .nE(w770) );
	vdp_slatch g772 (.D(w734), .C(w601), .nC(w602), .nQ(w6447) );
	vdp_slatch g773 (.D(REG_BUS[2]), .C(w1501), .nC(w1502), .nQ(w6458) );
	vdp_slatch g774 (.D(w734), .C(w605), .nC(w606), .nQ(w6476) );
	vdp_slatch g775 (.D(REG_BUS[2]), .C(w1422), .nC(w608), .nQ(w6465) );
	vdp_slatch g776 (.D(w734), .C(w1421), .nC(w1503), .nQ(w6481) );
	vdp_slatch g777 (.D(REG_BUS[2]), .C(w612), .nC(w613), .nQ(w6491) );
	vdp_slatch g778 (.D(w734), .C(w1420), .nC(w615), .nQ(w6509) );
	vdp_slatch g779 (.D(REG_BUS[2]), .C(w1419), .nC(w1418), .nQ(w6499) );
	vdp_slatch g780 (.D(VRAMA[14]), .C(w1417), .nC(w617), .nQ(w6515) );
	vdp_slatch g781 (.D(VRAMA[2]), .nC(w619), .C(w618), .nQ(w6526) );
	vdp_notif0 g782 (.nZ(VRAMA[2]), .nE(w823), .A(w6526) );
	vdp_notif0 g783 (.nZ(VRAMA[14]), .nE(w1416), .A(w6515) );
	vdp_notif0 g784 (.nZ(VRAMA[2]), .nE(w616), .A(w6499) );
	vdp_notif0 g785 (.nZ(VRAMA[14]), .nE(w1499), .A(w6509) );
	vdp_notif0 g786 (.nZ(VRAMA[2]), .nE(w611), .A(w6491) );
	vdp_notif0 g787 (.nZ(VRAMA[14]), .nE(w604), .A(w6476) );
	vdp_notif0 g788 (.nZ(VRAMA[2]), .nE(w1500), .A(w6465) );
	vdp_notif0 g789 (.nZ(VRAMA[14]), .nE(w609), .A(w6481) );
	vdp_notif0 g790 (.nZ(VRAMA[14]), .nE(w600), .A(w6447) );
	vdp_notif0 g791 (.nZ(VRAMA[2]), .nE(w822), .A(w6458) );
	vdp_bufif0 g792 (.A(w734), .Z(VRAMA[14]), .nE(w1451) );
	vdp_bufif0 g793 (.A(REG_BUS[2]), .Z(VRAMA[2]), .nE(w1453) );
	vdp_bufif0 g794 (.A(w714), .Z(VRAMA[13]), .nE(w1452) );
	vdp_bufif0 g795 (.A(w714), .Z(CA[13]), .nE(w825) );
	vdp_bufif0 g796 (.A(w735), .Z(VRAMA[2]), .nE(w1450) );
	vdp_bufif0 g797 (.A(w735), .Z(CA[2]), .nE(w824) );
	vdp_slatch g798 (.Q(w740), .D(REG_BUS[5]), .C(w1544), .nC(w1545) );
	vdp_not g799 (.A(REG_BUS[5]), .nZ(w736) );
	vdp_not g800 (.A(REG_BUS[2]), .nZ(w737) );
	vdp_cnt_bit_load g801 (.D(REG_BUS[5]), .nL(w1547), .L(w1556), .R(1'b0), .Q(w714), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w715), .CO(w746) );
	vdp_cnt_bit_load g802 (.D(REG_BUS[2]), .nL(w1387), .L(w782), .R(1'b0), .Q(w735), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w745), .CO(w713) );
	vdp_cnt_bit_load g803 (.D(w736), .nL(w1546), .L(w791), .R(1'b0), .Q(w744), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w723), .CO(w738) );
	vdp_cnt_bit_load g804 (.D(w737), .nL(w772), .L(w773), .R(1'b0), .Q(w742), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w748), .CO(w720) );
	vdp_nand3 g805 (.Z(w729), .B(w728), .A(w742), .C(w709) );
	vdp_bufif0 g806 (.A(w740), .Z(CA[21]), .nE(w770) );
	vdp_slatch g807 (.D(w753), .C(w601), .nC(w602), .nQ(w6446) );
	vdp_slatch g808 (.D(REG_BUS[1]), .C(w1501), .nC(w1502), .nQ(w6459) );
	vdp_slatch g809 (.D(w753), .C(w605), .nC(w606), .nQ(w6478) );
	vdp_slatch g810 (.D(REG_BUS[1]), .C(w1422), .nC(w608), .nQ(w6464) );
	vdp_slatch g811 (.D(w753), .C(w1421), .nC(w1503), .nQ(w6480) );
	vdp_slatch g812 (.D(REG_BUS[1]), .C(w612), .nC(w613), .nQ(w6494) );
	vdp_slatch g813 (.D(w753), .C(w1420), .nC(w615), .nQ(w6511) );
	vdp_slatch g814 (.D(REG_BUS[1]), .C(w1419), .nC(w1418), .nQ(w6498) );
	vdp_slatch g815 (.D(VRAMA[15]), .C(w1417), .nC(w617), .nQ(w6514) );
	vdp_slatch g816 (.D(VRAMA[1]), .C(w618), .nC(w619), .nQ(w6527) );
	vdp_notif0 g817 (.nZ(VRAMA[1]), .nE(w823), .A(w6527) );
	vdp_notif0 g818 (.nZ(VRAMA[15]), .nE(w1416), .A(w6514) );
	vdp_notif0 g819 (.nZ(VRAMA[1]), .nE(w616), .A(w6498) );
	vdp_notif0 g820 (.nZ(VRAMA[15]), .nE(w1499), .A(w6511) );
	vdp_notif0 g821 (.nZ(VRAMA[1]), .nE(w611), .A(w6494) );
	vdp_notif0 g822 (.nZ(VRAMA[15]), .nE(w604), .A(w6478) );
	vdp_notif0 g823 (.nZ(VRAMA[1]), .nE(w1500), .A(w6464) );
	vdp_notif0 g824 (.nZ(VRAMA[15]), .nE(w609), .A(w6480) );
	vdp_notif0 g825 (.nZ(VRAMA[15]), .nE(w600), .A(w6446) );
	vdp_notif0 g826 (.nZ(VRAMA[1]), .nE(w822), .A(w6459) );
	vdp_bufif0 g827 (.A(w753), .Z(VRAMA[15]), .nE(w1451) );
	vdp_bufif0 g828 (.A(REG_BUS[1]), .Z(VRAMA[1]), .nE(w1453) );
	vdp_bufif0 g829 (.A(w731), .Z(VRAMA[14]), .nE(w1452) );
	vdp_bufif0 g830 (.A(w731), .Z(CA[14]), .nE(w825) );
	vdp_bufif0 g831 (.A(w755), .Z(VRAMA[1]), .nE(w1450) );
	vdp_bufif0 g832 (.A(w755), .Z(CA[1]), .nE(w824) );
	vdp_slatch g833 (.Q(w1454), .D(REG_BUS[1]), .C(w1544), .nC(w1545) );
	vdp_not g834 (.A(REG_BUS[6]), .nZ(w758) );
	vdp_not g835 (.A(REG_BUS[1]), .nZ(w761) );
	vdp_cnt_bit_load g836 (.D(REG_BUS[6]), .nL(w1547), .L(w1556), .R(1'b0), .Q(w731), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w746), .CO(w762) );
	vdp_cnt_bit_load g837 (.D(REG_BUS[1]), .nL(w1387), .L(w782), .R(1'b0), .Q(w755), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w763), .CO(w745) );
	vdp_cnt_bit_load g838 (.D(w758), .nL(w1546), .L(w791), .R(1'b0), .Q(w743), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w738), .CO(w756) );
	vdp_cnt_bit_load g839 (.D(w761), .nL(w772), .L(w773), .R(1'b0), .Q(w760), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w759), .CO(w748) );
	vdp_nand3 g840 (.Z(w708), .B(w743), .A(w744), .C(w757) );
	vdp_bufif0 g841 (.A(w1454), .Z(CA[17]), .nE(w770) );
	vdp_slatch g842 (.nQ(w754), .D(w767), .C(w601), .nC(w602) );
	vdp_slatch g843 (.D(REG_BUS[0]), .C(w1501), .nC(w1502), .nQ(w6460) );
	vdp_slatch g844 (.D(w767), .C(w605), .nC(w606), .nQ(w6477) );
	vdp_slatch g845 (.D(REG_BUS[0]), .C(w1422), .nC(w608), .nQ(w6463) );
	vdp_slatch g846 (.D(w767), .C(w1421), .nC(w1503), .nQ(w6479) );
	vdp_slatch g847 (.D(REG_BUS[0]), .C(w612), .nC(w613), .nQ(w6493) );
	vdp_slatch g848 (.D(w767), .C(w1420), .nC(w615), .nQ(w6512) );
	vdp_slatch g849 (.D(REG_BUS[0]), .C(w1419), .nC(w1418), .nQ(w6497) );
	vdp_slatch g850 (.D(VRAMA[16]), .C(w1417), .nC(w617), .nQ(w6513) );
	vdp_slatch g851 (.Q(w6528), .D(VRAMA[0]), .C(w618), .nC(w619) );
	vdp_notif0 g852 (.nZ(VRAMA[0]), .nE(w823), .A(w6528) );
	vdp_notif0 g853 (.nZ(VRAMA[16]), .nE(w1416), .A(w6513) );
	vdp_notif0 g854 (.nZ(VRAMA[0]), .nE(w616), .A(w6497) );
	vdp_notif0 g855 (.nZ(VRAMA[16]), .nE(w1499), .A(w6512) );
	vdp_notif0 g856 (.nZ(VRAMA[0]), .nE(w611), .A(w6493) );
	vdp_notif0 g857 (.nZ(VRAMA[16]), .nE(w604), .A(w6477) );
	vdp_notif0 g858 (.nZ(VRAMA[0]), .nE(w1500), .A(w6463) );
	vdp_notif0 g859 (.nZ(VRAMA[16]), .nE(w609), .A(w6479) );
	vdp_notif0 g860 (.A(w754), .nZ(VRAMA[16]), .nE(w600) );
	vdp_notif0 g861 (.nZ(VRAMA[0]), .nE(w822), .A(w6460) );
	vdp_bufif0 g862 (.A(w767), .Z(VRAMA[16]), .nE(w1451) );
	vdp_bufif0 g863 (.A(REG_BUS[0]), .Z(VRAMA[0]), .nE(w1453) );
	vdp_bufif0 g864 (.A(w749), .Z(VRAMA[15]), .nE(w1452) );
	vdp_bufif0 g865 (.A(w749), .Z(CA[15]), .nE(w825) );
	vdp_bufif0 g866 (.A(w777), .Z(VRAMA[0]), .nE(w1450) );
	vdp_bufif0 g867 (.A(w777), .Z(CA[0]), .nE(w824) );
	vdp_slatch g868 (.Q(w768), .D(REG_BUS[0]), .C(w1544), .nC(w1545) );
	vdp_not g869 (.A(REG_BUS[7]), .nZ(w1548) );
	vdp_not g870 (.A(REG_BUS[0]), .nZ(w1424) );
	vdp_cnt_bit_load g871 (.D(REG_BUS[7]), .nL(w1547), .L(w1556), .R(1'b0), .Q(w749), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w762) );
	vdp_cnt_bit_load g872 (.D(REG_BUS[0]), .nL(w1387), .L(w782), .R(1'b0), .Q(w777), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w775), .CO(w763) );
	vdp_cnt_bit_load g873 (.D(w1548), .nL(w1546), .L(w791), .R(1'b0), .Q(w757), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w756) );
	vdp_cnt_bit_load g874 (.D(w1424), .nL(w772), .L(w773), .R(1'b0), .Q(w1423), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w775), .CO(w759) );
	vdp_nand3 g875 (.Z(w727), .B(w760), .A(w580), .C(w1382) );
	vdp_bufif0 g876 (.A(w768), .Z(CA[16]), .nE(w770) );
	vdp_slatch g877 (.D(VRAMA[8]), .C(w618), .nC(w619), .nQ(w6529) );
	vdp_slatch g878 (.D(w579), .C(w1419), .nC(w1418), .nQ(w6496) );
	vdp_slatch g879 (.D(w579), .C(w612), .nC(w613), .nQ(w6495) );
	vdp_slatch g880 (.D(w579), .C(w1422), .nC(w608), .nQ(w6462) );
	vdp_slatch g881 (.D(w579), .C(w1501), .nC(w1502), .nQ(w6461) );
	vdp_notif0 g882 (.nZ(VRAMA[8]), .nE(w822), .A(w6461) );
	vdp_notif0 g883 (.nZ(VRAMA[8]), .nE(w1500), .A(w6462) );
	vdp_notif0 g884 (.nZ(VRAMA[8]), .nE(w611), .A(w6495) );
	vdp_notif0 g885 (.nZ(VRAMA[8]), .nE(w616), .A(w6496) );
	vdp_notif0 g886 (.nZ(VRAMA[8]), .nE(w823), .A(w6529) );
	vdp_bufif0 g887 (.A(w768), .Z(VRAMA[16]), .nE(w1452) );
	vdp_not g888 (.A(w1415), .nZ(w1451) );
	vdp_not g889 (.A(w569), .nZ(w1453) );
	vdp_not g890 (.A(w31), .nZ(w1452) );
	vdp_not g891 (.A(w576), .nZ(w825) );
	vdp_not g892 (.A(w31), .nZ(w1450) );
	vdp_not g893 (.A(w576), .nZ(w824) );
	vdp_not g894 (.A(w576), .nZ(w770) );
	vdp_not g895 (.A(w1423), .nZ(w1382) );
	vdp_not g896 (.A(w771), .nZ(w1386) );
	vdp_not g897 (.A(M5), .nZ(w787) );
	vdp_and4 g898 (.Z(w783), .B(w663), .A(w792), .D(w579), .C(w793) );
	vdp_and4 g899 (.Z(w784), .B(w663), .A(w792), .D(w795), .C(w644) );
	vdp_and4 g900 (.B(w796), .A(w778), .D(w795), .C(w793), .Z(w786) );
	vdp_and4 g901 (.B(w796), .A(w778), .D(w579), .C(w793), .Z(w785) );
	vdp_and4 g902 (.Z(w780), .B(w793), .A(w579), .D(w797), .C(w663) );
	vdp_and4 g903 (.Z(w788), .B(w644), .A(w795), .D(w778), .C(w796) );
	vdp_and4 g904 (.Z(w779), .B(w644), .A(w579), .D(w797), .C(w663) );
	vdp_and4 g905 (.B(w800), .A(M5), .D(w686), .C(w801), .Z(w792) );
	vdp_comp_str g906 (.A(w803), .Z(w1544), .nZ(w1545) );
	vdp_comp_we g907 (.A(w1428), .Z(w1556), .nZ(w1547) );
	vdp_comp_we g908 (.A(w781), .Z(w782), .nZ(w1387) );
	vdp_comp_we g909 (.A(w804), .Z(w791), .nZ(w1546) );
	vdp_comp_we g910 (.A(w805), .Z(w773), .nZ(w772) );
	vdp_and g911 (.Z(w589), .B(w580), .A(w771) );
	vdp_and g912 (.Z(w775), .B(w580), .A(w1386) );
	vdp_or g913 (.Z(w803), .B(w779), .A(SYSRES) );
	vdp_or g914 (.Z(w781), .B(w780), .A(SYSRES) );
	vdp_or g915 (.Z(w1415), .B(w787), .A(w569) );
	vdp_or g916 (.B(w785), .A(SYSRES), .Z(w171) );
	vdp_or g917 (.B(w786), .A(SYSRES), .Z(w170) );
	vdp_or g918 (.Z(w169), .B(w784), .A(SYSRES) );
	vdp_or g919 (.Z(w168), .B(w783), .A(SYSRES) );
	vdp_or g920 (.B(w1425), .A(SYSRES), .Z(w164) );
	vdp_and4 g921 (.B(w663), .A(w794), .D(w579), .C(w644), .Z(w810) );
	vdp_or g922 (.B(w810), .A(SYSRES), .Z(w163) );
	vdp_and4 g923 (.B(w796), .A(w797), .D(w795), .C(w644), .Z(w809) );
	vdp_or g924 (.B(w809), .A(SYSRES), .Z(w162) );
	vdp_and4 g925 (.B(w796), .A(w797), .D(w579), .C(w793), .Z(w808) );
	vdp_or g926 (.B(w808), .A(SYSRES), .Z(w161) );
	vdp_and4 g927 (.B(w796), .A(w797), .D(w795), .C(w793), .Z(w1426) );
	vdp_or g928 (.B(w1426), .A(SYSRES), .Z(w167) );
	vdp_and4 g929 (.B(w663), .A(w794), .D(w795), .C(w644), .Z(w807) );
	vdp_or g930 (.B(w807), .A(SYSRES), .Z(w160) );
	vdp_and4 g931 (.B(w663), .A(w794), .D(w579), .C(w793), .Z(w806) );
	vdp_or g932 (.B(w806), .A(SYSRES), .Z(w159) );
	vdp_or g933 (.B(w811), .A(SYSRES), .Z(w165) );
	vdp_and4 g934 (.B(w663), .A(w794), .D(w795), .C(w793), .Z(w1425) );
	vdp_or g935 (.B(w812), .A(SYSRES), .Z(w166) );
	vdp_and4 g936 (.B(w796), .A(w794), .D(w579), .C(w644), .Z(w811) );
	vdp_and4 g937 (.B(w796), .A(w794), .D(w795), .C(w644), .Z(w812) );
	vdp_and4 g938 (.B(w793), .A(w579), .D(w794), .C(w796), .Z(w814) );
	vdp_or g939 (.B(w814), .A(SYSRES), .Z(w1100) );
	vdp_and4 g940 (.B(w793), .A(w795), .D(w794), .C(w796), .Z(w1427) );
	vdp_or g941 (.B(w1427), .A(SYSRES), .Z(w1138) );
	vdp_and4 g942 (.B(w793), .A(w795), .D(w792), .C(w663), .Z(w813) );
	vdp_or g943 (.B(w813), .A(SYSRES), .Z(w1101) );
	vdp_and4 g944 (.B(w644), .A(w795), .D(w797), .C(w663), .Z(w815) );
	vdp_or g945 (.B(w815), .A(SYSRES), .Z(w1428) );
	vdp_and4 g946 (.B(w644), .A(w579), .D(w792), .C(w796), .Z(w1429) );
	vdp_or g947 (.B(w1429), .A(SYSRES), .Z(w1062) );
	vdp_and4 g948 (.B(w793), .A(w795), .D(w797), .C(w663), .Z(w816) );
	vdp_or g949 (.B(w816), .A(SYSRES), .Z(w804) );
	vdp_and4 g950 (.B(w644), .A(w579), .D(w797), .C(w796), .Z(w817) );
	vdp_or g951 (.B(w817), .A(SYSRES), .Z(w805) );
	vdp_and4 g952 (.B(w644), .A(w579), .D(w792), .C(w663), .Z(w818) );
	vdp_or g953 (.B(w818), .A(SYSRES), .Z(w819) );
	vdp_and4 g954 (.B(w802), .A(w800), .D(M5), .C(w699), .Z(w797) );
	vdp_and3 g955 (.B(w801), .A(w800), .C(w686), .Z(w778) );
	vdp_and3 g956 (.B(w802), .A(w800), .C(w801), .Z(w794) );
	vdp_or g957 (.Z(w820), .B(w821), .A(w6431) );
	vdp_and g958 (.B(w799), .A(HCLK1), .Z(w800) );
	vdp_dlatch_inv g959 (.D(w798), .C(DCLK2), .nQ(w821), .nC(nDCLK2) );
	vdp_dlatch_inv g960 (.D(w6430), .C(HCLK2), .nQ(w799), .nC(nHCLK2) );
	vdp_not g961 (.A(w699), .nZ(w801) );
	vdp_not g962 (.A(w686), .nZ(w802) );
	vdp_not g963 (.A(w644), .nZ(w793) );
	vdp_not g964 (.A(w663), .nZ(w796) );
	vdp_not g965 (.A(w579), .nZ(w795) );
	vdp_slatch g966 (.D(REG_BUS[5]), .C(w612), .nC(w613), .nQ(w6489) );
	vdp_slatch g967 (.D(REG_BUS[4]), .C(w612), .nC(w613), .nQ(w6490) );
	vdp_sr_bit g968 (.D(w821), .C2(DCLK2), .C1(DCLK1), .Q(w6431), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_dlatch_inv g969 (.D(w820), .C(DCLK1), .nQ(w6430), .nC(nDCLK1) );
	vdp_comp_str g970 (.A(w857), .Z(w827), .nZ(w835) );
	vdp_fa g971 (.SUM(w854), .A(REG_BUS[6]), .B(w1521), .CO(w856), .CI(w852) );
	vdp_fa g972 (.SUM(w850), .A(REG_BUS[5]), .B(w851), .CO(w852), .CI(w849) );
	vdp_fa g973 (.SUM(w847), .A(REG_BUS[4]), .B(w848), .CO(w849), .CI(w844) );
	vdp_fa g974 (.SUM(w843), .A(REG_BUS[3]), .B(w846), .CO(w844), .CI(w841) );
	vdp_fa g975 (.SUM(w839), .A(REG_BUS[2]), .B(w840), .CO(w841), .CI(w838) );
	vdp_fa g976 (.SUM(w6434), .A(REG_BUS[1]), .B(w837), .CO(w838), .CI(w834) );
	vdp_fa g977 (.SUM(w6435), .A(REG_BUS[0]), .B(w831), .CO(w834), .CI(w829) );
	vdp_fa g978 (.SUM(w1430), .A(REG_BUS[7]), .B(w1520), .CO(w858), .CI(w856) );
	vdp_slatch g979 (.Q(w855), .D(DB[7]), .C(w827), .nC(w835) );
	vdp_aon22 g980 (.Z(w1531), .A1(w855), .A2(w826), .B1(w832), .B2(w1430) );
	vdp_slatch g981 (.Q(w853), .D(DB[6]), .C(w827), .nC(w835) );
	vdp_aon22 g982 (.Z(w1532), .A1(w853), .A2(w826), .B1(w832), .B2(w854) );
	vdp_slatch g983 (.Q(w1473), .D(DB[5]), .C(w827), .nC(w835) );
	vdp_aon22 g984 (.Z(w1533), .A1(w1473), .A2(w826), .B1(w832), .B2(w850) );
	vdp_slatch g985 (.Q(w845), .D(DB[4]), .C(w827), .nC(w835) );
	vdp_aon22 g986 (.Z(w1534), .A1(w845), .A2(w826), .B1(w832), .B2(w847) );
	vdp_slatch g987 (.Q(w842), .D(DB[3]), .C(w827), .nC(w835) );
	vdp_aon22 g988 (.Z(w1535), .A1(w842), .A2(w826), .B1(w832), .B2(w843) );
	vdp_slatch g989 (.Q(w836), .D(DB[2]), .C(w827), .nC(w835) );
	vdp_aon22 g990 (.Z(w1536), .A1(w836), .A2(w826), .B1(w832), .B2(w839) );
	vdp_slatch g991 (.Q(w833), .D(DB[1]), .C(w827), .nC(w835) );
	vdp_aon22 g992 (.Z(w1537), .A1(w833), .A2(w826), .B1(w832), .B2(w6434) );
	vdp_slatch g993 (.Q(w828), .D(DB[0]), .C(w827), .nC(w835) );
	vdp_aon22 g994 (.Z(w1538), .A1(w828), .A2(w826), .B1(w832), .B2(w6435) );
	vdp_dff g995 (.Q(REG_BUS[0]), .R(SYSRES), .C(w860), .D(w1538) );
	vdp_slatch g996 (.Q(w831), .D(REG_BUS[0]), .C(w859), .nC(w830) );
	vdp_dff g997 (.Q(REG_BUS[1]), .R(SYSRES), .D(w1537), .C(w860) );
	vdp_slatch g998 (.Q(w837), .D(REG_BUS[1]), .C(w859), .nC(w830) );
	vdp_dff g999 (.Q(REG_BUS[2]), .R(SYSRES), .C(w860), .D(w1536) );
	vdp_slatch g1000 (.Q(w840), .D(REG_BUS[2]), .C(w859), .nC(w830) );
	vdp_dff g1001 (.Q(REG_BUS[3]), .R(SYSRES), .D(w1535), .C(w860) );
	vdp_slatch g1002 (.Q(w846), .D(REG_BUS[3]), .C(w859), .nC(w830) );
	vdp_dff g1003 (.Q(REG_BUS[4]), .R(SYSRES), .C(w860), .D(w1534) );
	vdp_slatch g1004 (.Q(w848), .D(REG_BUS[4]), .C(w859), .nC(w830) );
	vdp_dff g1005 (.Q(REG_BUS[5]), .R(SYSRES), .C(w860), .D(w1533) );
	vdp_slatch g1006 (.Q(w851), .D(REG_BUS[5]), .C(w859), .nC(w830) );
	vdp_dff g1007 (.Q(REG_BUS[6]), .R(SYSRES), .C(w860), .D(w1532) );
	vdp_slatch g1008 (.Q(w1521), .D(REG_BUS[6]), .C(w859), .nC(w830) );
	vdp_dff g1009 (.Q(REG_BUS[7]), .R(SYSRES), .D(w1531), .C(w860) );
	vdp_slatch g1010 (.Q(w1520), .D(REG_BUS[7]), .C(w859), .nC(w830) );
	vdp_comp_str g1011 (.A(w819), .Z(w859), .nZ(w830) );
	vdp_comp_we g1012 (.A(w861), .Z(w826), .nZ(w832) );
	vdp_dff g1013 (.Q(w767), .R(w865), .C(w860), .D(w1522) );
	vdp_dff g1014 (.Q(w753), .R(w865), .C(w860), .D(w1523) );
	vdp_dff g1015 (.Q(w734), .R(w865), .C(w860), .D(w1524) );
	vdp_dff g1016 (.Q(w716), .R(SYSRES), .C(w860), .D(w1525) );
	vdp_dff g1017 (.Q(w699), .R(SYSRES), .C(w860), .D(w1526) );
	vdp_dff g1018 (.Q(w686), .R(SYSRES), .C(w860), .D(w1527) );
	vdp_dff g1019 (.Q(w663), .R(SYSRES), .C(w860), .D(w1528) );
	vdp_dff g1020 (.Q(w644), .R(SYSRES), .C(w860), .D(w1529) );
	vdp_dff g1021 (.Q(w579), .R(SYSRES), .C(w860), .D(w1530) );
	vdp_not g1022 (.A(w887), .nZ(w860) );
	vdp_or g1023 (.Z(w865), .B(SYSRES), .A(w829) );
	vdp_not g1024 (.A(M5), .nZ(w829) );
	vdp_slatch g1025 (.Q(w884), .D(w278), .C(w897), .nC(w875) );
	vdp_aon22 g1026 (.Z(w1530), .A1(w888), .A2(w895), .B1(w862), .B2(w886) );
	vdp_slatch g1027 (.Q(w888), .D(w243), .C(w897), .nC(w875) );
	vdp_comp_str g1028 (.A(w901), .Z(w897), .nZ(w875) );
	vdp_comp_we g1029 (.A(w861), .Z(w895), .nZ(w862) );
	vdp_ha g1030 (.SUM(w886), .A(w579), .B(w858), .CO(w883) );
	vdp_slatch g1031 (.Q(w882), .D(w251), .C(w897), .nC(w875) );
	vdp_aon22 g1032 (.Z(w1529), .A1(w884), .A2(w895), .B1(w862), .B2(w885) );
	vdp_ha g1033 (.SUM(w885), .A(w644), .B(w883), .CO(w1541) );
	vdp_slatch g1034 (.Q(w880), .D(w287), .C(w897), .nC(w875) );
	vdp_aon22 g1035 (.Z(w1528), .A1(w882), .A2(w895), .B1(w862), .B2(w881) );
	vdp_ha g1036 (.SUM(w881), .A(w663), .B(w1541), .CO(w879) );
	vdp_slatch g1037 (.Q(w877), .D(w260), .C(w897), .nC(w875) );
	vdp_aon22 g1038 (.Z(w1527), .A1(w880), .A2(w895), .B1(w862), .B2(w878) );
	vdp_ha g1039 (.SUM(w878), .A(w686), .B(w879), .CO(w1540) );
	vdp_slatch g1040 (.Q(w874), .D(w296), .C(w897), .nC(w875) );
	vdp_aon22 g1041 (.Z(w1526), .A1(w877), .A2(w895), .B1(w862), .B2(w876) );
	vdp_ha g1042 (.SUM(w876), .A(w699), .B(w1540), .CO(w873) );
	vdp_aon22 g1043 (.Z(w1525), .A1(w874), .A2(w895), .B1(w862), .B2(w871) );
	vdp_ha g1044 (.SUM(w871), .A(w716), .B(w873), .CO(w872) );
	vdp_comp_str g1045 (.A(w896), .Z(w894), .nZ(w864) );
	vdp_aon22 g1046 (.Z(w1524), .A1(w870), .A2(w895), .B1(w862), .B2(w1539) );
	vdp_ha g1047 (.SUM(w1539), .A(w734), .B(w872), .CO(w867) );
	vdp_slatch_r g1048 (.Q(w870), .D(DB[0]), .R(w865), .C(w894), .nC(w864) );
	vdp_slatch_r g1049 (.Q(w869), .D(DB[1]), .R(w865), .C(w894), .nC(w864) );
	vdp_aon22 g1050 (.Z(w1523), .A1(w869), .A2(w895), .B1(w862), .B2(w868) );
	vdp_ha g1051 (.SUM(w868), .A(w753), .B(w867), .CO(w866) );
	vdp_slatch_r g1052 (.Q(w863), .D(DB[2]), .R(w865), .C(w894), .nC(w864) );
	vdp_aon22 g1053 (.Z(w1522), .A1(w863), .A2(w895), .B1(w862), .B2(w1472) );
	vdp_ha g1054 (.SUM(w1472), .A(w767), .B(w866) );
	vdp_and3 g1055 (.C(w891), .A(w889), .B(w890), .Z(w893) );
	vdp_sr_bit g1056 (.D(w1436), .C2(HCLK2), .C1(HCLK1), .nQ(w98), .nC1(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1057 (.D(w909), .Q(w1436), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK2), .nC1(nHCLK1) );
	vdp_not g1058 (.A(w935), .nZ(w911) );
	vdp_not g1059 (.A(w457), .nZ(w1437) );
	vdp_not g1060 (.A(w458), .nZ(w922) );
	vdp_not g1061 (.A(w889), .nZ(w923) );
	vdp_not g1062 (.A(w920), .nZ(w928) );
	vdp_not g1063 (.A(w498), .nZ(w906) );
	vdp_not g1064 (.A(w573), .nZ(w917) );
	vdp_not g1065 (.A(w942), .nZ(w931) );
	vdp_not g1066 (.A(w1438), .nZ(w934) );
	vdp_not g1067 (.A(w932), .nZ(w902) );
	vdp_slatch g1068 (.Q(w484), .D(w899), .C(w900), .nC(w912) );
	vdp_slatch g1069 (.Q(w498), .D(w269), .C(w900), .nC(w912) );
	vdp_comp_str g1070 (.A(w901), .Z(w900), .nZ(w912) );
	vdp_dlatch_inv g1071 (.D(w581), .C(DCLK1), .nQ(w932), .nC(nDCLK1) );
	vdp_dlatch_inv g1072 (.D(w931), .C(DCLK1), .nQ(w930), .nC(nDCLK1) );
	vdp_dlatch_inv g1073 (.D(w944), .C(DCLK2), .nQ(w942), .nC(nDCLK2) );
	vdp_dlatch_inv g1074 (.D(w949), .C(DCLK1), .nQ(w944), .nC(nDCLK1) );
	vdp_slatch g1075 (.Q(w949), .D(w908), .C(DCLK2), .nC(nDCLK2) );
	vdp_slatch g1076 (.Q(w908), .D(w943), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g1077 (.D(w569), .C(HCLK1), .nQ(w907), .nC(nHCLK1) );
	vdp_rs_ff g1078 (.nQ(w904), .R(w951), .S(w950), .Q(w915) );
	vdp_rs_ff g1079 (.Q(w927), .R(w925), .S(w905) );
	vdp_and3 g1080 (.C(w412), .A(w458), .B(w1437), .Z(w910) );
	vdp_and3 g1081 (.C(w922), .A(w457), .B(w412), .Z(w97) );
	vdp_comp_dff g1082 (.D(w926), .C2(HCLK2), .C1(HCLK1), .Q(w919), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_comp_dff g1083 (.D(w916), .C2(HCLK2), .C1(HCLK1), .Q(w918), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g1084 (.C(w30), .A(w915), .B(FIFO_EMPTY), .Z(w916) );
	vdp_and g1085 (.A(DB[7]), .B(w896), .Z(w898) );
	vdp_and g1086 (.A(w907), .B(w949), .Z(w861) );
	vdp_and g1087 (.A(w918), .B(w917), .Z(w557) );
	vdp_and g1088 (.A(w573), .B(w918), .Z(w577) );
	vdp_and g1089 (.A(w919), .B(w917), .Z(w929) );
	vdp_and g1090 (.A(w573), .B(w919), .Z(w31) );
	vdp_or g1091 (.A(w919), .B(w940), .Z(w925) );
	vdp_or g1092 (.A(w919), .B(w557), .Z(w412) );
	vdp_or g1093 (.A(w573), .B(w440), .Z(w948) );
	vdp_aoi21 g1094 (.A1(w930), .B(SYSRES), .Z(w1438), .A2(w931) );
	vdp_or3 g1095 (.C(w903), .A(w924), .B(w893), .Z(w905) );
	vdp_or3 g1096 (.C(w577), .A(w929), .B(w571), .Z(w569) );
	vdp_or5 g1097 (.C(w913), .A(w902), .B(w569), .Z(w887), .D(w901), .E(w896) );
	vdp_nand3 g1098 (.C(w892), .A(w928), .B(w938), .Z(w798) );
	vdp_2a3oi g1099 (.A1(w891), .B(w945), .Z(w939), .A2(w938), .C(w890) );
	vdp_nand g1100 (.A(w484), .B(w906), .Z(w920) );
	vdp_nor g1101 (.A(w908), .B(w944), .Z(w892) );
	vdp_and4 g1102 (.C(w904), .A(FIFO_EMPTY), .B(w30), .Z(w926), .D(w927) );
	vdp_nor5 g1103 (.C(w498), .A(w952), .B(w939), .Z(w903), .D(w484), .E(w923) );
	vdp_and g1104 (.A(w573), .B(w952), .Z(w924) );
	vdp_not g1105 (.A(w562), .nZ(w1490) );
	vdp_not g1106 (.A(w1490), .nZ(w986) );
	vdp_not g1107 (.A(w967), .nZ(w1003) );
	vdp_not g1108 (.A(w944), .nZ(w1443) );
	vdp_not g1109 (.A(w949), .nZ(w988) );
	vdp_not g1110 (.A(w991), .nZ(w901) );
	vdp_not g1111 (.A(SEL0_M3), .nZ(w921) );
	vdp_not g1112 (.A(w976), .nZ(w984) );
	vdp_not g1113 (.A(M5), .nZ(w891) );
	vdp_rs_ff g1114 (.Q(w938), .R(w936), .S(w901) );
	vdp_rs_ff g1115 (.Q(w890), .R(w936), .S(w1011) );
	vdp_rs_ff g1116 (.Q(w945), .R(w936), .S(w896) );
	vdp_rs_ff g1117 (.nQ(w947), .R(w946), .S(w914) );
	vdp_rs_ff g1118 (.Q(w1008), .R(w934), .S(w941) );
	vdp_rs_ff g1119 (.Q(w552), .R(w934), .S(w1001) );
	vdp_rs_ff g1120 (.Q(w551), .R(w934), .S(w958) );
	vdp_or g1121 (.A(w958), .B(w1001), .Z(w1010) );
	vdp_and g1122 (.A(w1008), .B(w889), .Z(w559) );
	vdp_and g1123 (.A(w1007), .B(w1008), .Z(w562) );
	vdp_and g1124 (.A(w988), .B(w1443), .Z(w889) );
	vdp_and g1125 (.A(w988), .B(w942), .Z(w1007) );
	vdp_and g1126 (.A(w944), .B(w942), .Z(w974) );
	vdp_and g1127 (.A(w919), .B(w948), .Z(w950) );
	vdp_and g1128 (.A(w970), .B(w959), .Z(w403) );
	vdp_and g1129 (.A(w921), .B(w857), .Z(w1017) );
	vdp_and g1130 (.A(w994), .B(w993), .Z(w941) );
	vdp_or g1131 (.A(w918), .B(w940), .Z(w951) );
	vdp_or g1132 (.A(w987), .B(w990), .Z(w933) );
	vdp_or g1133 (.A(SYSRES), .B(w889), .Z(w946) );
	vdp_or g1134 (.A(SYSRES), .B(w949), .Z(w1014) );
	vdp_or g1135 (.A(w944), .B(w943), .Z(w1009) );
	vdp_or g1136 (.A(w970), .B(w994), .Z(w1015) );
	vdp_or g1137 (.A(w937), .B(SYSRES), .Z(w980) );
	vdp_or g1138 (.A(SYSRES), .B(w975), .Z(w1019) );
	vdp_or g1139 (.A(SYSRES), .B(w974), .Z(w936) );
	vdp_and g1140 (.A(w935), .B(w910), .Z(w119) );
	vdp_and g1141 (.A(w910), .B(w911), .Z(w96) );
	vdp_and g1142 (.A(w889), .B(w982), .Z(w1018) );
	vdp_nand g1143 (.A(w403), .B(w947), .Z(w999) );
	vdp_nor g1144 (.A(FIFO_FULL), .B(w986), .Z(w1000) );
	vdp_or5 g1145 (.C(w901), .A(w985), .B(w998), .Z(w997), .D(w857), .E(w1002) );
	vdp_or3 g1146 (.C(w989), .A(w970), .B(w398), .Z(w990) );
	vdp_nor g1147 (.A(w97), .B(w910), .Z(w909) );
	vdp_and3 g1148 (.C(w1020), .A(w1016), .B(w972), .Z(w992) );
	vdp_or4 g1149 (.C(w941), .A(w896), .B(w969), .Z(w937), .D(w403) );
	vdp_and4 g1150 (.C(w1016), .A(w994), .B(w977), .Z(w857), .D(w995) );
	vdp_aoi21 g1151 (.A1(w889), .B(SYSRES), .Z(w976), .A2(w983) );
	vdp_aoi21 g1152 (.A1(w857), .B(w992), .Z(w991), .A2(SEL0_M3) );
	vdp_or5 g1153 (.C(w403), .A(w969), .B(w896), .Z(w975), .D(w941), .E(w901) );
	vdp_and5 g1154 (.C(w981), .A(M5), .B(w1016), .Z(w896), .D(w995), .E(w994) );
	vdp_not g1155 (.A(CA[7]), .nZ(w963) );
	vdp_not g1156 (.A(w994), .nZ(w971) );
	vdp_not g1157 (.A(w971), .nZ(w956) );
	vdp_not g1158 (.A(w970), .nZ(w955) );
	vdp_not g1159 (.A(w955), .nZ(w954) );
	vdp_slatch g1160 (.Q(w996), .D(w957), .nC(w954), .C(w955) );
	vdp_slatch g1161 (.Q(w1016), .D(w957), .nC(w956), .C(w971), .nQ(w993) );
	vdp_rs_ff g1162 (.Q(w978), .R(w974), .S(w980) );
	vdp_rs_ff g1163 (.Q(w982), .R(w1019), .S(w1017), .nQ(w983) );
	vdp_rs_ff g1164 (.Q(w1020), .R(w984), .S(w1018), .nQ(w995) );
	vdp_rs_ff g1165 (.Q(w981), .R(w979), .S(w1434), .nQ(w977) );
	vdp_slatch_r g1166 (.Q(w952), .D(DB[6]), .C(w973), .nC(w953), .R(w865) );
	vdp_slatch_r g1167 (.Q(w458), .D(DB[5]), .R(w865), .C(w973), .nC(w953) );
	vdp_slatch_r g1168 (.Q(w457), .D(DB[4]), .R(w865), .C(w973), .nC(w953) );
	vdp_comp_str g1169 (.A(w896), .Z(w973), .nZ(w953) );
	vdp_not g1170 (.A(w1435), .nZ(w979) );
	vdp_aoi21 g1171 (.A1(w889), .B(SYSRES), .Z(w1435), .A2(w978) );
	vdp_and4 g1172 (.C(w920), .A(M5), .B(w938), .Z(w1434), .D(w889) );
	vdp_and g1173 (.A(w970), .B(w996), .Z(w1011) );
	vdp_rs_ff g1174 (.nQ(w1013), .R(w1012), .S(w1011) );
	vdp_rs_ff g1175 (.Q(w943), .R(w1014), .S(w1015) );
	vdp_not g1176 (.A(w957), .nZ(w1542) );
	vdp_not g1177 (.A(CA[2]), .nZ(w1043) );
	vdp_not g1178 (.A(CA[3]), .nZ(w1044) );
	vdp_aon22 g1179 (.Z(w957), .A1(CA[0]), .A2(w1069), .B1(SEL0_M3), .B2(CA[1]) );
	vdp_and4 g1180 (.C(w962), .A(w963), .B(CA[6]), .Z(w1006), .D(w961) );
	vdp_and4 g1181 (.C(w966), .A(w965), .B(CA[7]), .Z(w972), .D(w961) );
	vdp_and4 g1182 (.C(CA[3]), .A(w1003), .B(w1005), .Z(w989), .D(CA[9]) );
	vdp_and4 g1183 (.C(CA[2]), .A(w1003), .B(w1005), .Z(w394), .D(w1044) );
	vdp_and4 g1184 (.C(w967), .A(w1043), .B(CA[3]), .Z(w964), .D(w1005) );
	vdp_or g1185 (.A(w1006), .B(w394), .Z(w398) );
	vdp_and g1186 (.A(w941), .B(w1000), .Z(w998) );
	vdp_and g1187 (.A(w990), .B(w999), .Z(w1002) );
	vdp_and g1188 (.A(SEL0_M3), .B(w997), .Z(w1034) );
	vdp_or g1189 (.A(SYSRES), .B(w914), .Z(w1012) );
	vdp_or g1190 (.A(w972), .B(w960), .Z(w994) );
	vdp_or g1191 (.A(SYSRES), .B(w578), .Z(w940) );
	vdp_and3 g1192 (.C(w1042), .A(w896), .B(w1013), .Z(w985) );
	vdp_and3 g1193 (.C(w1045), .A(w1009), .B(w1170), .Z(w1005) );
	vdp_and5 g1194 (.C(CA[2]), .A(w967), .B(CA[3]), .Z(w1039), .D(w1542), .E(w1005) );
	vdp_and5 g1195 (.C(CA[2]), .A(w967), .B(w957), .Z(w1038), .D(CA[3]), .E(w1005) );
	vdp_and5 g1196 (.C(w1043), .A(w1010), .B(w1003), .Z(w968), .D(w1044), .E(w1005) );
	vdp_and5 g1197 (.C(w1044), .A(w1043), .B(w1010), .Z(w960), .D(w967), .E(w1005) );
	vdp_nor5 g1198 (.C(w1035), .A(w1038), .B(w1039), .Z(w1021), .D(w964), .E(w1034) );
	vdp_aon22 g1199 (.Z(w1032), .A1(w4), .A2(w1041), .B1(w37), .B2(SEL0_M3) );
	vdp_aon22 g1200 (.Z(VPOS_80), .A1(LSM0), .A2(VPOS[8]), .B1(w1029), .B2(VPOS[0]) );
	vdp_not g1201 (.A(LSM0), .nZ(w1029) );
	vdp_not g1202 (.A(SEL0_M3), .nZ(w1025) );
	vdp_not g1203 (.A(SEL0_M3), .nZ(w1041) );
	vdp_not g1204 (.A(w1487), .nZ(w101) );
	vdp_not g1205 (.A(CA[6]), .nZ(w965) );
	vdp_not g1206 (.A(w1432), .nZ(w1030) );
	vdp_not g1207 (.A(w957), .nZ(w959) );
	vdp_aoi21 g1208 (.A1(w958), .B(w1433), .Z(w1432), .A2(w964) );
	vdp_and4 g1209 (.C(w962), .A(w965), .B(CA[7]), .Z(w1431), .D(w961) );
	vdp_and4 g1210 (.C(w966), .A(w963), .B(CA[6]), .Z(w1433), .D(w961) );
	vdp_slatch g1211 (.Q(w103), .D(w962), .C(w1543), .nC(w1488) );
	vdp_comp_we g1212 (.A(PSG_Z80_CLK), .Z(w1543), .nZ(w1488) );
	vdp_and g1213 (.A(w47), .B(w1036), .Z(w1489) );
	vdp_and g1214 (.A(w957), .B(w970), .Z(w969) );
	vdp_or g1215 (.A(w968), .B(w1431), .Z(w970) );
	vdp_or g1216 (.A(w1035), .B(w1489), .Z(w1037) );
	vdp_or g1217 (.Z(w1031), .A(w38), .B(SYSRES) );
	vdp_and g1218 (.Z(V_INT_HAPPENED), .A(w58), .B(w1032) );
	vdp_rs_ff g1219 (.Q(w1027), .R(w1031), .S(V_INT_HAPPENED) );
	vdp_aoi221 g1220 (.Z(w1487), .A1(w100), .A2(1'b0), .B1(w1033), .B2(w1037), .C(w102) );
	vdp_aoi22 g1221 (.Z(w1022), .A1(w1028), .A2(w1025), .B1(SEL0_M3), .B2(w1027) );
	vdp_comp_str g1222 (.Z(w1055), .A(w58), .nZ(w1056) );
	vdp_comp_str g1223 (.Z(w1081), .A(w1062), .nZ(w1082) );
	vdp_comp_str g1224 (.Z(w1093), .A(w1101), .nZ(w1094) );
	vdp_comp_str g1225 (.Z(w1090), .A(w1100), .nZ(w1089) );
	vdp_not g1226 (.A(w1099), .nZ(w1102) );
	vdp_not g1227 (.A(w1091), .nZ(w1104) );
	vdp_not g1228 (.A(w1088), .nZ(w1103) );
	vdp_not g1229 (.A(w1103), .nZ(w1068) );
	vdp_not g1230 (.A(SEL0_M3), .nZ(w1069) );
	vdp_not g1231 (.A(w1104), .nZ(w1087) );
	vdp_not g1232 (.A(w1106), .nZ(w1086) );
	vdp_not g1233 (.A(w1105), .nZ(w1085) );
	vdp_aon222 g1234 (.C2(w1085), .B2(w1086), .A2(w1087), .C1(w1066), .B1(CA[15]), .A1(CA[7]), .Z(w1072) );
	vdp_aon222 g1235 (.C2(w1085), .B2(w1086), .A2(w1087), .C1(w1065), .B1(CA[13]), .A1(CA[6]), .Z(w1084) );
	vdp_aon222 g1236 (.C2(w1085), .B2(w1086), .A2(w1087), .C1(w1064), .B1(CA[12]), .A1(CA[5]), .Z(w1073) );
	vdp_aon222 g1237 (.C2(w1085), .B2(w1086), .A2(w1087), .C1(w1063), .B1(CA[11]), .A1(CA[4]), .Z(w1074) );
	vdp_aon222 g1238 (.C2(w1085), .B2(w1086), .A2(w1087), .C1(w1067), .B1(CA[10]), .A1(CA[3]), .Z(w1075) );
	vdp_aon222 g1239 (.C2(w1085), .B2(w1086), .A2(w1087), .C1(w1471), .B1(CA[9]), .A1(CA[2]), .Z(w1076) );
	vdp_aon222 g1240 (.C2(w1085), .B2(w1086), .A2(w1087), .C1(w1070), .B1(CA[8]), .A1(CA[1]), .Z(w1083) );
	vdp_aon222 g1241 (.C2(w1085), .B2(w1086), .A2(w1087), .C1(w1059), .B1(CA[14]), .A1(CA[0]), .Z(w1077) );
	vdp_aon222 g1242 (.C2(w1085), .B2(w1086), .A2(w1087), .C1(nHCLK1), .B1(1'b1), .A1(1'b0), .Z(w1088) );
	vdp_slatch g1243 (.Q(LSM0), .D(LSM0), .C(w1055), .nC(w1056) );
	vdp_slatch g1244 (.Q(LSM1), .D(LSM1), .C(w1055), .nC(w1056) );
	vdp_aon22 g1245 (.Z(w1058), .A1(COL[6]), .A2(w1095), .B1(w117), .B2(w1441) );
	vdp_not g1246 (.A(M2), .nZ(w1052) );
	vdp_not g1247 (.A(w1095), .nZ(w1441) );
	vdp_and g1248 (.Z(w1), .A(LSM1), .B(LSM0) );
	vdp_and g1249 (.Z(w1053), .A(M5), .B(w1052) );
	vdp_and g1250 (.Z(w1442), .A(M5), .B(M2) );
	vdp_and g1251 (.Z(VRAM128k), .A(M5), .B(w1079) );
	vdp_or3 g1252 (.Z(w1099), .A(w1096), .B(w1097), .C(w1349) );
	vdp_and g1253 (.Z(w1098), .A(w1096), .B(w1068) );
	vdp_nand g1254 (.Z(w1106), .A(w1104), .B(w1099) );
	vdp_nand g1255 (.Z(w1105), .A(w1104), .B(w1102) );
	vdp_slatch g1256 (.Q(LSCR), .D(REG_BUS[0]), .C(w1081), .nC(w1082) );
	vdp_slatch g1257 (.Q(HSCR), .D(REG_BUS[1]), .C(w1081), .nC(w1082) );
	vdp_slatch g1258 (.Q(VSCR), .D(REG_BUS[2]), .C(w1081), .nC(w1082) );
	vdp_slatch g1259 (.Q(IE2), .D(REG_BUS[3]), .C(w1081), .nC(w1082) );
	vdp_slatch g1260 (.Q(w116), .D(REG_BUS[4]), .C(w1081), .nC(w1082) );
	vdp_slatch g1261 (.Q(w82), .D(REG_BUS[5]), .C(w1081), .nC(w1082) );
	vdp_slatch g1262 (.Q(w1036), .D(REG_BUS[6]), .C(w1081), .nC(w1082) );
	vdp_slatch g1263 (.Q(w1091), .D(REG_BUS[7]), .C(w1081), .nC(w1082) );
	vdp_slatch g1264 (.Q(M2), .D(REG_BUS[3]), .C(w1090), .nC(w1089) );
	vdp_slatch g1265 (.Q(w1079), .D(REG_BUS[7]), .C(w1090), .nC(w1089) );
	vdp_slatch g1266 (.Q(w18), .D(REG_BUS[4]), .C(w1093), .nC(w1094) );
	vdp_slatch g1267 (.Q(S_TE), .D(REG_BUS[3]), .C(w1093), .nC(w1094) );
	vdp_slatch g1268 (.Q(LSM1), .D(REG_BUS[2]), .C(w1093), .nC(w1094) );
	vdp_slatch g1269 (.Q(LSM0), .D(REG_BUS[1]), .C(w1093), .nC(w1094) );
	vdp_slatch g1270 (.Q(H40), .D(REG_BUS[0]), .C(w1093), .nC(w1094) );
	vdp_slatch g1271 (.Q(w45), .D(REG_BUS[0]), .C(w1090), .nC(w1089) );
	vdp_slatch g1272 (.Q(w120), .D(REG_BUS[1]), .C(w1090), .nC(w1089) );
	vdp_slatch g1273 (.Q(M5), .D(REG_BUS[2]), .C(w1090), .nC(w1089) );
	vdp_slatch g1274 (.Q(M1), .D(REG_BUS[4]), .C(w1090), .nC(w1089) );
	vdp_slatch g1275 (.Q(IE0), .D(REG_BUS[5]), .C(w1090), .nC(w1089) );
	vdp_slatch g1276 (.Q(DISP), .D(REG_BUS[6]), .C(w1090), .nC(w1089) );
	vdp_and g1277 (.Z(w110), .A(w1038), .B(w1118) );
	vdp_and g1278 (.Z(w109), .A(w989), .B(w1118) );
	vdp_and g1279 (.Z(w111), .A(w1038), .B(w1119) );
	vdp_and g1280 (.Z(w112), .A(w989), .B(w1119) );
	vdp_and g1281 (.Z(w105), .A(w1038), .B(w1113) );
	vdp_and g1282 (.Z(w115), .A(w989), .B(w1113) );
	vdp_and g1283 (.Z(w57), .A(w1038), .B(w1114) );
	vdp_and g1284 (.Z(w48), .A(w989), .B(w1114) );
	vdp_and g1285 (.Z(w78), .A(w1038), .B(w1116) );
	vdp_and g1286 (.Z(w76), .A(w989), .B(w1116) );
	vdp_and g1287 (.Z(w80), .A(w1038), .B(w1117) );
	vdp_and g1288 (.Z(PSG_TEST_OE), .A(w989), .B(w1117) );
	vdp_and g1289 (.Z(w1134), .A(w1038), .B(w1121) );
	vdp_and g1290 (.Z(w1110), .A(w1038), .B(w1122) );
	vdp_and g1291 (.Z(w56), .A(w1038), .B(w1115) );
	vdp_and g1292 (.Z(w54), .A(w989), .B(w1115) );
	vdp_dlatch g1293 (.D(COL[0]), .C(HCLK1), .Q(w1059), .nC(nHCLK1) );
	vdp_dlatch g1294 (.D(COL[1]), .Q(w1070), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch g1295 (.D(COL[2]), .Q(w1471), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch g1296 (.D(COL[3]), .Q(w1067), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch g1297 (.D(COL[4]), .Q(w1063), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch g1298 (.D(COL[5]), .Q(w1064), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch g1299 (.D(w1058), .Q(w1065), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch g1300 (.D(COL[7]), .Q(w1066), .C(HCLK1), .nC(nHCLK1) );
	vdp_slatch g1301 (.Q(w52), .D(REG_BUS[5]), .C(w1094), .nC(w1093) );
	vdp_slatch g1302 (.Q(w39), .D(REG_BUS[6]), .C(w1094), .nC(w1093) );
	vdp_slatch g1303 (.Q(RS0), .D(REG_BUS[7]), .C(w1094), .nC(w1093) );
	vdp_slatch g1304 (.Q(w22), .D(REG_BUS[3]), .nC(w1141), .C(w1139) );
	vdp_slatch g1305 (.Q(w85), .D(REG_BUS[2]), .nC(w1141), .C(w1139) );
	vdp_slatch g1306 (.Q(M3), .D(REG_BUS[1]), .nC(w1141), .C(w1139) );
	vdp_slatch g1307 (.Q(w53), .D(REG_BUS[0]), .nC(w1141), .C(w1139) );
	vdp_slatch g1308 (.Q(w83), .D(REG_BUS[7]), .nC(w1141), .C(w1139) );
	vdp_slatch g1309 (.Q(w84), .D(REG_BUS[6]), .nC(w1141), .C(w1139) );
	vdp_slatch g1310 (.Q(w59), .D(REG_BUS[5]), .nC(w1141), .C(w1139) );
	vdp_slatch g1311 (.Q(w1380), .D(REG_BUS[4]), .nC(w1141), .C(w1139) );
	vdp_slatch_r g1312 (.Q(w106), .D(DB[14]), .nC(w1133), .R(w1128), .C(w1137) );
	vdp_slatch_r g1313 (.Q(w114), .D(DB[13]), .R(w1128), .nC(w1133), .C(w1137) );
	vdp_slatch_r g1314 (.Q(w107), .D(DB[12]), .R(w1128), .nC(w1133), .C(w1137) );
	vdp_comp_str g1315 (.Z(w1139), .A(w1138), .nZ(w1141) );
	vdp_comp_str g1316 (.Z(w1136), .A(w1110), .nZ(w1135) );
	vdp_not g1317 (.A(REG_BUS[6]), .nZ(w1439) );
	vdp_not g1318 (.A(REG_BUS[7]), .nZ(w1154) );
	vdp_not g1319 (.A(REG_BUS[4]), .nZ(w1142) );
	vdp_not g1320 (.A(REG_BUS[5]), .nZ(w1140) );
	vdp_not g1321 (.A(REG_BUS[2]), .nZ(w1155) );
	vdp_not g1322 (.A(REG_BUS[3]), .nZ(w1143) );
	vdp_not g1323 (.A(REG_BUS[0]), .nZ(w1149) );
	vdp_not g1324 (.A(REG_BUS[1]), .nZ(w1150) );
	vdp_not g1325 (.A(w1126), .nZ(w1145) );
	vdp_not g1326 (.A(w1127), .nZ(w1131) );
	vdp_not g1327 (.A(w1120), .nZ(w1144) );
	vdp_not g1328 (.A(w1132), .nZ(w1146) );
	vdp_comp_str g1329 (.Z(w1130), .nZ(w1129), .A(w1039) );
	vdp_slatch_r g1330 (.Q(w1132), .R(w1128), .D(DB[11]), .nC(w1129), .C(w1130) );
	vdp_slatch_r g1331 (.Q(w1120), .D(DB[10]), .nC(w1129), .R(w1128), .C(w1130) );
	vdp_and4 g1332 (.Z(w1448), .A(w1126), .B(w1127), .C(w1132), .D(w1120) );
	vdp_and4 g1333 (.Z(w1113), .A(w1132), .B(w1144), .C(w1131), .D(w1145) );
	vdp_and4 g1334 (.Z(w1119), .A(w1146), .B(w1120), .C(w1127), .D(w1126) );
	vdp_and4 g1335 (.Z(w1118), .A(w1146), .B(w1120), .C(w1127), .D(w1145) );
	vdp_and4 g1336 (.Z(w1117), .A(w1146), .B(w1120), .C(w1131), .D(w1126) );
	vdp_and4 g1337 (.Z(w1116), .A(w1146), .B(w1120), .C(w1131), .D(w1145) );
	vdp_and4 g1338 (.Z(w1114), .A(w1146), .B(w1144), .C(w1127), .D(w1126) );
	vdp_and4 g1339 (.Z(w1115), .A(w1146), .B(w1144), .C(w1127), .D(w1145) );
	vdp_and4 g1340 (.Z(w1122), .A(w1146), .B(w1144), .C(w1131), .D(w1126) );
	vdp_and4 g1341 (.Z(w1121), .A(w1146), .B(w1144), .C(w1131), .D(w1145) );
	vdp_nand g1342 (.Z(w1385), .A(w1448), .B(w1038) );
	vdp_slatch_r g1343 (.Q(w1126), .D(DB[8]), .R(w1128), .C(w1130), .nC(w1129) );
	vdp_slatch_r g1344 (.Q(w1125), .D(DB[11]), .R(w1128), .C(w1137), .nC(w1133) );
	vdp_slatch_r g1345 (.nC(w1129), .Q(w1127), .D(DB[9]), .R(w1128), .C(w1130) );
	vdp_slatch_r g1346 (.Q(w1124), .D(DB[10]), .R(w1128), .C(w1137), .nC(w1133) );
	vdp_slatch_r g1347 (.Q(w87), .D(DB[8]), .R(w1128), .C(w1137), .nC(w1133) );
	vdp_slatch_r g1348 (.Q(w1123), .D(DB[9]), .R(w1128), .C(w1137), .nC(w1133) );
	vdp_slatch_r g1349 (.Q(w86), .D(DB[7]), .R(w1128), .C(w1137), .nC(w1133) );
	vdp_slatch_r g1350 (.Q(w88), .D(DB[5]), .R(w1128), .C(w1137), .nC(w1133) );
	vdp_slatch_r g1351 (.Q(w89), .D(DB[6]), .R(w1128), .C(w1137), .nC(w1133) );
	vdp_slatch_r g1352 (.Q(w935), .D(DB[4]), .R(w1128), .C(w1137), .nC(w1133) );
	vdp_slatch_r g1353 (.Q(w1152), .D(DB[2]), .R(w1128), .C(w1137), .nC(w1133) );
	vdp_slatch_r g1354 (.Q(w1153), .D(DB[3]), .R(w1128), .C(w1137), .nC(w1133) );
	vdp_slatch_r g1355 (.Q(w1095), .D(DB[0]), .R(w1128), .C(w1137), .nC(w1133) );
	vdp_slatch_r g1356 (.Q(w771), .D(DB[1]), .R(w1128), .C(w1137), .nC(w1133) );
	vdp_slatch_r g1357 (.Q(w93), .D(DB[9]), .R(w1128), .C(w1136), .nC(w1135) );
	vdp_slatch_r g1358 (.Q(w94), .D(DB[10]), .R(w1128), .C(w1136), .nC(w1135) );
	vdp_slatch_r g1359 (.Q(w91), .D(DB[7]), .R(w1128), .C(w1136), .nC(w1135) );
	vdp_slatch_r g1360 (.Q(w92), .D(DB[8]), .R(w1128), .C(w1136), .nC(w1135) );
	vdp_slatch_r g1361 (.Q(w51), .D(DB[5]), .R(w1128), .C(w1136), .nC(w1135) );
	vdp_slatch_r g1362 (.Q(w41), .D(DB[6]), .R(w1128), .C(w1136), .nC(w1135) );
	vdp_slatch_r g1363 (.Q(w40), .D(DB[3]), .R(w1128), .C(w1136), .nC(w1135) );
	vdp_slatch_r g1364 (.Q(w42), .D(DB[4]), .R(w1128), .C(w1136), .nC(w1135) );
	vdp_slatch_r g1365 (.Q(w1440), .D(DB[1]), .R(w1128), .C(w1136), .nC(w1135) );
	vdp_slatch_r g1366 (.Q(w55), .D(DB[2]), .R(w1128), .C(w1136), .nC(w1135) );
	vdp_slatch_r g1367 (.Q(w43), .D(DB[0]), .R(w1128), .C(w1136), .nC(w1135) );
	vdp_comp_str g1368 (.Z(w1137), .nZ(w1133), .A(w1134) );
	vdp_notif0 g1369 (.A(VPOS[9]), .nZ(DB[10]), .nE(w1147) );
	vdp_notif0 g1370 (.A(VPOS[8]), .nZ(DB[9]), .nE(w1147) );
	vdp_bufif0 g1371 (.A(FIFO_EMPTY), .Z(DB[9]), .nE(w1178) );
	vdp_bufif0 g1372 (.A(FIFO_FULL), .Z(DB[8]), .nE(w1178) );
	vdp_bufif0 g1373 (.A(w1177), .Z(DB[1]), .nE(w1178) );
	vdp_bufif0 g1374 (.A(w1179), .Z(DB[0]), .nE(w1178) );
	vdp_bufif0 g1375 (.A(w1160), .Z(DB[7]), .nE(w1178) );
	vdp_bufif0 g1376 (.A(w1159), .Z(DB[6]), .nE(w1178) );
	vdp_bufif0 g1377 (.A(w1158), .Z(DB[5]), .nE(w1178) );
	vdp_bufif0 g1378 (.A(ODD_EVEN), .Z(DB[4]), .nE(w1178) );
	vdp_bufif0 g1379 (.A(w46), .Z(DB[3]), .nE(w1178) );
	vdp_bufif0 g1380 (.A(w20), .Z(DB[2]), .nE(w1178) );
	vdp_slatch_r g1381 (.Q(w72), .D(DB[4]), .R(w1128), .C(w1130), .nC(w1129) );
	vdp_slatch_r g1382 (.Q(w73), .D(DB[5]), .R(w1128), .C(w1130), .nC(w1129) );
	vdp_slatch_r g1383 (.Q(w75), .D(DB[7]), .R(w1128), .C(w1130), .nC(w1129) );
	vdp_slatch_r g1384 (.Q(w74), .D(DB[6]), .R(w1128), .C(w1130), .nC(w1129) );
	vdp_slatch_r g1385 (.Q(w68), .D(DB[0]), .R(w1128), .C(w1130), .nC(w1129) );
	vdp_slatch_r g1386 (.Q(w69), .D(DB[1]), .R(w1128), .C(w1130), .nC(w1129) );
	vdp_slatch_r g1387 (.Q(w71), .D(DB[3]), .R(w1128), .C(w1130), .nC(w1129) );
	vdp_slatch_r g1388 (.Q(w70), .D(DB[2]), .R(w1128), .C(w1130), .nC(w1129) );
	vdp_notif0 g1389 (.A(HPOS[0]), .nZ(DB[8]), .nE(w1147) );
	vdp_not g1390 (.A(SEL0_M3), .nZ(w1449) );
	vdp_comp_str g1391 (.Z(w1148), .A(w788), .nZ(w1151) );
	vdp_slatch_r g1392 (.Q(w1164), .D(w1149), .R(SYSRES), .C(w1148), .nC(w1151) );
	vdp_slatch_r g1393 (.Q(w1174), .D(w1155), .R(SYSRES), .C(w1148), .nC(w1151) );
	vdp_slatch_r g1394 (.Q(w1180), .D(w1150), .R(SYSRES), .C(w1148), .nC(w1151) );
	vdp_slatch_r g1395 (.Q(w1168), .D(w1439), .R(SYSRES), .C(w1148), .nC(w1151) );
	vdp_slatch_r g1396 (.Q(w1175), .D(w1143), .R(SYSRES), .C(w1148), .nC(w1151) );
	vdp_slatch_r g1397 (.Q(w1167), .D(w1140), .R(SYSRES), .C(w1148), .nC(w1151) );
	vdp_slatch_r g1398 (.Q(w1176), .D(w1142), .R(SYSRES), .C(w1148), .nC(w1151) );
	vdp_slatch_r g1399 (.Q(w1169), .D(w1154), .R(SYSRES), .C(w1148), .nC(w1151) );
	vdp_aon22 g1400 (.Z(w1177), .A1(FIFO_EMPTY), .A2(w1162), .B1(w1163), .B2(DMA_BUSY) );
	vdp_aon22 g1401 (.Z(w1179), .A1(FIFO_FULL), .A2(w1162), .B1(w1163), .B2(PAL) );
	vdp_and3 g1402 (.C(w1152), .A(w398), .B(w1449), .Z(w1157) );
	vdp_not g1403 (.A(w1157), .nZ(w1147) );
	vdp_not g1404 (.A(w969), .nZ(w1178) );
	vdp_cnt_bit_load g1405 (.V(w1169), .nL(w1184), .L(w1165), .R(1'b0), .Q(w1185), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1212) );
	vdp_cnt_bit_load g1406 (.V(w1168), .nL(w1184), .L(w1165), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1481), .CO(w1212) );
	vdp_cnt_bit_load g1407 (.V(w1167), .nL(w1184), .L(w1165), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1211), .CO(w1481) );
	vdp_cnt_bit_load g1408 (.V(w1176), .nL(w1184), .L(w1165), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1210), .CO(w1211) );
	vdp_cnt_bit_load g1409 (.V(w1175), .nL(w1184), .L(w1165), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1209), .CO(w1210) );
	vdp_cnt_bit_load g1410 (.V(w1174), .nL(w1184), .L(w1165), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1491), .CO(w1209) );
	vdp_cnt_bit_load g1411 (.V(w1180), .nL(w1184), .L(w1165), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1208), .CO(w1491) );
	vdp_cnt_bit_load g1412 (.V(w1164), .nL(w1184), .L(w1165), .R(1'b0), .CI(w1182), .CO(w1208), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g1413 (.D(w1445), .C2(HCLK2), .C1(HCLK1), .Q(w1186), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_rs_ff g1414 (.Q(w1159), .R(w1202), .S(w1203) );
	vdp_rs_ff g1415 (.Q(w1160), .R(w1201), .S(V_INT_HAPPENED) );
	vdp_rs_ff g1416 (.Q(w1158), .R(w1202), .S(COLLISION) );
	vdp_not g1417 (.A(M5), .nZ(w1200) );
	vdp_not g1418 (.A(w1160), .nZ(w1181) );
	vdp_not g1419 (.A(w1166), .nZ(w1171) );
	vdp_not g1420 (.A(CA[21]), .nZ(w1446) );
	vdp_not g1421 (.A(SEL0_M3), .nZ(w1172) );
	vdp_not g1422 (.A(w1205), .nZ(w1173) );
	vdp_comp_we g1423 (.Z(w1184), .A(w1444), .nZ(w1165) );
	vdp_or g1424 (.A(w1205), .B(w1186), .Z(w1444) );
	vdp_and g1425 (.A(w1173), .B(w1185), .Z(w1445) );
	vdp_and g1426 (.A(w1181), .B(SPRITE_OVF), .Z(w1203) );
	vdp_or g1427 (.A(w1153), .B(w4), .Z(w1182) );
	vdp_not g1428 (.A(w1162), .nZ(w1163) );
	vdp_nor3 g1429 (.A(SEL0_M3), .B(w1200), .Z(w1162), .C(CA[1]) );
	vdp_nor3 g1430 (.A(w1153), .B(w5), .Z(w1205), .C(w29) );
	vdp_nor g1431 (.A(w1207), .B(w1187), .Z(w1170) );
	vdp_or5 g1432 (.A(w1172), .B(CA[4]), .C(CA[5]), .D(CA[15]), .Z(w1207), .E(CA[6]) );
	vdp_or5 g1433 (.A(CA[16]), .B(CA[17]), .C(CA[20]), .D(w1171), .Z(w1187), .E(w1446) );
	vdp_rs_ff g1434 (.Q(w1193), .R(w1244), .S(w1445) );
	vdp_rs_ff g1435 (.Q(w1245), .R(w1228), .S(w1447) );
	vdp_dff g1436 (.Q(w1247), .R(w1206), .C(w1196), .D(w1189) );
	vdp_dff g1437 (.Q(w1246), .R(w1206), .C(w1196), .D(w1188) );
	vdp_dff g1438 (.Q(w1248), .R(w1206), .C(w1196), .D(w1190) );
	vdp_rs_ff g1439 (.Q(w1497), .R(w1243), .S(w1496) );
	vdp_rs_ff g1440 (.Q(w1216), .R(w1217), .S(w1494) );
	vdp_dlatch_inv g1441 (.D(w1223), .Q(w1224), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g1442 (.D(w1217), .C(DCLK1), .Q(w1223), .nC(nDCLK1) );
	vdp_dlatch_inv g1443 (.D(w1226), .Q(w1202), .C(HCLK1), .nC(nHCLK1) );
	vdp_not g1444 (.A(w1239), .nZ(w1213) );
	vdp_not g1445 (.A(w653), .nZ(w1192) );
	vdp_not g1446 (.A(w1195), .nZ(w1190) );
	vdp_not g1447 (.A(w1194), .nZ(w1189) );
	vdp_not g1448 (.A(w1204), .nZ(w1206) );
	vdp_not g1449 (.A(w1220), .nZ(w1196) );
	vdp_not g1450 (.A(w1197), .nZ(w50) );
	vdp_not g1451 (.A(w1198), .nZ(w1199) );
	vdp_sr_bit g1452 (.D(w1225), .C2(HCLK2), .C1(HCLK1), .Q(w1243), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and g1453 (.A(M5), .B(w1216), .Z(w1220) );
	vdp_and g1454 (.A(SEL0_M3), .B(w1215), .Z(w1045) );
	vdp_and g1455 (.A(w1197), .B(w1045), .Z(w1495) );
	vdp_or g1456 (.A(w987), .B(w1495), .Z(w1494) );
	vdp_or g1457 (.A(w969), .B(SYSRES), .Z(w1496) );
	vdp_and g1458 (.A(w1200), .B(w1202), .Z(w1227) );
	vdp_or g1459 (.A(w1246), .B(w1227), .Z(w1228) );
	vdp_and g1460 (.A(M5), .B(w460), .Z(w1447) );
	vdp_and g1461 (.A(M1), .B(M5), .Z(w1191) );
	vdp_or g1462 (.A(w1248), .B(w1227), .Z(w1201) );
	vdp_or g1463 (.A(w1247), .B(w1227), .Z(w1244) );
	vdp_comp_dff g1464 (.D(w1497), .C2(HCLK2), .C1(HCLK1), .Q(w1225), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_comp_dff g1465 (.D(w1220), .C2(DCLK2), .C1(DCLK1), .Q(w1217), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_nor g1466 (.A(w1225), .B(SYSRES), .Z(w1519) );
	vdp_nand g1467 (.A(w1243), .B(w1519), .Z(w1226) );
	vdp_nand g1468 (.A(w1160), .B(IE0), .Z(w1195) );
	vdp_and3 g1469 (.A(w1191), .B(w898), .Z(w1238), .C(w1192) );
	vdp_and3 g1470 (.A(w1191), .B(w898), .Z(w1237), .C(w653) );
	vdp_and4 g1471 (.A(w1194), .B(IE2), .C(w1195), .D(w1245), .Z(w1188) );
	vdp_nand3 g1472 (.C(w1193), .A(w1195), .B(w1380), .Z(w1194) );
	vdp_aoi21 g1473 (.A1(w1224), .B(SYSRES), .Z(w1204), .A2(w1223) );
	vdp_dff g1474 (.Q(w1267), .R(w1253), .C(w1250), .D(w1236) );
	vdp_dff g1475 (.Q(w1263), .R(w1253), .C(w1250), .D(w1262) );
	vdp_dff g1476 (.Q(w1233), .R(w1253), .C(w1250), .D(w1231) );
	vdp_dff g1477 (.Q(w1241), .R(w1253), .C(w1250), .D(w1240) );
	vdp_dff g1478 (.Q(w1242), .R(w1253), .C(w1250), .D(w1230) );
	vdp_dff g1479 (.Q(w1221), .R(w1253), .C(w1250), .D(w1258) );
	vdp_dff g1480 (.Q(w1218), .R(w1253), .C(w1250), .D(w1256) );
	vdp_dff g1481 (.Q(w1249), .R(1'b0), .C(w1250), .D(w1214) );
	vdp_ha g1482 (.SUM(w1256), .A(w1218), .B(w1213), .CO(w1219) );
	vdp_ha g1483 (.SUM(w1258), .A(w1221), .B(w1219), .CO(w1222) );
	vdp_ha g1484 (.SUM(w1230), .A(w1242), .B(w1222), .CO(w1229) );
	vdp_ha g1485 (.SUM(w1240), .A(w1241), .B(w1229), .CO(w1234) );
	vdp_ha g1486 (.SUM(w1231), .A(w1233), .B(w1234), .CO(w1232) );
	vdp_ha g1487 (.SUM(w1236), .A(w1267), .B(w1232), .CO(w1235) );
	vdp_ha g1488 (.SUM(w1262), .A(w1263), .B(w1235) );
	vdp_and3 g1489 (.A(w1263), .B(w1233), .Z(w1260), .C(w1267) );
	vdp_and4 g1490 (.C(w1221), .A(w1241), .B(w1260), .Z(w1266), .D(w1242) );
	vdp_nand g1491 (.A(w1249), .B(SEL0_M3), .Z(w1383) );
	vdp_dff g1492 (.Q(w1274), .R(1'b0), .C(w1250), .D(w1255) );
	vdp_dff g1493 (.Q(w1255), .R(w1257), .C(w1250), .D(w1279) );
	vdp_dff g1494 (.Q(w1279), .R(w1257), .C(w1277), .D(w1259) );
	vdp_dff g1495 (.Q(w1259), .R(w1257), .C(w1250), .D(w1283) );
	vdp_dff g1496 (.Q(w1283), .R(w1257), .C(w1250), .D(w1284) );
	vdp_dff g1497 (.Q(w1284), .R(w1257), .C(w1250), .D(1'b1) );
	vdp_dff g1498 (.Q(w1484), .R(w1293), .C(w1268), .D(w1260) );
	vdp_dff g1499 (.Q(w1268), .R(1'b0), .C(w1250), .D(w1266) );
	vdp_dff g1500 (.Q(w1286), .R(w1265), .C(w1287), .D(w1260) );
	vdp_dff g1501 (.Q(w1264), .R(w1278), .C(w1291), .D(1'b1) );
	vdp_or g1502 (.A(SYSRES), .B(w1264), .Z(w1265) );
	vdp_or g1503 (.A(w1257), .B(w1274), .Z(w1289) );
	vdp_not g1504 (.A(w1274), .nZ(w1252) );
	vdp_not g1505 (.A(w1484), .nZ(w1257) );
	vdp_nand3 g1506 (.A(SEL0_M3), .B(w1272), .Z(w1253), .C(w1252) );
	vdp_not g1507 (.nZ(w1277), .A(w1273) );
	vdp_not g1508 (.nZ(w1250), .A(w1251) );
	vdp_dff g1509 (.Q(w1276), .R(1'b0), .C(w1277), .D(w1298) );
	vdp_dff g1510 (.Q(w1301), .R(w1278), .C(w1277), .D(w1282) );
	vdp_dff g1511 (.Q(w1282), .R(w1278), .C(w1250), .D(w1303) );
	vdp_dff g1512 (.Q(w1303), .R(w1278), .C(w1277), .D(w1281) );
	vdp_dff g1513 (.Q(w1281), .R(w1278), .C(w1277), .D(w1292) );
	vdp_dff g1514 (.Q(w1292), .R(w1278), .C(w1250), .D(w47) );
	vdp_dff g1515 (.Q(w1308), .R(w1307), .C(w1277), .D(w1097) );
	vdp_dff g1516 (.Q(w1097), .R(w1307), .C(w1250), .D(w1288) );
	vdp_not g1517 (.A(w1295), .nZ(w100) );
	vdp_not g1518 (.A(w967), .nZ(w1271) );
	vdp_not g1519 (.A(w1282), .nZ(w1280) );
	vdp_not g1520 (.A(w1279), .nZ(w1492) );
	vdp_not g1521 (.A(w1288), .nZ(w1307) );
	vdp_not g1522 (.A(w1045), .nZ(w1291) );
	vdp_not g1523 (.A(w1197), .nZ(w1485) );
	vdp_and g1524 (.A(w1289), .B(w1045), .Z(w1288) );
	vdp_and g1525 (.A(w1290), .B(w1288), .Z(w1287) );
	vdp_and g1526 (.A(w1308), .B(w1287), .Z(w47) );
	vdp_and g1527 (.A(w1283), .B(w1492), .Z(w1299) );
	vdp_and g1528 (.A(w1284), .B(w1492), .Z(w1300) );
	vdp_and g1529 (.A(w1275), .B(w958), .Z(w1297) );
	vdp_and g1530 (.A(w1275), .B(w1001), .Z(w1270) );
	vdp_and g1531 (.A(w967), .B(w1276), .Z(w1275) );
	vdp_and g1532 (.A(w100), .B(w1097), .Z(w1033) );
	vdp_nand g1533 (.A(w1281), .B(w1280), .Z(w1272) );
	vdp_nor g1534 (.A(w1278), .B(w1292), .Z(w1302) );
	vdp_or3 g1535 (.C(w1286), .A(SYSRES), .B(w1274), .Z(w1293) );
	vdp_oai21 g1536 (.A1(w1001), .B(w1271), .Z(w1295), .A2(w958) );
	vdp_dff g1537 (.Q(w1315), .R(1'b0), .C(w1250), .D(w1198) );
	vdp_rs_ff g1538 (.nQ(w1042), .R(w1316), .S(w1313) );
	vdp_not g1539 (.A(w1321), .nZ(PSG_Z80_CLK) );
	vdp_not g1540 (.A(REG_BUS[7]), .nZ(w1312) );
	vdp_and3 g1541 (.C(w1312), .A(w803), .B(M5), .Z(w1313) );
	vdp_or g1542 (.A(w1198), .B(SYSRES), .Z(w1316) );
	vdp_and g1543 (.A(w1333), .B(w576), .Z(w1334) );
	vdp_not g1544 (.A(w1290), .nZ(w1336) );
	vdp_and4 g1545 (.C(CA[21]), .A(w1166), .B(CA[20]), .Z(w1290), .D(w1485) );
	vdp_dff g1546 (.Q(w1373), .R(1'b0), .C(w1321), .D(w1358) );
	vdp_dff g1547 (.Q(w1353), .R(1'b0), .C(w1321), .D(w1352) );
	vdp_dff g1548 (.Q(w1296), .R(1'b0), .C(w1339), .D(w1340) );
	vdp_dff g1549 (.Q(w1352), .R(1'b0), .C(w1339), .D(w1296) );
	vdp_dff g1550 (.Q(w1365), .R(w1366), .C(HCLK2), .D(w1368) );
	vdp_dff g1551 (.Q(DMA_BUSY), .R(w1366), .C(HCLK2), .D(w1365) );
	vdp_rs_ff g1552 (.Q(w1239), .R(w1366), .S(w1305) );
	vdp_rs_ff g1553 (.Q(w1486), .R(w1366), .S(w1237) );
	vdp_rs_ff g1554 (.Q(w1214), .R(w1306), .S(w1238) );
	vdp_sr_bit g1555 (.D(w576), .Q(w1333), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1556 (.D(w1493), .Q(w1364), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_dlatch_inv g1557 (.D(w1332), .nQ(w1311), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g1558 (.D(w1331), .nQ(w1332), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g1559 (.D(w1318), .C(HCLK1), .nQ(w1331), .nC(nHCLK1) );
	vdp_aon22 g1560 (.Z(w1360), .A2(w1310), .B1(w1331), .B2(w1369), .A1(w1311) );
	vdp_sr_bit g1561 (.D(w1370), .Q(w1375), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1562 (.D(w1335), .Q(w1370), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1563 (.D(VRAM_REFRESH), .C2(HCLK2), .C1(HCLK1), .Q(w1335), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_aon22 g1564 (.Z(w1348), .A2(w1302), .B1(w1376), .B2(w1377), .A1(w1346) );
	vdp_not g1565 (.A(w1483), .nZ(w1035) );
	vdp_not g1566 (.A(w1302), .nZ(w1377) );
	vdp_not g1567 (.A(w1364), .nZ(w1369) );
	vdp_not g1568 (.A(w1309), .nZ(w1347) );
	vdp_not g1569 (.A(w1286), .nZ(w1278) );
	vdp_or g1570 (.A(w1239), .B(w1486), .Z(w1368) );
	vdp_or g1571 (.A(SYSRES), .B(w578), .Z(w1366) );
	vdp_or g1572 (.A(w1305), .B(w1366), .Z(w1306) );
	vdp_or g1573 (.A(w1190), .B(w1188), .Z(w277) );
	vdp_or g1574 (.A(w1190), .B(w1189), .Z(w252) );
	vdp_and g1575 (.A(w1364), .B(w629), .Z(w1310) );
	vdp_or g1576 (.A(w1311), .B(w1370) );
	vdp_and g1577 (.A(w1272), .B(w1287), .Z(w1346) );
	vdp_and g1578 (.A(w1303), .B(w1287), .Z(w1376) );
	vdp_and g1579 (.A(w1287), .B(w1278), .Z(w102) );
	vdp_and g1580 (.A(w962), .B(w103), .Z(w1359) );
	vdp_or g1581 (.A(w1297), .B(w966), .Z(w1355) );
	vdp_aon22 g1582 (.Z(w1363), .A2(w1036), .B1(w1304), .B2(w1351), .A1(w1350) );
	vdp_and g1583 (.A(w1358), .B(w1373), .Z(w1096) );
	vdp_and g1584 (.A(w1371), .B(w1378), .Z(w1361) );
	vdp_and g1585 (.A(w1378), .B(w1374), .Z(w1358) );
	vdp_not g1586 (.A(w1374), .nZ(w1371) );
	vdp_not g1587 (.A(w1372), .nZ(w1378) );
	vdp_not g1588 (.A(w1332), .nZ(w1367) );
	vdp_not g1589 (.A(w1344), .nZ(w1362) );
	vdp_and g1590 (.A(w1356), .B(w1323), .Z(w1322) );
	vdp_and g1591 (.A(w1356), .B(w1325), .Z(w961) );
	vdp_and g1592 (.A(w1356), .B(w1327), .Z(w966) );
	vdp_and g1593 (.A(w1356), .B(w1324), .Z(w962) );
	vdp_and g1594 (.A(w1356), .B(w1326), .Z(w1340) );
	vdp_and g1595 (.A(w961), .B(w1340), .Z(w987) );
	vdp_and g1596 (.A(SEL0_M3), .B(w1337), .Z(w958) );
	vdp_and g1597 (.A(SEL0_M3), .B(w1328), .Z(w1001) );
	vdp_not g1598 (.A(SEL0_M3), .nZ(w1356) );
	vdp_nand g1599 (.A(w1352), .B(w1353), .Z(w1374) );
	vdp_nand g1600 (.A(FIFO_FULL), .B(w1320), .Z(w1319) );
	vdp_nand g1601 (.A(SEL0_M3), .B(w252), .Z(w1330) );
	vdp_nand g1602 (.A(w277), .B(SEL0_M3), .Z(w1329) );
	vdp_or3 g1603 (.C(w1190), .A(w1189), .B(w1188), .Z(w1028) );
	vdp_and3 g1604 (.C(w1311), .A(w576), .B(w1364), .Z(w581) );
	vdp_aoi21 g1605 (.A2(w1310), .B(w1367), .Z(w1309), .A1(w1331) );
	vdp_nor g1606 (.A(w1335), .B(w1375), .Z(w1320) );
	vdp_nand g1607 (.A(w100), .B(w1336), .Z(w1344) );
	vdp_nand3 g1608 (.C(w1319), .A(w3), .B(w1334), .Z(w1318) );
	vdp_2a3oi g1609 (.A1(w1367), .B(w654), .Z(w1317), .A2(w1331), .C(w1364) );
	vdp_nor4 g1610 (.C(VRAM_REFRESH), .A(w1370), .B(w1335), .Z(w1493), .D(w1375) );
	vdp_comb1 g1611 (.A1(CA[15]), .B(w1371), .Z(w1372), .A2(CA[14]), .C(w1322) );
	vdp_aon22 g1612 (.Z(w1294), .A2(w1036), .B1(w1304), .B2(w1345), .A1(w1482) );
	vdp_not g1613 (.A(w1036), .nZ(w1304) );
	vdp_or4 g1614 (.C(w1347), .A(w1378), .B(w1346), .Z(w1482), .D(w1299) );
	vdp_or4 g1615 (.C(w1311), .A(w1362), .B(w1359), .Z(w1351), .D(w1311) );
	vdp_or3 g1616 (.C(w1348), .A(w1358), .B(w1349), .Z(w1345) );
	vdp_comb1 g1617 (.A1(w1097), .B(w1282), .Z(w1483), .A2(w1302), .C(w1287) );
	vdp_and6 g1618 (.C(w1342), .A(w1249), .B(w1341), .Z(w1305), .D(w1315), .E(SEL0_M3), .F(w1291) );
	vdp_or5 g1619 (.C(w1360), .A(w1352), .B(w47), .Z(w1350), .D(w1300), .E(w1098) );
	vdp_or5 g1620 (.C(w1311), .A(w1361), .B(w101), .Z(w1354), .D(w1299), .E(w1359) );
	vdp_aoi22 g1621 (.Z(w1298), .A2(w47), .B1(w1301), .B2(w1287), .A1(w1302) );
	vdp_n_fet g1622 (.Z(w305), .A(w415) );
	vdp_n_fet g1623 (.Z(w262), .A(w415) );
	vdp_n_fet g1624 (.A(w415), .Z(w297) );
	vdp_n_fet g1625 (.A(w415), .Z(w254) );
	vdp_n_fet g1626 (.Z(w288), .A(w415) );
	vdp_n_fet g1627 (.Z(w245), .A(w415) );
	vdp_n_fet g1628 (.Z(w279), .A(w415) );
	vdp_n_fet g1629 (.Z(w237), .A(w415) );
	vdp_aon22 g1630 (.Z(w1349), .A2(w1310), .B1(w1310), .B2(w1367), .A1(w1311) );
	vdp_comp_we g1631 (.nZ(w1321), .Z(w1339), .A(w1357) );
	vdp_comp_we g1632 (.nZ(w1251), .Z(w1273), .A(w1384) );
	vdp_not g1633 (.nZ(w1574), .A(w1906) );
	vdp_not g1634 (.nZ(w1576), .A(w1577) );
	vdp_sr_bit g1635 (.Q(w5), .D(w1901), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1636 (.Q(w1582), .D(VPLA7), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1637 (.Q(w1558), .D(VPLA6), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1638 (.Q(w1605), .D(w1579), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1639 (.Q(w1559), .D(VPLA5), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1640 (.Q(w1563), .D(VPLA4), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1641 (.Q(w1745), .D(VPLA0), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1642 (.Q(w1590), .D(w1588), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1643 (.Q(w1587), .D(VPLA2), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1644 (.Q(w1564), .D(VPLA3), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1645 (.Q(w1597), .D(w1784), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1646 (.Q(w1595), .D(w1592), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1647 (.Q(w1592), .D(w1917), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1648 (.Q(w1596), .D(w1599), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1649 (.Q(w1569), .D(w1866), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_not g1650 (.nZ(w1588), .A(VPLA1) );
	vdp_not g1651 (.nZ(w58), .A(w1587) );
	vdp_not g1652 (.nZ(w1573), .A(w1587) );
	vdp_not g1653 (.nZ(w1566), .A(ODD_EVEN) );
	vdp_not g1654 (.nZ(w1575), .A(LSM0) );
	vdp_not g1655 (.nZ(w1917), .A(w1902) );
	vdp_not g1656 (.nZ(w1601), .A(w1602) );
	vdp_not g1657 (.nZ(w1589), .A(w1903) );
	vdp_not g1658 (.nZ(w1594), .A(w1595) );
	vdp_not g1659 (.nZ(w1571), .A(w53) );
	vdp_and g1660 (.Z(w1593), .A(w1780), .B(w1597) );
	vdp_nor g1661 (.Z(w1591), .A(SYSRES), .B(w1563) );
	vdp_oai21 g1662 (.Z(w1902), .B(w1591), .A2(w1601), .A1(w1592) );
	vdp_oai21 g1663 (.Z(w1602), .B(w1600), .A2(w1599), .A1(w1784) );
	vdp_aoi21 g1664 (.Z(w1903), .B(SYSRES), .A2(w1596), .A1(w1780) );
	vdp_and g1665 (.Z(w1570), .A(w1573), .B(w37) );
	vdp_and3 g1666 (.Z(w1780), .A(w1594), .B(w53), .C(w1592) );
	vdp_or g1667 (.Z(w1572), .A(SYSRES), .B(w1573) );
	vdp_and g1668 (.Z(w1866), .A(w1567), .B(w1577) );
	vdp_and g1669 (.Z(w1578), .A(w1570), .B(w1571) );
	vdp_and g1670 (.Z(w1567), .A(w1570), .B(w53) );
	vdp_and g1671 (.Z(w1562), .A(w1557), .B(w1564) );
	vdp_or g1672 (.Z(w1561), .A(SYSRES), .B(w1562) );
	vdp_2A3OI g1673 (.Z(w1906), .A1(w1576), .A2(w1567), .C(SYSRES), .B(w1575) );
	vdp_or g1674 (.Z(w1557), .A(w1565), .B(w1566) );
	vdp_or g1675 (.Z(w1560), .A(SYSRES), .B(w1603) );
	vdp_and g1676 (.Z(w1603), .A(w1557), .B(w1559) );
	vdp_and g1677 (.Z(w1583), .A(w1557), .B(w1582) );
	vdp_and g1678 (.Z(w1581), .A(w1557), .B(w1558) );
	vdp_or g1679 (.Z(w1855), .A(w1603), .B(SYSRES) );
	vdp_and g1680 (.Z(w1786), .A(w1579), .B(M5) );
	vdp_not g1681 (.nZ(w46), .A(w1585) );
	vdp_not g1682 (.nZ(w1585), .A(w1584) );
	vdp_not g1683 (.nZ(w1609), .A(w1584) );
	vdp_not g1684 (.nZ(w1901), .A(w1756) );
	vdp_and g1685 (.Z(w1675), .A(M5), .B(w1580) );
	vdp_or g1686 (.Z(w1586), .A(SYSRES), .B(w1583) );
	vdp_oai21 g1687 (.Z(w1584), .B(DISP), .A2(w29), .A1(w5) );
	vdp_rs_ff g1688 (.Q(w1580), .S(w1581), .R(w1586) );
	vdp_rs_ff g1689 (.Q(w1568), .R(w1560), .S(w1562) );
	vdp_rs_ff g1690 (.Q(w29), .S(w1590), .R(w1572) );
	vdp_rs_ff g1691 (.Q(w19), .R(w1563), .S(w1561) );
	vdp_tff g1692 (.C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .CI(w1578), .R(w1574), .A(w1569), .Q(ODD_EVEN) );
	vdp_cnt_bit_load g1693 (.D(w1776), .Q(w1641), .nL(w1884), .L(w1761), .CI(w1778), .nC1(nHCLK1), .CO(w1853), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g1694 (.Q(w1565), .D(HPLA13), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1695 (.Q(w1915), .D(HPLA0), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1696 (.Q(w30), .D(w1930), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1697 (.Q(w37), .D(HPLA14), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1698 (.Q(VRAM_REFRESH), .D(HPLA23), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1699 (.Q(w1643), .D(HPLA25), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1700 (.Q(w1637), .D(HPLA24), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1701 (.Q(w1613), .D(HPLA15), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1702 (.Q(w1638), .D(w1652), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1703 (.Q(w1599), .D(HPLA1), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1704 (.Q(w1783), .D(HPLA12), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1705 (.Q(w1667), .D(HPLA11), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1706 (.Q(w1784), .D(HPLA2), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1707 (.Q(w1652), .D(w1894), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1708 (.Q(w1793), .D(HPLA16), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1709 (.Q(w1647), .D(HPLA26), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1710 (.Q(w1666), .D(HPLA27), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1711 (.Q(w1928), .D(w1932), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1712 (.Q(w1699), .D(w1695), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1713 (.Q(w1649), .D(w1796), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1714 (.Q(w8), .D(HPLA28), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1715 (.Q(w1664), .D(HPLA17), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1716 (.Q(w1661), .D(w1842), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1717 (.Q(w1680), .D(HPLA10), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1718 (.Q(w1672), .D(HPLA3), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1719 (.Q(w1728), .D(w1676), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1720 (.Q(w27), .D(HPLA36), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1721 (.Q(w21), .D(HPLA29), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1722 (.Q(w1694), .D(HPLA18), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1723 (.Q(w1896), .D(w1734), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1724 (.Q(w1730), .D(HPLA9), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1725 (.Q(w1690), .D(HPLA4), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1726 (.Q(w1714), .D(HPLA35), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1727 (.Q(w28), .D(HPLA34), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1728 (.Q(w1716), .D(HPLA19), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1729 (.Q(w1717), .D(HPLA20), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1730 (.Q(w1743), .D(HPLA8), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1731 (.Q(w1691), .D(HPLA5), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1732 (.Q(w1604), .D(w1922), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1733 (.Q(w1678), .D(w1921), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1734 (.Q(w1729), .D(HPLA7), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1735 (.Q(w1692), .D(HPLA6), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1736 (.Q(w1733), .D(HPLA21), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1737 (.Q(w1711), .D(HPLA32), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1738 (.Q(w24), .D(HPLA31), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1739 (.Q(w1712), .D(w1604), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1740 (.Q(w1744), .D(w1700), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1741 (.Q(w1787), .D(HPLA22), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_not g1742 (.nZ(w1633), .A(M5) );
	vdp_not g1743 (.nZ(w6), .A(w1868) );
	vdp_not g1744 (.nZ(w38), .A(w1613) );
	vdp_not g1745 (.nZ(w1794), .A(w1608) );
	vdp_not g1746 (.nZ(w1617), .A(w53) );
	vdp_not g1747 (.nZ(w1619), .A(w1863) );
	vdp_not g1748 (.nZ(w1705), .A(w1) );
	vdp_not g1749 (.nZ(w1657), .A(w1625) );
	vdp_not g1750 (.nZ(w1639), .A(w1638) );
	vdp_not g1751 (.nZ(w1650), .A(w1613) );
	vdp_not g1752 (.nZ(w1651), .A(VSCR) );
	vdp_not g1753 (.nZ(w7), .A(w1645) );
	vdp_not g1754 (.nZ(w1635), .A(w39) );
	vdp_not g1755 (.nZ(w1927), .A(w53) );
	vdp_not g1756 (.nZ(w12), .A(w1890) );
	vdp_not g1757 (.nZ(w1891), .A(w1661) );
	vdp_not g1758 (.nZ(w1894), .A(w1671) );
	vdp_not g1759 (.nZ(w1704), .A(w1630) );
	vdp_not g1760 (.nZ(w1913), .A(w1629) );
	vdp_not g1761 (.nZ(w1655), .A(H40) );
	vdp_not g1762 (.nZ(w13), .A(w1702) );
	vdp_not g1763 (.nZ(w1883), .A(w1616) );
	vdp_not g1764 (.nZ(w1740), .A(w1674) );
	vdp_not g1765 (.nZ(w1718), .A(w1706) );
	vdp_not g1766 (.nZ(w1735), .A(w52) );
	vdp_not g1767 (.nZ(w1682), .A(w1838) );
	vdp_not g1768 (.nZ(w11), .A(w1869) );
	vdp_not g1769 (.nZ(w1746), .A(w1744) );
	vdp_not g1770 (.nZ(w1648), .A(w42) );
	vdp_not g1771 (.nZ(w1665), .A(w51) );
	vdp_not g1772 (.nZ(w1614), .A(w41) );
	vdp_not g1773 (.nZ(w1854), .A(w18) );
	vdp_not g1774 (.nZ(w1914), .A(w45) );
	vdp_not g1775 (.nZ(w1916), .A(M5) );
	vdp_not g1776 (.nZ(w1909), .A(w1683) );
	vdp_not g1777 (.nZ(w1760), .A(w1876) );
	vdp_not g1778 (.nZ(w1887), .A(w1861) );
	vdp_not g1779 (.nZ(w1762), .A(w1053) );
	vdp_not g1780 (.nZ(w1779), .A(w1777) );
	vdp_not g1781 (.nZ(w1773), .A(w1442) );
	vdp_not g1782 (.nZ(w1774), .A(PAL) );
	vdp_aon22 g1783 (.Z(w1937), .B1(w1764), .A1(w1763), .A2(DB[4]), .B2(w1762) );
	vdp_aon22 g1784 (.Z(w1875), .B1(w1764), .A1(w1763), .A2(DB[5]), .B2(w1750) );
	vdp_aon22 g1785 (.Z(w1877), .B1(w1764), .A1(w1763), .B2(w1887), .A2(DB[6]) );
	vdp_aon22 g1786 (.Z(w1872), .B2(1'b1), .A2(DB[7]), .B1(w1764), .A1(w1763) );
	vdp_aon22 g1787 (.Z(w1871), .B2(1'b1), .A2(DB[8]), .B1(w1764), .A1(w1763) );
	vdp_aon22 g1788 (.Z(w1753), .B2(1'b1), .B1(w1615), .A2(DB[8]), .A1(w1931) );
	vdp_aon22 g1789 (.Z(w1886), .B2(w1749), .A2(DB[3]), .B1(w1764), .A1(w1763) );
	vdp_aon22 g1790 (.Z(w1771), .A2(DB[2]), .B2(w1774), .B1(w1764), .A1(w1763) );
	vdp_aon22 g1791 (.Z(w1772), .A2(DB[1]), .B2(w1748), .B1(w1764), .A1(w1763) );
	vdp_aon22 g1792 (.Z(w1878), .A1(w1931), .B1(w1615), .B2(1'b1), .A2(DB[7]) );
	vdp_aon22 g1793 (.Z(w20), .A1(w1916), .B2(w1751), .B1(M5), .A2(w1728) );
	vdp_aon22 g1794 (.Z(w1721), .B1(w1615), .A1(w1931), .A2(DB[6]), .B2(1'b1) );
	vdp_aon22 g1795 (.Z(w1698), .B1(w1712), .B2(w1713), .A2(w1788), .A1(w1710) );
	vdp_not g1796 (.nZ(w1713), .A(w1710) );
	vdp_aon22 g1797 (.Z(w1879), .B1(w1615), .A1(w1931), .B2(1'b0), .A2(DB[5]) );
	vdp_not g1798 (.nZ(w1741), .A(w1738) );
	vdp_aon22 g1799 (.Z(w1923), .B1(w1615), .A1(w1931), .B2(w1883), .A2(DB[4]) );
	vdp_aon22 g1800 (.Z(w1880), .B2(w1882), .B1(w1615), .A2(DB[3]), .A1(w1931) );
	vdp_aon22 g1801 (.Z(w1696), .A2(w1633), .B2(M5), .A1(w1698), .B1(w1697) );
	vdp_aon22 g1802 (.Z(w1881), .A2(DB[2]), .B2(w1668), .A1(w1931), .B1(w1615) );
	vdp_aon22 g1803 (.Z(w1892), .B2(w1793), .B1(VSCR), .A2(w1651), .A1(w1650) );
	vdp_aon22 g1804 (.Z(w1642), .B1(w1867), .A1(HCLK2), .B2(w1635), .A2(w39) );
	vdp_aon22 g1805 (.Z(w1907), .A1(w1931), .B1(w1615), .B2(w1653), .A2(DB[1]) );
	vdp_aon22 g1806 (.Z(w1620), .A2(DB[0]), .B1(w1615), .B2(w1616), .A1(w1931) );
	vdp_not g1807 (.nZ(w4), .A(w1783) );
	vdp_not g1808 (.nZ(w3), .A(w1649) );
	vdp_rs_ff g1809 (.Q(w1693), .S(w1742), .R(w1857) );
	vdp_rs_ff g1810 (.Q(w1739), .R(w1730), .S(w1732) );
	vdp_rs_ff g1811 (.Q(w1676), .S(w1897), .R(w1692) );
	vdp_rs_ff g1812 (.Q(w1856), .R(w1926), .S(w1672) );
	vdp_rs_ff g1813 (.Q(w1677), .R(w1667), .S(w1920) );
	vdp_aon22 g1814 (.Z(w1776), .A2(DB[0]), .B2(w1747), .B1(w1764), .A1(w1763) );
	vdp_notif0 g1815 (.nZ(DB[1]), .A(VRAM_REFRESH), .nE(w1631) );
	vdp_notif0 g1816 (.nZ(DB[0]), .A(w30), .nE(w1631) );
	vdp_notif0 g1817 (.nZ(DB[7]), .A(w37), .nE(w1632) );
	vdp_notif0 g1818 (.A(w38), .nZ(DB[6]), .nE(w1632) );
	vdp_notif0 g1819 (.A(w6), .nZ(DB[2]), .nE(w1631) );
	vdp_notif0 g1820 (.A(w7), .nZ(DB[3]), .nE(w1631) );
	vdp_notif0 g1821 (.nZ(DB[5]), .A(w13), .nE(w1631) );
	vdp_notif0 g1822 (.A(w12), .nZ(DB[4]), .nE(w1631) );
	vdp_notif0 g1823 (.A(w15), .nZ(DB[5]), .nE(w1632) );
	vdp_notif0 g1824 (.nZ(DB[7]), .A(w8), .nE(w1631) );
	vdp_notif0 g1825 (.nZ(DB[6]), .A(w3), .nE(w1631) );
	vdp_notif0 g1826 (.nZ(DB[4]), .A(w16), .nE(w1632) );
	vdp_notif0 g1827 (.nZ(DB[9]), .A(w27), .nE(w1631) );
	vdp_notif0 g1828 (.nZ(DB[8]), .A(w21), .nE(w1631) );
	vdp_notif0 g1829 (.nZ(DB[3]), .A(w10), .nE(w1632) );
	vdp_notif0 g1830 (.nZ(DB[2]), .A(w26), .nE(w1632) );
	vdp_notif0 g1831 (.nZ(DB[10]), .A(w28), .nE(w1631) );
	vdp_notif0 g1832 (.nZ(DB[11]), .A(w11), .nE(w1631) );
	vdp_notif0 g1833 (.nZ(DB[12]), .A(w23), .nE(w1631) );
	vdp_notif0 g1834 (.nZ(DB[13]), .A(w24), .nE(w1631) );
	vdp_notif0 g1835 (.nZ(DB[1]), .A(w14), .nE(w1632) );
	vdp_notif0 g1836 (.nZ(DB[0]), .A(w9), .nE(w1632) );
	vdp_not g1837 (.nZ(VPOS[9]), .A(w1874) );
	vdp_not g1838 (.nZ(VPOS[8]), .A(w1873) );
	vdp_not g1839 (.nZ(VPOS[7]), .A(w1684) );
	vdp_not g1840 (.nZ(HPOS[7]), .A(w1909) );
	vdp_not g1841 (.nZ(HPOS[8]), .A(w1760) );
	vdp_not g1842 (.nZ(HPOS[6]), .A(w1682) );
	vdp_not g1843 (.nZ(VPOS[6]), .A(w1910) );
	vdp_not g1844 (.nZ(VPOS[5]), .A(w1911) );
	vdp_not g1845 (.nZ(HPOS[5]), .A(w1718) );
	vdp_not g1846 (.nZ(HPOS[4]), .A(w1740) );
	vdp_not g1847 (.nZ(VPOS[4]), .A(w1912) );
	vdp_not g1848 (.nZ(HPOS[3]), .A(w1913) );
	vdp_not g1849 (.nZ(VPOS[3]), .A(w1669) );
	vdp_not g1850 (.nZ(HPOS[2]), .A(w1704) );
	vdp_not g1851 (.nZ(VPOS[2]), .A(w1658) );
	vdp_not g1852 (.nZ(HPOS[1]), .A(w1657) );
	vdp_not g1853 (.nZ(VPOS[1]), .A(w1618) );
	vdp_not g1854 (.nZ(HPOS[0]), .A(w1619) );
	vdp_not g1855 (.nZ(VPOS[0]), .A(w1612) );
	vdp_aoi22 g1856 (.Z(w1867), .A1(w1605), .B1(w1634), .B2(M5), .A2(w1633) );
	vdp_aon22 g1857 (.Z(w1659), .A2(w1633), .B1(w1660), .B2(M5), .A1(w1700) );
	vdp_aoi22 g1858 (.Z(w1612), .B2(w1705), .B1(w1641), .A1(ODD_EVEN), .A2(w1) );
	vdp_aoi22 g1859 (.Z(w1618), .B2(w1705), .B1(w1781), .A1(w1641), .A2(w1) );
	vdp_aoi22 g1860 (.Z(w1658), .A2(w1), .A1(w1781), .B2(w1705), .B1(w1860) );
	vdp_aoi22 g1861 (.Z(w1669), .A1(w1860), .B2(w1705), .A2(w1), .B1(w1766) );
	vdp_aoi22 g1862 (.Z(w1912), .B1(w1859), .A1(w1766), .A2(w1), .B2(w1705) );
	vdp_aoi22 g1863 (.Z(w1911), .B1(w1720), .A1(w1859), .A2(w1), .B2(w1705) );
	vdp_aoi22 g1864 (.Z(w1910), .A2(w1), .B2(w1705), .B1(w1685), .A1(w1720) );
	vdp_aoi22 g1865 (.Z(w1684), .B2(w1705), .A1(w1685), .B1(w1755), .A2(w1) );
	vdp_aoi22 g1866 (.Z(w1873), .B2(w1705), .A2(w1), .A1(w1755), .B1(w1782) );
	vdp_aoi22 g1867 (.Z(w1874), .B1(1'b0), .A2(w1), .B2(w1705), .A1(w1782) );
	vdp_comp_dff g1868 (.Q(w1600), .D(w1636), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_comp_dff g1869 (.Q(w1736), .D(w1898), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_cnt_bit g1870 (.CI(w1900), .Q(w1788), .nEN(SYSRES), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g1871 (.nZ(w1870), .A(w55) );
	vdp_and g1872 (.Z(w1723), .A(w1738), .B(w1677) );
	vdp_and g1873 (.Z(w1724), .A(w1738), .B(w1677) );
	vdp_and g1874 (.Z(w1726), .A(w1925), .B(w1739) );
	vdp_and g1875 (.Z(w1727), .A(w1739), .B(w1741) );
	vdp_and g1876 (.Z(w1725), .A(w1786), .B(w1693) );
	vdp_and g1877 (.Z(w1925), .A(w1785), .B(w1675) );
	vdp_and g1878 (.Z(w1668), .A(w53), .B(w1655) );
	vdp_and g1879 (.Z(w15), .A(w1892), .B(w1646) );
	vdp_and g1880 (.Z(w1653), .A(w1617), .B(w1655) );
	vdp_and g1881 (.Z(w25), .A(w1585), .B(w1856) );
	vdp_and g1882 (.Z(w1654), .A(w52), .B(w1736) );
	vdp_and g1883 (.Z(w1679), .A(w1854), .B(w53) );
	vdp_and g1884 (.Z(w14), .A(w1646), .B(w1733) );
	vdp_and g1885 (.Z(w1865), .A(w1914), .B(w1679) );
	vdp_and g1886 (.Z(w9), .A(w1787), .B(w1646) );
	vdp_and g1887 (.Z(w1885), .A(w1745), .B(w4) );
	vdp_or g1888 (.Z(w1750), .A(w1858), .B(w1861) );
	vdp_or g1889 (.Z(w1749), .A(w1888), .B(w1861) );
	vdp_and g1890 (.Z(w1710), .A(M5), .B(w22) );
	vdp_and g1891 (.Z(w1900), .A(w1746), .B(w1700) );
	vdp_or g1892 (.Z(w1732), .A(SYSRES), .B(w1731) );
	vdp_or g1893 (.Z(w26), .A(w1717), .B(w1716) );
	vdp_or g1894 (.Z(w23), .A(w1711), .B(w1717) );
	vdp_or g1895 (.Z(w1922), .A(w1723), .B(w1727) );
	vdp_or g1896 (.Z(w1742), .A(w1729), .B(w1690) );
	vdp_or g1897 (.Z(w1857), .A(SYSRES), .B(w1731) );
	vdp_or g1898 (.Z(w1731), .A(w1680), .B(w1743) );
	vdp_or g1899 (.Z(w1897), .A(w1691), .B(SYSRES) );
	vdp_or g1900 (.Z(w1882), .A(w1616), .B(w1924) );
	vdp_or g1901 (.Z(w1926), .A(SYSRES), .B(w1690) );
	vdp_or g1902 (.Z(w1895), .A(w1654), .B(w1600) );
	vdp_or g1903 (.Z(w1842), .A(w1896), .B(w1734) );
	vdp_and g1904 (.Z(w10), .A(w1694), .B(w1646) );
	vdp_and g1905 (.Z(w1734), .A(w1606), .B(w1679) );
	vdp_or g1906 (.Z(w1920), .A(SYSRES), .B(w1680) );
	vdp_not g1907 (.nZ(w1632), .A(w54) );
	vdp_not g1908 (.nZ(w1631), .A(w48) );
	vdp_aon33 g1909 (.Z(w1778), .A3(w1777), .A2(w1870), .A1(w4), .B1(w55), .B3(1'b1), .B2(w1199) );
	vdp_aoi21 g1910 (.Z(w1868), .A1(w1637), .A2(w1646), .B(w1607) );
	vdp_aoi21 g1911 (.Z(w1645), .A1(w1643), .B(w1644), .A2(w1646) );
	vdp_aoi21 g1912 (.Z(w1608), .A1(w40), .A2(w50), .B(w1640) );
	vdp_aoi21 g1913 (.Z(w1671), .A1(w1652), .B(w1893), .A2(w1895) );
	vdp_aoi21 g1914 (.Z(w1890), .A1(w1646), .B(w1889), .A2(w1647) );
	vdp_aoi21 g1915 (.Z(w1702), .B(w1899), .A1(w1646), .A2(w1666) );
	vdp_aoi21 g1916 (.Z(w1869), .A1(w1646), .A2(w1714), .B(w1715) );
	vdp_xor g1917 (.Z(w1700), .B(w1605), .A(w1678) );
	vdp_xor g1918 (.Z(w1747), .A(ODD_EVEN), .B(w1774) );
	vdp_and3 g1919 (.Z(w1607), .A(w1665), .B(w42), .C(w1614) );
	vdp_and3 g1920 (.Z(w1930), .A(w1929), .B(w1792), .C(w1662) );
	vdp_and3 g1921 (.Z(w1644), .A(w1648), .B(w51), .C(w1614) );
	vdp_and3 g1922 (.Z(w1889), .A(w51), .B(w1614), .C(w42) );
	vdp_and3 g1923 (.Z(w1899), .A(w1648), .B(w1665), .C(w1717) );
	vdp_and3 g1924 (.Z(w1715), .A(w42), .B(w1665), .C(w41) );
	vdp_or3 g1925 (.Z(w1921), .A(w1725), .B(w1726), .C(w1724) );
	vdp_and3 g1926 (.Z(w1924), .A(w53), .B(w1655), .C(M5) );
	vdp_and3 g1927 (.Z(w1803), .A(w1652), .B(w53), .C(w1639) );
	vdp_and3 g1928 (.Z(w1616), .A(H40), .B(M5), .C(w1617) );
	vdp_nor4 g1929 (.Z(w1662), .A(HPLA33), .B(HPLA35), .C(HPLA29), .D(HPLA36) );
	vdp_nor4 g1930 (.Z(w1777), .A(w56), .B(w1780), .D(w1885), .C(SYSRES) );
	vdp_comp_we g1931 (.Z(w1761), .nZ(w1884), .A(w1779) );
	vdp_comp_we g1932 (.Z(w1763), .nZ(w1764), .A(w56) );
	vdp_comp_we g1933 (.Z(w1931), .nZ(w1615), .A(w57) );
	vdp_comp_we g1934 (.Z(w1622), .nZ(w1621), .A(w1606) );
	vdp_and3 g1935 (.Z(w17), .A(DISP), .B(w1856), .C(w29) );
	vdp_or4 g1936 (.Z(w1606), .A(w57), .B(SYSRES), .C(w1803), .D(w1915) );
	vdp_nor3 g1937 (.Z(w1792), .A(HPLA28), .B(HPLA30), .C(HPLA27) );
	vdp_nor3 g1938 (.Z(w1738), .A(w1675), .B(w1786), .C(w1785) );
	vdp_nand g1939 (.Z(w1695), .A(w1696), .B(w1735) );
	vdp_nand g1940 (.Z(w1932), .A(w1659), .B(w1927) );
	vdp_nand g1941 (.Z(w1796), .A(w1891), .B(HPLA30) );
	vdp_nor3 g1942 (.Z(w1646), .A(w42), .B(w51), .C(w41) );
	vdp_nor g1943 (.Z(w1861), .A(w1774), .B(M5) );
	vdp_nor g1944 (.Z(w1748), .A(ODD_EVEN), .B(w1774) );
	vdp_nor g1945 (.Z(w1858), .A(w1762), .B(PAL) );
	vdp_nor g1946 (.Z(w1888), .A(w1762), .B(w1774) );
	vdp_nor g1947 (.Z(w1893), .A(w1599), .B(SYSRES) );
	vdp_SDELAY8 g1948 (.Q(w1751), .D(w1728), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2), .nC3(nHCLK1), .C3(HCLK1), .nC4(nHCLK2), .C4(HCLK2), .nC5(nHCLK1), .C5(HCLK1), .nC6(nHCLK2), .C6(HCLK2), .nC7(nHCLK1), .C7(HCLK1), .nC8(nHCLK2), .C8(HCLK2), .nC9(nHCLK1), .C9(HCLK1), .nC10(nHCLK2), .C10(HCLK2), .nC11(nHCLK1), .C11(HCLK1), .nC12(nHCLK2), .C12(HCLK2), .nC13(nHCLK1), .C13(HCLK1), .nC14(nHCLK2), .C14(HCLK2), .nC15(nHCLK1), .C15(HCLK1), .nC16(nHCLK2), .C16(HCLK2) );
	vdp_SDELAY7 g1949 (.Q(w1697), .D(w1698), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .nC4(nHCLK2), .C5(HCLK1), .nC5(nHCLK1), .C6(HCLK2), .nC6(nHCLK2), .C7(HCLK1), .nC7(nHCLK1), .C8(HCLK2), .nC8(nHCLK2), .C9(HCLK1), .nC9(nHCLK1), .C10(HCLK2), .nC10(nHCLK2), .C11(HCLK1), .nC11(nHCLK1), .C12(HCLK2), .nC12(nHCLK2), .C13(HCLK1), .nC13(nHCLK1), .C14(HCLK2), .nC14(nHCLK2), .C3(HCLK1) );
	vdp_SDELAY8 g1950 (.Q(w1660), .D(w1700), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2), .C3(HCLK1), .nC4(nHCLK2), .C4(HCLK2), .nC5(nHCLK1), .C5(HCLK1), .nC6(nHCLK2), .C6(HCLK2), .nC7(nHCLK1), .C7(HCLK1), .nC8(nHCLK2), .C8(HCLK2), .nC9(nHCLK1), .C9(HCLK1), .nC10(nHCLK2), .C10(HCLK2), .C11(HCLK1), .nC12(nHCLK2), .C12(HCLK2), .nC13(nHCLK1), .C13(HCLK1), .nC14(nHCLK2), .C14(HCLK2), .nC15(nHCLK1), .C15(HCLK1), .nC16(nHCLK2), .C16(HCLK2), .nC3(nHCLK1), .nC11(nHCLK1) );
	vdp_SDELAY8 g1951 (.Q(w1634), .D(w1605), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2), .C3(HCLK1), .nC4(nHCLK2), .C4(HCLK2), .nC5(nHCLK1), .C5(HCLK1), .nC6(nHCLK2), .C6(HCLK2), .nC7(nHCLK1), .C7(HCLK1), .nC8(nHCLK2), .C8(HCLK2), .nC9(nHCLK1), .C9(HCLK1), .nC10(nHCLK2), .C10(HCLK2), .nC11(nHCLK1), .C11(HCLK1), .nC12(nHCLK2), .C12(HCLK2), .nC13(nHCLK1), .C13(HCLK1), .nC14(nHCLK2), .C14(HCLK2), .nC15(nHCLK1), .C15(HCLK1), .nC16(nHCLK2), .C16(HCLK2), .nC3(nHCLK1) );
	vdp_cnt_bit_load g1952 (.D(w1772), .Q(w1781), .nL(w1884), .L(w1761), .CI(w1853), .nC1(nHCLK1), .CO(w1934), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1953 (.D(w1771), .Q(w1860), .nL(w1884), .L(w1761), .CI(w1934), .nC1(nHCLK1), .CO(w1935), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1954 (.D(w1886), .Q(w1766), .nL(w1884), .L(w1761), .CI(w1935), .nC1(nHCLK1), .CO(w1936), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1955 (.D(w1937), .Q(w1859), .nL(w1884), .L(w1761), .CI(w1936), .nC1(nHCLK1), .CO(w1791), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1956 (.D(w1875), .Q(w1720), .nL(w1884), .L(w1761), .CI(w1791), .nC1(nHCLK1), .CO(w1790), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1957 (.D(w1877), .Q(w1685), .nL(w1884), .L(w1761), .CI(w1790), .nC1(nHCLK1), .CO(w1938), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1958 (.D(w1872), .Q(w1755), .nL(w1884), .L(w1761), .CI(w1938), .nC1(nHCLK1), .CO(w1789), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1959 (.D(w1871), .Q(w1782), .nL(w1884), .L(w1761), .CI(w1789), .nC1(nHCLK1), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1960 (.D(w1753), .Q(w1876), .nL(w1621), .L(w1622), .CI(w1754), .nC1(nHCLK1), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1961 (.D(w1878), .Q(w1683), .nL(w1621), .L(w1622), .CI(w1681), .nC1(nHCLK1), .CO(w1754), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1962 (.D(w1721), .Q(w1838), .nL(w1621), .L(w1622), .CI(w1719), .nC1(nHCLK1), .CO(w1681), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1963 (.D(w1879), .Q(w1706), .nL(w1621), .L(w1622), .CI(w1707), .nC1(nHCLK1), .CO(w1719), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1964 (.D(w1923), .Q(w1674), .nL(w1621), .L(w1622), .CI(w1673), .nC1(nHCLK1), .CO(w1707), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1965 (.D(w1880), .Q(w1629), .nL(w1621), .L(w1622), .CI(w1670), .nC1(nHCLK1), .CO(w1673), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1966 (.D(w1881), .Q(w1630), .nL(w1621), .L(w1622), .CI(w1656), .nC1(nHCLK1), .CO(w1670), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1967 (.D(w1907), .Q(w1625), .nL(w1621), .L(w1622), .CI(w1933), .nC1(nHCLK1), .CO(w1656), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1968 (.D(w1620), .Q(w1863), .nL(w1621), .L(w1622), .CI(w1794), .nC1(nHCLK1), .CO(w1933), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_or8 g1969 (.Z(VPLA7), .A(w1804), .B(w1805), .C(w1806), .D(w1807), .E(w1850), .F(w1851), .G(w1852), .H(w1808) );
	vdp_or8 g1970 (.Z(VPLA6), .A(w1809), .B(w1849), .C(w1848), .D(w1831), .E(w1847), .F(w1810), .G(w1811), .H(w1846) );
	vdp_or8 g1971 (.Z(VPLA5), .A(w1939), .B(w1918), .C(w1919), .D(w1905), .E(w1830), .F(w1829), .G(w1904), .H(w1828) );
	vdp_or5 g1972 (.Z(VPLA4), .A(w1824), .B(w1825), .C(w1826), .D(w1827), .E(w6542) );
	vdp_or7 g1973 (.Z(VPLA3), .A(w6619), .B(w6620), .C(w6618), .D(w1823), .E(w6539), .F(w6540), .G(w6541) );
	vdp_or7 g1974 (.Z(VPLA0), .A(w1812), .B(w1813), .C(w1814), .D(w1815), .E(w1816), .F(w1817), .G(w1818) );
	vdp_nor g1975 (.Z(w1640), .A(w1606), .B(w40) );
	vdp_and g1976 (.Z(w16), .A(w1646), .B(w1664) );
	vdp_not g1977 (.nZ(VPLA1), .A(w1819) );
	vdp_nor3 g1978 (.Z(VPLA2), .A(w1822), .B(w1821), .C(w1820) );
	vdp_rs_ff g1979 (.S(w1855), .R(w1581), .Q(w1579) );
	vdp_rs_ff g1980 (.S(w1593), .R(w1589), .Q(w1577) );
	vdp_and g1981 (.Z(w1785), .A(w1568), .B(M5) );
	vdp_nor4 g1982 (.Z(w1929), .A(HPLA23), .B(HPLA25), .C(HPLA24), .D(HPLA26) );
	vdp_nand3 g1983 (.A(w2060), .B(w2059), .C(w2057), .Z(w2053) );
	vdp_nand3 g1984 (.A(w2057), .B(w2059), .C(w2062), .Z(w2048) );
	vdp_nand3 g1985 (.A(w2057), .B(w2060), .C(w2061), .Z(w2049) );
	vdp_nand3 g1986 (.A(w2061), .B(w2057), .C(w2062), .Z(w2050) );
	vdp_nand3 g1987 (.A(w2061), .B(w2058), .C(w2062), .Z(w2045) );
	vdp_nand3 g1988 (.A(w2058), .B(w2060), .C(w2061), .Z(w2044) );
	vdp_nand3 g1989 (.A(w2059), .B(w2058), .C(w2062), .Z(w2052) );
	vdp_nand3 g1990 (.A(w2060), .B(w2059), .C(w2058), .Z(w2051) );
	vdp_nand3 g1991 (.A(w2033), .B(w2034), .C(w2029), .Z(w2043) );
	vdp_nand3 g1992 (.A(w2029), .B(w2034), .C(w2032), .Z(w2042) );
	vdp_nand3 g1993 (.A(w2031), .B(w2030), .C(w2032), .Z(w2036) );
	vdp_nand3 g1994 (.A(w2030), .B(w2033), .C(w2031), .Z(w2037) );
	vdp_nand3 g1995 (.A(w2034), .B(w2030), .C(w2032), .Z(w2038) );
	vdp_nand3 g1996 (.A(w2033), .B(w2034), .C(w2030), .Z(w2039) );
	vdp_nand3 g1997 (.A(w2031), .B(w2029), .C(w2032), .Z(w2040) );
	vdp_nand3 g1998 (.A(w2029), .B(w2033), .C(w2031), .Z(w2041) );
	vdp_nand3 g1999 (.A(w2021), .B(w2019), .C(w2017), .Z(w2014) );
	vdp_nand3 g2000 (.A(w2017), .B(w2019), .C(w2022), .Z(w2013) );
	vdp_nand3 g2001 (.A(w2020), .B(w2018), .C(w2022), .Z(w2007) );
	vdp_nand3 g2002 (.A(w2018), .B(w2021), .C(w2020), .Z(w2008) );
	vdp_nand3 g2003 (.A(w2019), .B(w2018), .C(w2022), .Z(w2009) );
	vdp_nand3 g2004 (.A(w2021), .B(w2019), .C(w2018), .Z(w2010) );
	vdp_nand3 g2005 (.A(w2020), .B(w2017), .C(w2022), .Z(w2011) );
	vdp_nand3 g2006 (.A(w2017), .B(w2021), .C(w2020), .Z(w2012) );
	vdp_nand3 g2007 (.A(w1960), .B(w1957), .C(w1961), .Z(w1954) );
	vdp_nand3 g2008 (.A(w1961), .B(w1957), .C(w1959), .Z(w1953) );
	vdp_nand3 g2009 (.A(w1958), .B(w1956), .C(w1959), .Z(w1947) );
	vdp_nand3 g2010 (.A(w1956), .B(w1960), .C(w1958), .Z(w1948) );
	vdp_nand3 g2011 (.A(w1957), .B(w1956), .C(w1959), .Z(w1949) );
	vdp_nand3 g2012 (.A(w1960), .B(w1957), .C(w1956), .Z(w1950) );
	vdp_nand3 g2013 (.A(w1958), .B(w1961), .C(w1959), .Z(w1951) );
	vdp_nand3 g2014 (.A(w1961), .B(w1960), .C(w1958), .Z(w1952) );
	vdp_not g2015 (.nZ(w1955), .A(w1942) );
	vdp_not g2016 (.nZ(w2015), .A(w1943) );
	vdp_not g2017 (.nZ(w2023), .A(w1940) );
	vdp_not g2018 (.nZ(w2054), .A(w1941) );
	vdp_nand g2019 (.Z(w1945), .B(w1946), .A(w1955) );
	vdp_nand g2020 (.Z(w1946), .B(w1955), .A(w1962) );
	vdp_nand g2021 (.Z(w2005), .B(w2006), .A(w2015) );
	vdp_nand g2022 (.Z(w2006), .B(w2015), .A(w1966) );
	vdp_comp_we g2023 (.A(w2016), .Z(w2018), .nZ(w2017) );
	vdp_comp_we g2024 (.A(w2076), .Z(w2020), .nZ(w2019) );
	vdp_comp_we g2025 (.A(w2075), .Z(w2022), .nZ(w2021) );
	vdp_comp_we g2026 (.A(w1963), .Z(w1956), .nZ(w1961) );
	vdp_comp_we g2027 (.A(w1964), .Z(w1958), .nZ(w1957) );
	vdp_comp_we g2028 (.A(w1965), .Z(w1959), .nZ(w1960) );
	vdp_nand g2029 (.Z(w2024), .B(w2023), .A(w2027) );
	vdp_comp_we g2030 (.A(w2026), .Z(w2030), .nZ(w2029) );
	vdp_comp_we g2031 (.A(w2028), .Z(w2031), .nZ(w2034) );
	vdp_comp_we g2032 (.A(w2035), .Z(w2032), .nZ(w2033) );
	vdp_nand g2033 (.Z(w2025), .B(w2024), .A(w2023) );
	vdp_nand g2034 (.Z(w2046), .B(w2054), .A(w2055) );
	vdp_comp_we g2035 (.A(w2056), .Z(w2058), .nZ(w2057) );
	vdp_comp_we g2036 (.A(w2063), .Z(w2061), .nZ(w2059) );
	vdp_comp_we g2037 (.A(w2064), .Z(w2062), .nZ(w2060) );
	vdp_nand g2038 (.Z(w2047), .B(w2046), .A(w2054) );
	vdp_comp_str g2039 (.A(w2087), .Z(w2088), .nZ(w2086) );
	vdp_comp_str g2040 (.A(w2104), .Z(w2077), .nZ(w2078) );
	vdp_comp_str g2041 (.A(w2113), .Z(w2068), .nZ(w2067) );
	vdp_comp_str g2042 (.A(w2114), .Z(w1969), .nZ(w1968) );
	vdp_comp_str g2043 (.A(w1977), .Z(w1978), .nZ(w1979) );
	vdp_comp_str g2044 (.A(w2151), .Z(w2337), .nZ(w2214) );
	vdp_comp_str g2045 (.A(w2362), .Z(w2330), .nZ(w2329) );
	vdp_comp_str g2046 (.A(w2333), .Z(w2343), .nZ(w2331) );
	vdp_comp_str g2047 (.A(w2122), .Z(w2334), .nZ(w2332) );
	vdp_comp_str g2048 (.A(w2242), .Z(w1985), .nZ(w1989) );
	vdp_comp_str g2049 (.A(w2363), .Z(w1986), .nZ(w1990) );
	vdp_comp_str g2050 (.A(w2120), .Z(w1988), .nZ(w1991) );
	vdp_slatch g2051 (.Q(w2347), .C(w1988), .D(w2115), .nC(w1991) );
	vdp_slatch g2052 (.Q(w2346), .C(w1986), .D(w2115), .nC(w1990) );
	vdp_slatch g2053 (.Q(w2309), .C(w1988), .D(w2249), .nC(w1991) );
	vdp_slatch g2054 (.Q(w2345), .C(w1985), .D(w2115), .nC(w1989) );
	vdp_slatch g2055 (.Q(w2350), .C(w1988), .D(w2250), .nC(w1991) );
	vdp_slatch g2056 (.Q(w2308), .C(w1985), .D(w2249), .nC(w1989) );
	vdp_slatch g2057 (.Q(w2310), .C(w1986), .D(w2249), .nC(w1990) );
	vdp_slatch g2058 (.Q(w2244), .C(w1988), .D(w2252), .nC(w1991) );
	vdp_slatch g2059 (.Q(w2348), .C(w1985), .D(w2250), .nC(w1989) );
	vdp_slatch g2060 (.Q(w2349), .C(w1986), .D(w2250), .nC(w1990) );
	vdp_slatch g2061 (.Q(w1998), .C(w1988), .D(w1987), .nC(w1991) );
	vdp_slatch g2062 (.Q(w2243), .C(w1985), .D(w2252), .nC(w1989) );
	vdp_slatch g2063 (.Q(w2245), .C(w1986), .D(w2252), .nC(w1990) );
	vdp_slatch g2064 (.Q(w1995), .C(w1985), .D(w1987), .nC(w1989) );
	vdp_slatch g2065 (.Q(w1997), .C(w1986), .D(w1987), .nC(w1990) );
	vdp_slatch g2066 (.Q(w1992), .C(w1988), .D(w1984), .nC(w1991) );
	vdp_slatch g2067 (.Q(w2004), .C(w1985), .D(w1984), .nC(w1989) );
	vdp_slatch g2068 (.Q(w1993), .C(w1986), .D(w1984), .nC(w1990) );
	vdp_slatch g2069 (.Q(w2323), .C(w2334), .D(w2115), .nC(w2332) );
	vdp_slatch g2070 (.Q(w2322), .C(w2343), .D(w2115), .nC(w2331) );
	vdp_slatch g2071 (.Q(w2328), .C(w2334), .D(w2249), .nC(w2332) );
	vdp_slatch g2072 (.Q(w2324), .C(w2330), .D(w2115), .nC(w2329) );
	vdp_slatch g2073 (.Q(w2316), .C(w2334), .D(w2250), .nC(w2332) );
	vdp_slatch g2074 (.Q(w2326), .C(w2330), .D(w2249), .nC(w2329) );
	vdp_slatch g2075 (.Q(w2327), .C(w2343), .D(w2249), .nC(w2331) );
	vdp_slatch g2076 (.Q(w2313), .C(w2334), .D(w2252), .nC(w2332) );
	vdp_slatch g2077 (.Q(w2314), .C(w2330), .D(w2250), .nC(w2329) );
	vdp_slatch g2078 (.Q(w2315), .C(w2343), .D(w2250), .nC(w2331) );
	vdp_slatch g2079 (.Q(w2311), .C(w2330), .D(w2252), .nC(w2329) );
	vdp_slatch g2080 (.Q(w2312), .C(w2343), .D(w2252), .nC(w2331) );
	vdp_slatch g2081 (.Q(w2198), .C(w2337), .D(w2250), .nC(w2214) );
	vdp_slatch g2082 (.Q(w2340), .C(w2337), .D(w2249), .nC(w2214) );
	vdp_slatch g2083 (.Q(w2341), .C(w2337), .D(w2115), .nC(w2214) );
	vdp_and g2084 (.Z(w2158), .A(w2341), .B(w2340) );
	vdp_and g2085 (.Z(w2325), .A(w2340), .B(w2338) );
	vdp_and g2086 (.Z(w2307), .A(w2341), .B(w2339) );
	vdp_and g2087 (.Z(w2253), .A(w2338), .B(w2339) );
	vdp_slatch g2088 (.Q(w2090), .C(w2088), .D(w2084), .nC(w2086) );
	vdp_or g2089 (.Z(w2064), .A(w2089), .B(w2090) );
	vdp_notif0 g2090 (.A(w2064), .nZ(DB[0]), .nE(w1970) );
	vdp_slatch g2091 (.Q(w2365), .C(w2088), .D(w2081), .nC(w2086) );
	vdp_or g2092 (.Z(w2063), .A(w2089), .B(w2365) );
	vdp_notif0 g2093 (.A(w2063), .nZ(DB[1]), .nE(w1970) );
	vdp_slatch g2094 (.Q(w2366), .C(w2088), .D(w2083), .nC(w2086) );
	vdp_or g2095 (.Z(w2056), .A(w2089), .B(w2366) );
	vdp_notif0 g2096 (.A(w2056), .nZ(DB[2]), .nE(w1970) );
	vdp_slatch g2097 (.Q(w2094), .C(w2088), .D(w2095), .nC(w2086) );
	vdp_or g2098 (.Z(w2055), .A(w2089), .B(w2094) );
	vdp_notif0 g2099 (.A(w2055), .nZ(DB[3]), .nE(w1970) );
	vdp_slatch g2100 (.Q(w2085), .C(w2077), .D(w2084), .nC(w2078) );
	vdp_or g2101 (.Z(w2035), .A(w2082), .B(w2085) );
	vdp_notif0 g2102 (.A(w2035), .nZ(DB[4]), .nE(w1970) );
	vdp_slatch g2103 (.Q(w2080), .C(w2077), .D(w2081), .nC(w2078) );
	vdp_or g2104 (.Z(w2028), .A(w2082), .B(w2080) );
	vdp_notif0 g2105 (.A(w2028), .nZ(DB[5]), .nE(w1970) );
	vdp_slatch g2106 (.Q(w2079), .C(w2077), .D(w2083), .nC(w2078) );
	vdp_or g2107 (.Z(w2026), .A(w2082), .B(w2079) );
	vdp_notif0 g2108 (.A(w2026), .nZ(DB[6]), .nE(w1970) );
	vdp_slatch g2109 (.Q(w2074), .C(w2077), .D(w2095), .nC(w2078) );
	vdp_or g2110 (.Z(w2027), .A(w2082), .B(w2074) );
	vdp_notif0 g2111 (.A(w2027), .nZ(DB[7]), .nE(w1970) );
	vdp_slatch g2112 (.Q(w2364), .C(w2068), .D(w2084), .nC(w2067) );
	vdp_or g2113 (.Z(w2075), .A(w2069), .B(w2364) );
	vdp_notif0 g2114 (.A(w2075), .nZ(DB[8]), .nE(w1970) );
	vdp_slatch g2115 (.Q(w2073), .C(w2068), .D(w2081), .nC(w2067) );
	vdp_or g2116 (.Z(w2076), .A(w2069), .B(w2073) );
	vdp_notif0 g2117 (.A(w2076), .nZ(DB[9]), .nE(w1970) );
	vdp_slatch g2118 (.Q(w2066), .C(w2068), .D(w2083), .nC(w2067) );
	vdp_or g2119 (.Z(w2016), .A(w2069), .B(w2066) );
	vdp_notif0 g2120 (.A(w2016), .nZ(DB[10]), .nE(w1970) );
	vdp_slatch g2121 (.Q(w2065), .C(w2068), .D(w2095), .nC(w2067) );
	vdp_or g2122 (.Z(w1966), .A(w2069), .B(w2065) );
	vdp_notif0 g2123 (.A(w1966), .nZ(DB[11]), .nE(w1970) );
	vdp_slatch g2124 (.Q(w1971), .C(w1969), .D(w2084), .nC(w1968) );
	vdp_or g2125 (.Z(w1965), .A(w1967), .B(w1971) );
	vdp_notif0 g2126 (.A(w1965), .nZ(DB[12]), .nE(w1970) );
	vdp_slatch g2127 (.Q(w1972), .C(w1969), .D(w2081), .nC(w1968) );
	vdp_or g2128 (.Z(w1964), .A(w1967), .B(w1972) );
	vdp_notif0 g2129 (.A(w1964), .nZ(DB[13]), .nE(w1970) );
	vdp_slatch g2130 (.Q(w1973), .C(w1969), .D(w2083), .nC(w1968) );
	vdp_or g2131 (.Z(w1963), .A(w1967), .B(w1973) );
	vdp_notif0 g2132 (.A(w1963), .nZ(DB[14]), .nE(w1970) );
	vdp_slatch g2133 (.Q(w1974), .C(w1969), .D(w2095), .nC(w1968) );
	vdp_or g2134 (.Z(w1962), .A(w1967), .B(w1974) );
	vdp_notif0 g2135 (.A(w1962), .nZ(DB[15]), .nE(w1970) );
	vdp_not g2136 (.A(PSG_TEST_OE), .nZ(w1970) );
	vdp_not g2137 (.nZ(w2143), .A(PSG_Z80_CLK) );
	vdp_clkgen g2138 (.PH(w2143), .CLK1(w2144), .nCLK1(w2145), .CLK2(w2146), .nCLK2(w2147) );
	vdp_comp_dff g2139 (.D(SYSRES), .nC1(w2145), .C1(w2144), .C2(w2146), .nC2(w2147), .Q(w2175) );
	vdp_sr_bit g2140 (.D(w2175), .nC1(w2145), .nC2(w2147), .C1(w2144), .C2(w2146), .Q(w2177) );
	vdp_sr_bit g2141 (.D(w2150), .nC1(w2145), .nC2(w2147), .C1(w2144), .C2(w2146), .Q(w2149) );
	vdp_not g2142 (.nZ(w2176), .A(w2177) );
	vdp_and g2143 (.Z(w2148), .A(w2175), .B(w2176) );
	vdp_nor g2144 (.Z(w2150), .A(w2149), .B(w2148) );
	vdp_cnt_bit g2145 (.CI(w2149), .R(w2148), .C1(w2144), .nC1(w2145), .nC2(w2147), .C2(w2146), .Q(w2174) );
	vdp_dlatch_inv g2146 (.nQ(w2173), .D(w2174), .nC(w2145), .C(w2144) );
	vdp_not g2147 (.nZ(w2172), .A(w2173) );
	vdp_nand g2148 (.Z(w2171), .A(w2149), .B(w2173) );
	vdp_not g2149 (.nZ(w2170), .A(w2171) );
	vdp_not g2150 (.nZ(w2169), .A(w2168) );
	vdp_not g2151 (.nZ(PSG_CLK1), .A(w2171) );
	vdp_not g2152 (.nZ(PSG_nCLK1), .A(w2170) );
	vdp_not g2153 (.nZ(PSG_nCLK2), .A(w2169) );
	vdp_not g2154 (.nZ(PSG_CLK2), .A(w2168) );
	vdp_nand g2155 (.Z(w2168), .A(w2149), .B(w2172) );
	vdp_sr_bit g2156 (.D(w2278), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2134) );
	vdp_sr_bit g2157 (.D(w2279), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2278) );
	vdp_sr_bit g2158 (.D(w2277), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2279) );
	vdp_sr_bit g2159 (.D(w2138), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2277) );
	vdp_sr_bit g2160 (.D(w2276), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2137) );
	vdp_sr_bit g2161 (.D(w2275), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2276) );
	vdp_sr_bit g2162 (.D(w2274), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2275) );
	vdp_sr_bit g2163 (.D(w2142), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2274) );
	vdp_sr_bit g2164 (.D(w2273), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2141) );
	vdp_sr_bit g2165 (.D(w2272), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2273) );
	vdp_sr_bit g2166 (.D(w2271), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2272) );
	vdp_sr_bit g2167 (.D(w2204), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2271) );
	vdp_sr_bit g2168 (.D(w2269), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2203) );
	vdp_sr_bit g2169 (.D(w2270), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2269) );
	vdp_sr_bit g2170 (.D(w2268), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2270) );
	vdp_sr_bit g2171 (.D(w2202), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2268) );
	vdp_sr_bit g2172 (.D(w2267), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2201) );
	vdp_sr_bit g2173 (.D(w2266), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2267) );
	vdp_sr_bit g2174 (.D(w2265), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2266) );
	vdp_sr_bit g2175 (.D(w2190), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2265) );
	vdp_sr_bit g2176 (.D(w2264), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2189) );
	vdp_sr_bit g2177 (.D(w2263), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2264) );
	vdp_sr_bit g2178 (.D(w2260), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2263) );
	vdp_sr_bit g2179 (.D(w2187), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2260) );
	vdp_sr_bit g2180 (.D(w2261), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2188) );
	vdp_sr_bit g2181 (.D(w2262), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2261) );
	vdp_sr_bit g2182 (.D(w2288), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2262) );
	vdp_sr_bit g2183 (.D(w2256), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2288) );
	vdp_sr_bit g2184 (.D(w2287), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2257) );
	vdp_sr_bit g2185 (.D(w2289), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2287) );
	vdp_sr_bit g2186 (.D(w2290), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2289) );
	vdp_sr_bit g2187 (.D(w2225), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2290) );
	vdp_sr_bit g2188 (.D(w2215), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2224) );
	vdp_sr_bit g2189 (.D(w2216), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2215) );
	vdp_sr_bit g2190 (.D(w2217), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2216) );
	vdp_sr_bit g2191 (.D(w2226), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2217) );
	vdp_sr_bit g2192 (.D(w2132), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2222) );
	vdp_sr_bit g2193 (.D(w2131), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2132) );
	vdp_sr_bit g2194 (.D(w2130), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2131) );
	vdp_sr_bit g2195 (.D(w2128), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2130) );
	vdp_aon2222 g2196 (.Z(w2000), .D2(1'b0), .C2(w2004), .C1(w1996), .D1(w2003), .B1(w1993), .A2(w1992), .A1(w1994), .B2(w2002) );
	vdp_cgi2a g2197 (.Z(w2342), .A(w2000), .C(w2354), .B(w2134) );
	vdp_aon2222 g2198 (.Z(w2001), .D2(1'b0), .C2(w1995), .C1(w1996), .D1(w2003), .B1(w1997), .A2(w1998), .A1(w1994), .B2(w2002) );
	vdp_cgi2a g2199 (.Z(w2354), .A(w2001), .C(w2353), .B(w2137) );
	vdp_aon2222 g2200 (.Z(w2248), .D2(1'b0), .C2(w2243), .C1(w1996), .D1(w2003), .B1(w2245), .A2(w2244), .A1(w1994), .B2(w2002) );
	vdp_cgi2a g2201 (.Z(w2353), .A(w2248), .C(w2352), .B(w2141) );
	vdp_aon2222 g2202 (.Z(w2247), .D2(w2325), .C2(w2348), .C1(w1996), .D1(w2003), .B1(w2349), .A2(w2350), .A1(w1994), .B2(w2002) );
	vdp_cgi2a g2203 (.Z(w2352), .A(w2247), .C(w2254), .B(w2203) );
	vdp_aon2222 g2204 (.Z(w2246), .D2(w2307), .C2(w2308), .C1(w1996), .D1(w2003), .B1(w2310), .A2(w2309), .A1(w1994), .B2(w2002) );
	vdp_cgi2a g2205 (.Z(w2254), .A(w2246), .C(w2255), .B(w2201) );
	vdp_aon2222 g2206 (.Z(w2318), .D2(w2253), .C2(w2345), .C1(w1996), .D1(w2003), .B1(w2346), .A2(w2347), .A1(w1994), .B2(w2002) );
	vdp_cgi2a g2207 (.Z(w2255), .A(w2318), .C(w2351), .B(w2189) );
	vdp_aon2222 g2208 (.Z(w2317), .D2(1'b0), .C2(w2311), .C1(w1996), .D1(w2003), .B1(w2312), .A2(w2313), .A1(w1994), .B2(w2002) );
	vdp_cgi2a g2209 (.Z(w2351), .A(w2317), .C(w2344), .B(w2188) );
	vdp_aon2222 g2210 (.Z(w2319), .D2(1'b0), .C2(w2314), .C1(w1996), .D1(w2003), .B1(w2315), .A2(w2316), .A1(w1994), .B2(w2002) );
	vdp_cgi2a g2211 (.Z(w2344), .A(w2319), .C(w2218), .B(w2257) );
	vdp_aon2222 g2212 (.Z(w2320), .D2(1'b0), .C2(w2326), .C1(w1996), .D1(w2003), .B1(w2327), .A2(w2328), .A1(w1994), .B2(w2002) );
	vdp_cgi2a g2213 (.Z(w2218), .A(w2320), .C(w2219), .B(w2224) );
	vdp_aon2222 g2214 (.Z(w2221), .D2(1'b0), .C2(w2324), .C1(w1996), .D1(w2003), .B1(w2322), .A2(w2323), .A1(w1994), .B2(w2002) );
	vdp_cgi2a g2215 (.Z(w2219), .A(w2221), .C(1'b1), .B(w2222) );
	vdp_not g2216 (.nZ(w2003), .A(w2321) );
	vdp_sr_bit g2217 (.D(w2302), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .Q(w2223) );
	vdp_nand g2218 (.Z(w2321), .A(w2297), .B(w2223) );
	vdp_not g2219 (.nZ(w1996), .A(w2303) );
	vdp_sr_bit g2220 (.D(w2298), .Q(w2302), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_nand g2221 (.Z(w2303), .A(w2297), .B(w2302) );
	vdp_not g2222 (.nZ(w2002), .A(w2301) );
	vdp_sr_bit g2223 (.D(w2234), .Q(w2298), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_nand g2224 (.Z(w2301), .A(w2297), .B(w2298) );
	vdp_not g2225 (.nZ(w1994), .A(w2299) );
	vdp_sr_bit g2226 (.D(w2300), .Q(w2234), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_nand g2227 (.Z(w2299), .A(w2297), .B(w2234) );
	vdp_sr_bit g2228 (.D(w2124), .Q(w2205), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_sr_bit g2229 (.D(w2306), .Q(w2304), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_sr_bit g2230 (.D(w2305), .Q(w2306), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_sr_bit g2231 (.D(w2233), .Q(w2305), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_sr_bit g2232 (.D(w2342), .Q(w2233), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_not g2233 (.nZ(w2297), .A(w2205) );
	vdp_nor4 g2234 (.Z(w2300), .A(w2302), .B(w2298), .D(w2234), .C(w2124) );
	vdp_nor4 g2235 (.Z(w2195), .A(w2237), .B(w2238), .D(w2235), .C(w2236) );
	vdp_nor4 g2236 (.Z(w2197), .A(w2230), .B(w2231), .D(w2210), .C(w2211) );
	vdp_nor3 g2237 (.Z(w2196), .A(w2206), .B(w2207), .C(w2208) );
	vdp_not g2238 (.nZ(w1982), .A(w2205) );
	vdp_nand4 g2239 (.Z(w2194), .A(w2195), .B(w2197), .D(w2165), .C(w2196) );
	vdp_nand g2240 (.Z(w2199), .A(w2133), .B(w2198) );
	vdp_nand g2241 (.Z(w2200), .A(w2194), .B(w2199) );
	vdp_lfsr_bit g2242 (.Q(w2230), .A(w2200), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2228), .B(w2229) );
	vdp_lfsr_bit g2243 (.Q(w2231), .A(w2230), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2228), .B(w2229) );
	vdp_lfsr_bit g2244 (.Q(w2211), .A(w2231), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2228), .B(w2229) );
	vdp_lfsr_bit g2245 (.Q(w2210), .A(w2211), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2228), .B(w2229) );
	vdp_lfsr_bit g2246 (.Q(w2206), .A(w2210), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2228), .B(w2229) );
	vdp_lfsr_bit g2247 (.Q(w2207), .A(w2206), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2228), .B(w2229) );
	vdp_lfsr_bit g2248 (.Q(w2208), .A(w2207), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2228), .B(w2229) );
	vdp_lfsr_bit g2249 (.Q(w2235), .A(w2208), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2228), .B(w2229) );
	vdp_lfsr_bit g2250 (.Q(w2236), .A(w2235), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2228), .B(w2229) );
	vdp_lfsr_bit g2251 (.Q(w2237), .A(w2236), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2228), .B(w2229) );
	vdp_lfsr_bit g2252 (.Q(w2238), .A(w2237), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2228), .B(w2229) );
	vdp_lfsr_bit g2253 (.Q(w2239), .A(w2238), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2228), .B(w2229) );
	vdp_lfsr_bit g2254 (.Q(w2240), .A(w2239), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2228), .B(w2229) );
	vdp_lfsr_bit g2255 (.Q(w2227), .A(w2240), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2228), .B(w2229) );
	vdp_lfsr_bit g2256 (.Q(w2127), .A(w2227), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2228), .B(w2229) );
	vdp_lfsr_bit g2257 (.Q(w2241), .A(w2127), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2228), .B(w2229) );
	vdp_xor g2258 (.Z(w2133), .A(w2240), .B(w2241) );
	vdp_and g2259 (.Z(w2286), .A(w2129), .B(w2222) );
	vdp_ha g2260 (.SUM(w2128), .CO(w2184), .B(w2286), .A(1'b1) );
	vdp_and g2261 (.Z(w2259), .A(w2129), .B(w2224) );
	vdp_ha g2262 (.SUM(w2226), .CO(w2183), .B(w2259), .A(w2184) );
	vdp_and g2263 (.Z(w2258), .A(w2129), .B(w2257) );
	vdp_ha g2264 (.SUM(w2225), .CO(w2182), .B(w2258), .A(w2183) );
	vdp_and g2265 (.Z(w2186), .A(w2129), .B(w2188) );
	vdp_ha g2266 (.SUM(w2256), .CO(w2181), .B(w2186), .A(w2182) );
	vdp_and g2267 (.Z(w2285), .A(w2129), .B(w2189) );
	vdp_ha g2268 (.SUM(w2187), .CO(w2180), .B(w2285), .A(w2181) );
	vdp_and g2269 (.Z(w2284), .A(w2129), .B(w2201) );
	vdp_ha g2270 (.SUM(w2190), .CO(w2179), .B(w2284), .A(w2180) );
	vdp_and g2271 (.Z(w2283), .A(w2129), .B(w2203) );
	vdp_ha g2272 (.SUM(w2202), .CO(w2178), .B(w2283), .A(w2179) );
	vdp_and g2273 (.Z(w2282), .A(w2129), .B(w2141) );
	vdp_ha g2274 (.SUM(w2204), .CO(w2140), .B(w2282), .A(w2178) );
	vdp_and g2275 (.Z(w2281), .A(w2129), .B(w2137) );
	vdp_ha g2276 (.SUM(w2142), .CO(w2139), .B(w2281), .A(w2140) );
	vdp_and g2277 (.Z(w2280), .A(w2129), .B(w2134) );
	vdp_ha g2278 (.SUM(w2138), .B(w2280), .A(w2139) );
	vdp_and g2279 (.Z(w2209), .A(w2234), .B(w2304) );
	vdp_cnt_bit g2280 (.CI(w2209), .R(w2205), .C1(PSG_CLK1), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C2(PSG_CLK2), .Q(w2335) );
	vdp_and g2281 (.Z(w2213), .A(w2234), .B(w2306) );
	vdp_cnt_bit g2282 (.CI(w2213), .R(w2205), .C1(PSG_CLK1), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C2(PSG_CLK2), .Q(w2336) );
	vdp_and g2283 (.Z(w2212), .A(w2234), .B(w2305) );
	vdp_cnt_bit g2284 (.CI(w2212), .R(w2205), .C1(PSG_CLK1), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C2(PSG_CLK2), .Q(w2159) );
	vdp_and g2285 (.Z(w2232), .A(w2234), .B(w2233) );
	vdp_cnt_bit g2286 (.CI(w2232), .R(w2205), .C1(PSG_CLK1), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C2(PSG_CLK2), .Q(w2152) );
	vdp_nor g2287 (.Z(w2129), .A(w2342), .B(w2205) );
	vdp_slatch g2288 (.Q(w1983), .C(w1980), .D(DB[7]), .nC(w1981) );
	vdp_comp_str g2289 (.A(w1030), .Z(w1980), .nZ(w1981) );
	vdp_and g2290 (.Z(w1975), .A(w1982), .B(w1983) );
	vdp_and g2291 (.Z(w1977), .A(w1976), .B(w1975) );
	vdp_and g2292 (.Z(w2361), .A(w1982), .B(w2360) );
	vdp_slatch g2293 (.Q(w2360), .C(w1980), .D(DB[6]), .nC(w1981) );
	vdp_slatch g2294 (.Q(w2103), .C(w1978), .D(w2361), .nC(w1979) );
	vdp_and g2295 (.Z(w1984), .A(w1982), .B(w2071) );
	vdp_slatch g2296 (.Q(w2071), .C(w1980), .D(DB[5]), .nC(w1981) );
	vdp_slatch g2297 (.Q(w2072), .C(w1978), .D(w1984), .nC(w1979) );
	vdp_and g2298 (.Z(w1987), .A(w1982), .B(w2070) );
	vdp_slatch g2299 (.Q(w2070), .C(w1980), .D(DB[4]), .nC(w1981) );
	vdp_slatch g2300 (.Q(w2102), .C(w1978), .D(w1987), .nC(w1979) );
	vdp_and g2301 (.Z(w2252), .A(w1982), .B(w2109) );
	vdp_slatch g2302 (.Q(w2109), .C(w1980), .D(DB[3]), .nC(w1981) );
	vdp_or g2303 (.Z(w2095), .A(w2110), .B(w2252) );
	vdp_and g2304 (.Z(w2250), .A(w1982), .B(w2359) );
	vdp_or g2305 (.Z(w2083), .A(w2110), .B(w2250) );
	vdp_slatch g2306 (.Q(w2359), .C(w1980), .D(DB[2]), .nC(w1981) );
	vdp_not g2307 (.nZ(w2110), .A(w1982) );
	vdp_and g2308 (.Z(w2249), .A(w1982), .B(w2251) );
	vdp_or g2309 (.Z(w2081), .A(w2110), .B(w2249) );
	vdp_slatch g2310 (.Q(w2251), .C(w1980), .D(DB[1]), .nC(w1981) );
	vdp_and g2311 (.Z(w2115), .A(w1982), .B(w2116) );
	vdp_or g2312 (.Z(w2084), .A(w2110), .B(w2115) );
	vdp_slatch g2313 (.Q(w2116), .C(w1980), .D(DB[0]), .nC(w1981) );
	vdp_not g2314 (.nZ(w2114), .A(w2112) );
	vdp_aoi21 g2315 (.Z(w2112), .B(w2124), .A1(w2117), .A2(w2111) );
	vdp_and3 g2316 (.Z(w2111), .A(w2092), .B(w2091), .C(w2102) );
	vdp_not g2317 (.nZ(w2113), .A(w2357) );
	vdp_aoi21 g2318 (.Z(w2357), .B(w2124), .A1(w2117), .A2(w2358) );
	vdp_and3 g2319 (.Z(w2358), .A(w2092), .B(w2072), .C(w2102) );
	vdp_not g2320 (.nZ(w2367), .A(w2356) );
	vdp_aoi21 g2321 (.Z(w2356), .B(w2124), .A1(w2117), .A2(w2355) );
	vdp_and3 g2322 (.Z(w2355), .A(w2103), .B(w2091), .C(w2093) );
	vdp_not g2323 (.nZ(w2121), .A(w1975) );
	vdp_or g2324 (.Z(w2123), .A(w1975), .B(w2124) );
	vdp_and g2325 (.Z(w2362), .A(w2123), .B(w2367) );
	vdp_and g2326 (.Z(w2242), .A(w2121), .B(w2367) );
	vdp_and g2327 (.Z(w2333), .A(w2123), .B(w2108) );
	vdp_and g2328 (.Z(w2363), .A(w2121), .B(w2108) );
	vdp_not g2329 (.nZ(w2108), .A(w2107) );
	vdp_aoi21 g2330 (.Z(w2107), .B(w2124), .A1(w2117), .A2(w2106) );
	vdp_and3 g2331 (.Z(w2106), .A(w2092), .B(w2072), .C(w2093) );
	vdp_not g2332 (.nZ(w2104), .A(w2105) );
	vdp_aoi21 g2333 (.Z(w2105), .B(w2124), .A1(w2117), .A2(w2119) );
	vdp_and3 g2334 (.Z(w2119), .A(w2103), .B(w2091), .C(w2102) );
	vdp_and g2335 (.Z(w2122), .A(w2123), .B(w2118) );
	vdp_and g2336 (.Z(w2120), .A(w2121), .B(w2118) );
	vdp_not g2337 (.nZ(w2118), .A(w2101) );
	vdp_aoi21 g2338 (.Z(w2101), .B(w2124), .A1(w2117), .A2(w2100) );
	vdp_and3 g2339 (.Z(w2100), .A(w2092), .B(w2091), .C(w2093) );
	vdp_and3 g2340 (.Z(w2099), .A(w2103), .B(w2072), .C(w2102) );
	vdp_not g2341 (.nZ(w2087), .A(w2098) );
	vdp_aoi21 g2342 (.Z(w2098), .B(w2124), .A1(w2117), .A2(w2099) );
	vdp_and3 g2343 (.Z(w2096), .A(w2103), .B(w2072), .C(w2093) );
	vdp_not g2344 (.nZ(w2151), .A(w2097) );
	vdp_aoi21 g2345 (.Z(w2097), .B(w2124), .A1(w2117), .A2(w2096) );
	vdp_not g2346 (.nZ(w2338), .A(w2341) );
	vdp_not g2347 (.nZ(w2339), .A(w2340) );
	vdp_not g2348 (.nZ(w2093), .A(w2102) );
	vdp_not g2349 (.nZ(w2091), .A(w2072) );
	vdp_not g2350 (.nZ(w2092), .A(w2103) );
	vdp_nor g2351 (.Z(w1967), .A(w2335), .B(w1123) );
	vdp_nor g2352 (.Z(w2069), .A(w2336), .B(w1123) );
	vdp_nor g2353 (.Z(w2082), .A(w2159), .B(w1123) );
	vdp_nor g2354 (.Z(w2089), .A(w2127), .B(w1123) );
	vdp_aon22 g2355 (.Z(w2154), .A2(w2159), .A1(w2158), .B2(w2153), .B1(w2152) );
	vdp_sr_bit g2356 (.D(w2154), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2155) );
	vdp_not g2357 (.nZ(w2153), .A(w2158) );
	vdp_not g2358 (.nZ(w2156), .A(w2155) );
	vdp_not g2359 (.nZ(w2292), .A(w1124) );
	vdp_not g2360 (.nZ(w2291), .A(w1125) );
	vdp_not g2361 (.nZ(w2192), .A(w2191) );
	vdp_sr_bit g2362 (.D(w1976), .nC1(w2145), .nC2(w2147), .C1(w2144), .C2(w2146), .Q(w2117) );
	vdp_nand g2363 (.Z(w2293), .A(w1124), .B(w2291) );
	vdp_nand g2364 (.Z(w2157), .A(w1125), .B(w6537) );
	vdp_nand g2365 (.Z(w2294), .A(w2291), .B(w2292) );
	vdp_nand g2366 (.Z(w2295), .A(w1125), .B(w2292) );
	vdp_and g2367 (.Z(w2161), .A(w2154), .B(w2156) );
	vdp_and g2368 (.Z(w1941), .A(w1123), .B(w2157) );
	vdp_and g2369 (.Z(w1943), .A(w1123), .B(w2293) );
	vdp_and g2370 (.Z(w1942), .A(w1123), .B(w2294) );
	vdp_and g2371 (.Z(w1940), .A(w1123), .B(w2295) );
	vdp_nor4 g2372 (.Z(w2165), .A(w2227), .B(w2240), .D(w2239), .C(w2127) );
	vdp_not g2373 (.nZ(w2162), .A(w2161) );
	vdp_not g2374 (.nZ(w2229), .A(w2163) );
	vdp_not g2375 (.nZ(w2228), .A(w2296) );
	vdp_not g2376 (.nZ(w2124), .A(w2192) );
	vdp_nand g2377 (.Z(w2163), .A(w2160), .B(w2162) );
	vdp_nand g2378 (.Z(w2296), .A(w2160), .B(w2161) );
	vdp_nor g2379 (.Z(w2160), .A(w2124), .B(w2164) );
	vdp_rs_ff g2380 (.S(w2151), .R(w2164), .Q(w2193) );
	vdp_rs_ff g2381 (.S(w1976), .R(w1030), .Q(w2166) );
	vdp_nor g2382 (.Z(w2167), .A(w1030), .B(w2166) );
	vdp_comp_dff g2383 (.D(w2167), .nC1(w2145), .C1(w2144), .C2(w2146), .nC2(w2147), .Q(w1976) );
	vdp_comp_dff g2384 (.D(SYSRES), .nC1(PSG_nCLK1), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC2(PSG_nCLK2), .Q(w2191) );
	vdp_comp_dff g2385 (.D(w2193), .nC1(PSG_nCLK1), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC2(PSG_nCLK2), .Q(w2164) );
	vdp_sr_bit g2386 (.Q(w2535), .D(w2529), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2387 (.nZ(AD_RD_DIR), .A(w2528) );
	vdp_sr_bit g2388 (.Q(w2536), .D(w2399), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2389 (.Q(w2464), .D(w2412), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2390 (.Q(w2519), .D(w31), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2391 (.Q(w2391), .D(w33), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2392 (.nZ(w2531), .A(w2389) );
	vdp_or g2393 (.Z(w2399), .A(w33), .B(w2391) );
	vdp_sr_bit g2394 (.Q(w2408), .D(w2410), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_sr_bit g2395 (.Q(w2532), .D(w2521), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2396 (.nZ(w2463), .A(w2532) );
	vdp_or g2397 (.Z(w2387), .A(w2391), .B(w2390) );
	vdp_sr_bit g2398 (.Q(w2390), .D(w540), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2399 (.Q(w2388), .D(w30), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2400 (.Q(w2523), .D(w2388), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2401 (.Q(w2522), .D(w2400), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2402 (.Q(w2517), .D(w2519), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2403 (.Q(w2534), .D(w2539), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_not g2404 (.nZ(w2513), .A(w2581) );
	vdp_not g2405 (.nZ(w2411), .A(VRAM128k) );
	vdp_sr_bit g2406 (.Q(w2400), .D(VRAM_REFRESH), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2407 (.nZ(w2471), .A(w2386) );
	vdp_not g2408 (.nZ(w2537), .A(w2524) );
	vdp_not g2409 (.nZ(w2406), .A(w2398) );
	vdp_oai21 g2410 (.Z(w2386), .B(w2406), .A1(w2537), .A2(w2525) );
	vdp_or g2411 (.Z(w2398), .A(w2531), .B(w2530) );
	vdp_or g2412 (.Z(w2529), .A(w2390), .B(w540) );
	vdp_not g2413 (.nZ(w2538), .A(w2392) );
	vdp_not g2414 (.nZ(w2573), .A(w2539) );
	vdp_dlatch_inv g2415 (.nQ(w2539), .D(w3), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2416 (.nQ(w2533), .D(w2407), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g2417 (.nQ(w2407), .D(w2534), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g2418 (.nQ(w2389), .D(w2387), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2419 (.nQ(w2530), .D(w2389), .C(HCLK2), .nC(nHCLK2) );
	vdp_dlatch_inv g2420 (.nQ(w2527), .D(w2526), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2421 (.nQ(w2524), .D(w2523), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2422 (.nQ(w2525), .D(w2524), .C(HCLK2), .nC(nHCLK2) );
	vdp_aon22 g2423 (.Z(nCAS1), .A1(w2407), .B1(w2396), .B2(1'b1), .A2(w2532) );
	vdp_and3 g2424 (.Z(nWE1), .A(w2395), .B(w2536), .C(w2396) );
	vdp_and3 g2425 (.Z(nWE0), .A(w2396), .B(w2395), .C(w2535) );
	vdp_aoi222 g2426 (.Z(w2528), .A1(1'b1), .B1(w2393), .B2(1'b1), .A2(w88), .C1(w2398), .C2(w2396) );
	vdp_aon333 g2427 (.Z(nOE1), .A1(w2471), .A2(w2534), .A3(w2396), .B1(w2527), .B2(w2527), .B3(w2538), .C1(w2527), .C2(w2527), .C3(w2393) );
	vdp_or3 g2428 (.Z(w2526), .A(w2521), .B(w2523), .C(w2388) );
	vdp_sr_bit g2429 (.Q(w2393), .D(w2573), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_dlatch_inv g2430 (.nQ(w2395), .D(w2393), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g2431 (.nQ(w2520), .D(w2395), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g2432 (.nQ(w2396), .D(w2394), .C(DCLK1), .nC(nDCLK1) );
	vdp_not g2433 (.nZ(w2394), .A(w2520) );
	vdp_nand g2434 (.Z(w2607), .A(w2520), .B(w2393) );
	vdp_nand g2435 (.Z(w2606), .A(w2393), .B(w2533) );
	vdp_nand g2436 (.Z(w2402), .A(w2534), .B(1'b1) );
	vdp_aoi33 g2437 (.Z(w2587), .A1(w2517), .A2(w32), .A3(w32), .B1(w2413), .B2(w2414), .B3(w3) );
	vdp_and g2438 (.Z(w2409), .A(w2396), .B(w2395) );
	vdp_not g2439 (.nZ(w2403), .A(w2464) );
	vdp_comp_strong g2440 (.nZ(w2420), .Z(w2419), .A(w2426) );
	vdp_comp_strong g2441 (.nZ(w2486), .Z(w2508), .A(w2509) );
	vdp_comp_strong g2442 (.nZ(w2421), .Z(w2465), .A(w2509) );
	vdp_comp_strong g2443 (.nZ(w2469), .Z(w2468), .A(w2426) );
	vdp_comp_strong g2444 (.nZ(w2427), .Z(w2470), .A(w2423) );
	vdp_comp_strong g2445 (.nZ(w2473), .Z(w2514), .A(w2423) );
	vdp_not g2446 (.nZ(w2429), .A(w2393) );
	vdp_not g2447 (.nZ(w2414), .A(w32) );
	vdp_not g2448 (.nZ(w2413), .A(w34) );
	vdp_comp_strong g2449 (.nZ(w2467), .Z(w6538), .A(w2409) );
	vdp_comp_strong g2450 (.nZ(w2404), .Z(w2510), .A(w2409) );
	vdp_or g2451 (.Z(w2521), .A(w2400), .B(w2522) );
	vdp_and g2452 (.Z(w2410), .A(VRAM128k), .B(HCLK1) );
	vdp_comp_we g2453 (.nZ(w2511), .Z(w2512), .A(w88) );
	vdp_comp_we g2454 (.nZ(w2422), .Z(w2585), .A(w2430) );
	vdp_not g2455 (.nZ(w2586), .A(w2464) );
	vdp_not g2456 (.nZ(w2425), .A(w2607) );
	vdp_not g2457 (.nZ(w6543), .A(w2606) );
	vdp_not g2458 (.nZ(w6544), .A(w2402) );
	vdp_comp_we g2459 (.nZ(w6545), .Z(w2516), .A(M5) );
	vdp_comp_we g2460 (.nZ(w2472), .Z(w2428), .A(VRAM128k) );
	vdp_and g2461 (.Z(w2412), .A(w98), .B(w3) );
	vdp_and g2462 (.Z(w2423), .A(w3), .B(HCLK1) );
	vdp_and g2463 (.Z(w2426), .A(HCLK2), .B(w2518) );
	vdp_and g2464 (.Z(w2509), .A(w3), .B(HCLK1) );
	vdp_oai21 g2465 (.Z(w2581), .A1(HCLK2), .A2(w2411), .B(DCLK1) );
	vdp_notif0 g2466 (.nZ(AD_DATA[0]), .A(w2417), .nE(w2403) );
	vdp_aon22 g2467 (.Z(nYS), .A1(VRAMA[16]), .A2(w2512), .B1(w2511), .B2(w2569) );
	vdp_aon22 g2468 (.Z(w2553), .A1(VRAMA[15]), .B1(w2511), .A2(w2512), .B2(w2492) );
	vdp_aon22 g2469 (.Z(w2551), .A1(VRAMA[14]), .B1(w2511), .A2(w2512), .B2(w2378) );
	vdp_aon22 g2470 (.Z(w2603), .A1(VRAMA[6]), .B1(w2511), .A2(w2512), .B2(w2552) );
	vdp_aon22 g2471 (.Z(w2491), .A1(VRAMA[7]), .B1(w2511), .A2(w2512), .B2(w2370) );
	vdp_aon22 g2472 (.Z(w2570), .A1(VRAMA[13]), .B1(w2511), .A2(w2512), .B2(w2385) );
	vdp_aon22 g2473 (.Z(w2592), .A1(VRAMA[5]), .B1(w2511), .A2(w2512), .B2(w2589) );
	vdp_aon22 g2474 (.Z(w2556), .A1(VRAMA[12]), .B1(w2511), .A2(w2512), .B2(w2453) );
	vdp_aon22 g2475 (.Z(w2605), .A1(VRAMA[4]), .B1(w2511), .A2(w2512), .B2(w2460) );
	vdp_aon22 g2476 (.Z(w2555), .A1(VRAMA[11]), .B1(w2511), .A2(w2512), .B2(w2596) );
	vdp_aon22 g2477 (.Z(w2597), .A1(VRAMA[3]), .B1(w2511), .A2(w2512), .B2(w2590) );
	vdp_aon22 g2478 (.Z(w2571), .A1(VRAMA[10]), .B1(w2511), .A2(w2512), .B2(w2504) );
	vdp_aon22 g2479 (.Z(w2595), .A1(VRAMA[2]), .B1(w2511), .A2(w2512), .B2(w2449) );
	vdp_aon22 g2480 (.Z(w2415), .A1(VRAMA[8]), .B1(w2511), .A2(w2512), .B2(w2418) );
	vdp_aon22 g2481 (.Z(w2593), .A1(VRAMA[0]), .B1(w2511), .A2(w2512), .B2(w2441) );
	vdp_aon22 g2482 (.Z(w2594), .A1(VRAMA[9]), .B1(w2511), .A2(w2512), .B2(w2487) );
	vdp_aon22 g2483 (.Z(w2604), .A1(VRAMA[1]), .B1(w2511), .A2(w2512), .B2(w2445) );
	vdp_notif0 g2484 (.nZ(AD_DATA[1]), .A(w2436), .nE(w2403) );
	vdp_notif0 g2485 (.nZ(AD_DATA[2]), .A(w2489), .nE(w2403) );
	vdp_notif0 g2486 (.nZ(AD_DATA[3]), .A(w2446), .nE(w2403) );
	vdp_notif0 g2487 (.nZ(AD_DATA[5]), .A(w2384), .nE(w2403) );
	vdp_notif0 g2488 (.nZ(AD_DATA[4]), .A(w2466), .nE(w2403) );
	vdp_notif0 g2489 (.nZ(AD_DATA[6]), .A(w2379), .nE(w2403) );
	vdp_notif0 g2490 (.nZ(AD_DATA[7]), .A(w2377), .nE(w2403) );
	vdp_slatch g2491 (.nQ(w2417), .D(w2416), .nC(w2404), .C(w2510) );
	vdp_slatch g2492 (.nQ(w2436), .D(w2435), .nC(w2404), .C(w2510) );
	vdp_slatch g2493 (.nQ(w2489), .D(w2443), .nC(w2404), .C(w2510) );
	vdp_slatch g2494 (.nQ(w2446), .D(w2447), .nC(w2404), .C(w2510) );
	vdp_slatch g2495 (.nQ(w2466), .D(w2401), .nC(w2404), .C(w2510) );
	vdp_slatch g2496 (.nQ(w2384), .D(w2609), .nC(w2404), .C(w2510) );
	vdp_slatch g2497 (.nQ(w2379), .D(w2455), .nC(w2404), .C(w2510) );
	vdp_slatch g2498 (.nQ(w2377), .D(w2554), .nC(w2404), .C(w2510) );
	vdp_slatch g2499 (.nQ(w2372), .D(w2371), .nC(w2467), .C(w6538) );
	vdp_slatch g2500 (.nQ(w2458), .D(w2454), .nC(w2467), .C(w6538) );
	vdp_slatch g2501 (.nQ(w2495), .D(w2582), .nC(w2467), .C(w6538) );
	vdp_slatch g2502 (.nQ(w2496), .D(w2383), .nC(w2467), .C(w6538) );
	vdp_slatch g2503 (.nQ(w2557), .D(w2456), .nC(w2467), .C(w6538) );
	vdp_slatch g2504 (.nQ(w2450), .D(w2448), .nC(w2467), .C(w6538) );
	vdp_slatch g2505 (.nQ(w2444), .D(w2490), .nC(w2467), .C(w6538) );
	vdp_slatch g2506 (.nQ(w2474), .D(w2572), .nC(w2467), .C(w6538) );
	vdp_slatch g2507 (.Q(w2418), .D(w2477), .nC(w2420), .C(w2419) );
	vdp_slatch g2508 (.Q(w2487), .D(w2599), .nC(w2420), .C(w2419) );
	vdp_slatch g2509 (.Q(w2596), .D(w2560), .nC(w2420), .C(w2419) );
	vdp_slatch g2510 (.Q(w2504), .D(w2488), .nC(w2420), .C(w2419) );
	vdp_slatch g2511 (.Q(w2385), .D(w2476), .nC(w2420), .C(w2419) );
	vdp_slatch g2512 (.Q(w2453), .D(w2561), .nC(w2420), .C(w2419) );
	vdp_slatch g2513 (.Q(w2492), .D(w2564), .nC(w2420), .C(w2419) );
	vdp_slatch g2514 (.Q(w2378), .D(w2475), .nC(w2420), .C(w2419) );
	vdp_slatch g2515 (.nQ(w2563), .D(w355), .nC(w2486), .C(w2508) );
	vdp_slatch g2516 (.nQ(w2565), .D(RD_DATA[6]), .nC(w2486), .C(w2508) );
	vdp_slatch g2517 (.nQ(w2562), .D(RD_DATA[5]), .nC(w2486), .C(w2508) );
	vdp_slatch g2518 (.nQ(w2601), .D(RD_DATA[4]), .nC(w2486), .C(w2508) );
	vdp_slatch g2519 (.nQ(w2559), .D(w321), .nC(w2486), .C(w2508) );
	vdp_slatch g2520 (.nQ(w2602), .D(RD_DATA[2]), .nC(w2486), .C(w2508) );
	vdp_slatch g2521 (.nQ(w2600), .D(RD_DATA[0]), .nC(w2486), .C(w2508) );
	vdp_slatch g2522 (.nQ(w2558), .D(RD_DATA[1]), .nC(w2486), .C(w2508) );
	vdp_notif0 g2523 (.nZ(w355), .A(w2372), .nE(w2586) );
	vdp_notif0 g2524 (.nZ(RD_DATA[6]), .A(w2458), .nE(w2586) );
	vdp_notif0 g2525 (.nZ(RD_DATA[5]), .A(w2495), .nE(w2586) );
	vdp_notif0 g2526 (.nZ(RD_DATA[4]), .A(w2496), .nE(w2586) );
	vdp_notif0 g2527 (.nZ(w321), .A(w2557), .nE(w2586) );
	vdp_notif0 g2528 (.nZ(RD_DATA[2]), .A(w2450), .nE(w2586) );
	vdp_notif0 g2529 (.nZ(RD_DATA[1]), .A(w2444), .nE(w2586) );
	vdp_notif0 g2530 (.nZ(RD_DATA[0]), .A(w2474), .nE(w2586) );
	vdp_slatch g2531 (.nQ(w2575), .D(AD_DATA[7]), .nC(w2421), .C(w2465) );
	vdp_slatch g2532 (.nQ(w2574), .D(AD_DATA[6]), .nC(w2421), .C(w2465) );
	vdp_slatch g2533 (.nQ(w2598), .D(AD_DATA[5]), .nC(w2421), .C(w2465) );
	vdp_slatch g2534 (.nQ(w2577), .D(AD_DATA[3]), .nC(w2421), .C(w2465) );
	vdp_slatch g2535 (.nQ(w2578), .D(AD_DATA[2]), .nC(w2421), .C(w2465) );
	vdp_slatch g2536 (.nQ(w2580), .D(AD_DATA[1]), .nC(w2421), .C(w2465) );
	vdp_slatch g2537 (.nQ(w2579), .D(AD_DATA[0]), .nC(w2421), .C(w2465) );
	vdp_slatch g2538 (.Q(w2376), .D(w2485), .nC(w2469), .C(w2468) );
	vdp_slatch g2539 (.Q(w2382), .D(w2484), .nC(w2469), .C(w2468) );
	vdp_slatch g2540 (.Q(w2457), .D(w2483), .nC(w2469), .C(w2468) );
	vdp_slatch g2541 (.Q(w2583), .D(w2480), .nC(w2469), .C(w2468) );
	vdp_slatch g2542 (.Q(w2507), .D(w2481), .nC(w2469), .C(w2468) );
	vdp_slatch g2543 (.Q(w2442), .D(w2479), .nC(w2469), .C(w2468) );
	vdp_slatch g2544 (.Q(w2494), .D(w2375), .nC(w2427), .C(w2470) );
	vdp_slatch g2545 (.Q(w2588), .D(w2381), .nC(w2427), .C(w2470) );
	vdp_slatch g2546 (.Q(w2567), .D(w2434), .nC(w2427), .C(w2470) );
	vdp_slatch g2547 (.Q(w2498), .D(w2433), .nC(w2427), .C(w2470) );
	vdp_slatch g2548 (.Q(w2505), .D(w2506), .nC(w2427), .C(w2470) );
	vdp_slatch g2549 (.Q(w2584), .D(w2439), .nC(w2427), .C(w2470) );
	vdp_slatch g2550 (.Q(w2503), .D(w2405), .nC(w2427), .C(w2470) );
	vdp_slatch g2551 (.Q(w2591), .D(w2440), .nC(w2427), .C(w2470) );
	vdp_slatch g2552 (.Q(w2515), .D(w2438), .nC(w2473), .C(w2514) );
	vdp_slatch g2553 (.Q(w2502), .D(w2613), .nC(w2473), .C(w2514) );
	vdp_slatch g2554 (.Q(w2451), .D(w2432), .nC(w2473), .C(w2514) );
	vdp_slatch g2555 (.Q(w2499), .D(w2608), .nC(w2473), .C(w2514) );
	vdp_slatch g2556 (.Q(w2461), .D(w2380), .nC(w2473), .C(w2514) );
	vdp_slatch g2557 (.Q(w2497), .D(w2431), .nC(w2473), .C(w2514) );
	vdp_slatch g2558 (.Q(w2459), .D(w2374), .nC(w2473), .C(w2514) );
	vdp_slatch g2559 (.Q(w2493), .D(w2373), .nC(w2473), .C(w2514) );
	vdp_sr_bit g2560 (.Q(w2430), .D(w32), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2561 (.nZ(w2619), .A(w116) );
	vdp_not g2562 (.nZ(w2500), .A(w2501) );
	vdp_not g2563 (.nZ(w6546), .A(M5) );
	vdp_not g2564 (.nZ(w2437), .A(w2429) );
	vdp_not g2565 (.nZ(w2392), .A(w2437) );
	vdp_aoi21 g2566 (.Z(w2501), .B(w2568), .A2(VRAMA[9]), .A1(w6546) );
	vdp_aoi22 g2567 (.Z(w2599), .A1(w2444), .B1(w2422), .B2(w2558), .A2(w2585) );
	vdp_aoi22 g2568 (.Z(w2560), .A1(w2557), .B1(w2422), .B2(w2559), .A2(w2585) );
	vdp_aoi22 g2569 (.Z(w2488), .A1(w2450), .B1(w2422), .B2(w2602), .A2(w2585) );
	vdp_aoi22 g2570 (.Z(w2476), .A1(w2495), .B1(w2422), .B2(w2562), .A2(w2585) );
	vdp_aoi22 g2571 (.Z(w2561), .A1(w2496), .B1(w2422), .B2(w2601), .A2(w2585) );
	vdp_aoi22 g2572 (.Z(w2564), .A1(w2372), .B1(w2422), .B2(w2563), .A2(w2585) );
	vdp_aoi22 g2573 (.Z(w2475), .A1(w2458), .B1(w2422), .B2(w2565), .A2(w2585) );
	vdp_slatch g2574 (.Q(w2424), .D(w2478), .nC(w2469), .C(w2468) );
	vdp_slatch g2575 (.nQ(w2576), .D(AD_DATA[4]), .nC(w2421), .C(w2465) );
	vdp_slatch g2576 (.Q(w2452), .D(w2482), .nC(w2469), .C(w2468) );
	vdp_aoi22 g2577 (.Z(w2478), .A1(w2417), .B1(w2422), .B2(w2579), .A2(w2585) );
	vdp_aoi22 g2578 (.Z(w2479), .A1(w2436), .B1(w2422), .B2(w2580), .A2(w2585) );
	vdp_aoi22 g2579 (.Z(w2480), .A1(w2489), .B1(w2422), .B2(w2578), .A2(w2585) );
	vdp_aoi22 g2580 (.Z(w2481), .A1(w2446), .B1(w2422), .B2(w2577), .A2(w2585) );
	vdp_aoi22 g2581 (.Z(w2482), .A1(w2466), .B1(w2422), .B2(w2576), .A2(w2585) );
	vdp_aoi22 g2582 (.Z(w2483), .A1(w2384), .B1(w2422), .B2(w2598), .A2(w2585) );
	vdp_aoi22 g2583 (.Z(w2485), .A1(w2377), .B1(w2422), .B2(w2575), .A2(w2585) );
	vdp_aoi22 g2584 (.Z(w2484), .A1(w2379), .B1(w2422), .B2(w2574), .A2(w2585) );
	vdp_aon22 g2585 (.Z(w2440), .A1(VRAMA[2]), .B1(w6545), .B2(VRAMA[1]), .A2(w2516) );
	vdp_aon22 g2586 (.Z(w2439), .A1(VRAMA[3]), .B1(w6545), .B2(VRAMA[2]), .A2(w2516) );
	vdp_aon22 g2587 (.Z(w2405), .A1(VRAMA[4]), .B1(w6545), .B2(VRAMA[3]), .A2(w2516) );
	vdp_aon22 g2588 (.Z(w2506), .A1(VRAMA[5]), .B1(w6545), .B2(VRAMA[4]), .A2(w2516) );
	vdp_aon22 g2589 (.Z(w2433), .A1(VRAMA[6]), .B1(w6545), .B2(VRAMA[5]), .A2(w2516) );
	vdp_aon22 g2590 (.Z(w2434), .A1(VRAMA[7]), .B1(w6545), .B2(VRAMA[6]), .A2(w2516) );
	vdp_aon22 g2591 (.Z(w2381), .A1(VRAMA[8]), .B1(w6545), .B2(VRAMA[7]), .A2(w2516) );
	vdp_aon22 g2592 (.Z(w2375), .A1(VRAMA[9]), .B1(w6545), .B2(VRAMA[8]), .A2(w2516) );
	vdp_and g2593 (.Z(w2568), .A(VRAMA[1]), .B(M5) );
	vdp_aon22 g2594 (.Z(w2373), .A1(w2566), .B1(w2472), .B2(VRAMA[15]), .A2(w2428) );
	vdp_aon22 g2595 (.Z(w2374), .A1(VRAMA[15]), .B1(w2472), .B2(VRAMA[14]), .A2(w2428) );
	vdp_aon22 g2596 (.Z(w2380), .A1(VRAMA[14]), .B1(w2472), .B2(VRAMA[13]), .A2(w2428) );
	vdp_aon22 g2597 (.Z(w2608), .A1(VRAMA[12]), .B1(w2472), .B2(VRAMA[11]), .A2(w2428) );
	vdp_aon22 g2598 (.Z(w2431), .A1(VRAMA[13]), .B1(w2472), .B2(VRAMA[12]), .A2(w2428) );
	vdp_aon22 g2599 (.Z(w2432), .A1(VRAMA[11]), .B1(w2472), .B2(VRAMA[10]), .A2(w2428) );
	vdp_aon22 g2600 (.Z(w2613), .A1(VRAMA[10]), .B1(w2472), .B2(w2500), .A2(w2428) );
	vdp_aon22 g2601 (.Z(w2438), .A1(w2568), .B1(w2472), .B2(VRAMA[0]), .A2(w2428) );
	vdp_aon22 g2602 (.Z(w2566), .A1(w2619), .B1(w116), .B2(w82), .A2(VRAMA[16]) );
	vdp_aon222 g2603 (.Z(w2441), .A1(w2425), .A2(w2424), .B1(w6543), .B2(w2591), .C1(w6544), .C2(w2515) );
	vdp_aon222 g2604 (.Z(w2445), .A1(w2425), .A2(w2442), .B1(w6543), .B2(w2584), .C1(w6544), .C2(w2502) );
	vdp_aon222 g2605 (.Z(w2449), .A1(w2425), .A2(w2583), .B1(w6543), .B2(w2503), .C1(w6544), .C2(w2451) );
	vdp_aon222 g2606 (.Z(w2590), .A1(w2425), .A2(w2507), .B1(w6543), .B2(w2505), .C1(w6544), .C2(w2499) );
	vdp_aon222 g2607 (.Z(w2460), .A1(w2425), .A2(w2452), .B1(w6543), .B2(w2498), .C1(w6544), .C2(w2497) );
	vdp_aon222 g2608 (.Z(w2589), .A1(w2425), .A2(w2457), .B1(w6543), .B2(w2567), .C1(w6544), .C2(w2461) );
	vdp_aon222 g2609 (.Z(w2552), .A1(w2425), .A2(w2382), .B1(w6543), .B2(w2588), .C1(w6544), .C2(w2459) );
	vdp_aon222 g2610 (.Z(w2370), .A1(w2425), .A2(w2376), .B1(w6543), .B2(w2494), .C1(w6544), .C2(w2493) );
	vdp_dlatch_inv g2611 (.nQ(w2518), .D(w2587), .C(HCLK1), .nC(nHCLK1) );
	vdp_comp_we g2612 (.Z(w2462), .A(w2520) );
	vdp_aon22 g2613 (.Z(nRAS1), .A1(1'b1), .B1(w2463), .B2(w2407), .A2(w2462) );
	vdp_aoi22 g2614 (.Z(w2477), .A1(w2474), .B1(w2422), .B2(w2600), .A2(w2585) );
	vdp_and g2615 (.Z(w2540), .B(w2618), .A(DCLK2) );
	vdp_nor g2616 (.Z(w2614), .A(w2542), .B(RES) );
	vdp_sr_bit g2617 (.Q(w2542), .D(w2614), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_dlatch_inv g2618 (.nQ(w2615), .D(w2543), .C(DCLK1), .nC(nDCLK1) );
	vdp_and g2619 (.Z(w2616), .A(DCLK2), .B(w2615) );
	vdp_dlatch_inv g2620 (.nQ(w2618), .D(w2542), .C(DCLK1), .nC(nDCLK1) );
	vdp_not g2621 (.nZ(w2546), .A(w2548) );
	vdp_not g2622 (.nZ(w2545), .A(w2617) );
	vdp_neg_dff g2623 (.Q(w2548), .C(DCLK1), .D(1'b1), .R(w2540) );
	vdp_not g2624 (.A(w2542), .nZ(w2543) );
	vdp_neg_dff g2625 (.Q(w2617), .R(w2616), .C(DCLK1), .D(1'b1) );
	vdp_sr_bit g2626 (.Q(w2694), .D(w2686), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2627 (.Q(w2690), .D(w2689), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2628 (.Q(w2878), .D(w2690), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2629 (.Q(w2708), .D(w2878), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2630 (.Q(w2663), .D(RD_DATA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2631 (.Q(w2664), .D(RD_DATA[2]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2632 (.Q(w2665), .D(w321), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2633 (.Q(w2857), .D(w2881), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2634 (.Q(w2881), .D(w2882), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2635 (.Q(w2882), .D(w2883), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2636 (.Q(w2883), .D(w2884), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2637 (.Q(w2884), .D(w2885), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2638 (.Q(w2885), .D(w2886), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2639 (.Q(w2886), .D(w2887), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2640 (.Q(w2887), .D(w17), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2641 (.Q(w2672), .D(w2700), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2642 (.Q(w2670), .D(w2890), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2643 (.Q(w2914), .D(w2892), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2644 (.Q(w2892), .D(w2646), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2645 (.Q(w2646), .D(w96), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2646 (.Q(w2621), .D(w2620), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2647 (.Q(w2626), .D(w2760), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2648 (.Q(w2684), .D(w2872), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2649 (.Q(w2688), .D(w2889), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2650 (.Q(w2704), .D(w2696), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2651 (.Q(w2620), .D(w2699), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2652 (.Q(w2725), .D(w2702), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2653 (.Q(w2724), .D(w2761), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2654 (.Q(PLANE_A_PRIO), .D(w2716), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2655 (.Q(PLANE_B_PRIO), .D(w2717), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2656 (.Q(w2680), .D(w2718), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2657 (.Q(w2723), .D(w2722), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2658 (.Q(w2642), .D(w2721), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2659 (.Q(w2721), .D(COL[7]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2660 (.Q(w2643), .D(w2916), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2661 (.Q(w2916), .D(w117), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2662 (.Q(w2734), .D(w2707), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2663 (.Q(w2720), .D(w2719), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2664 (.Q(SPR_PRIO), .D(w2864), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2665 (.Q(w2731), .D(w173), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2666 (.Q(w2730), .D(w172), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2667 (.Q(w2635), .D(w2651), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2668 (.Q(w2640), .D(w2652), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2669 (.Q(w2637), .D(w2662), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2670 (.Q(w2628), .D(w2653), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2671 (.Q(w2647), .D(w2659), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2672 (.Q(w2627), .D(w2654), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2673 (.Q(w2622), .D(w2757), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2674 (.Q(w2632), .D(w2655), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2675 (.Q(w2638), .D(w2649), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_slatch g2676 (.nQ(w2912), .D(w2651), .C(w2648), .nC(w2645) );
	vdp_slatch g2677 (.nQ(w2913), .D(w2649), .C(w2648), .nC(w2645) );
	vdp_slatch g2678 (.nQ(w2911), .D(w2652), .C(w2648), .nC(w2645) );
	vdp_slatch g2679 (.nQ(w2910), .D(w2662), .C(w2648), .nC(w2645) );
	vdp_slatch g2680 (.nQ(w2909), .D(w2653), .C(w2648), .nC(w2645) );
	vdp_slatch g2681 (.nQ(w2908), .D(w2659), .C(w2648), .nC(w2645) );
	vdp_slatch g2682 (.nQ(w2907), .D(w2654), .C(w2648), .nC(w2645) );
	vdp_slatch g2683 (.nQ(w2906), .D(w2757), .C(w2648), .nC(w2645) );
	vdp_slatch g2684 (.nQ(w2905), .D(w2655), .C(w2648), .nC(w2645) );
	vdp_slatch g2685 (.Q(w2706), .D(REG_BUS[7]), .nC(w2683), .C(w2693) );
	vdp_slatch g2686 (.Q(w2703), .D(REG_BUS[5]), .nC(w2683), .C(w2693) );
	vdp_slatch g2687 (.Q(w2695), .D(REG_BUS[4]), .nC(w2683), .C(w2693) );
	vdp_slatch g2688 (.Q(w2691), .D(REG_BUS[3]), .nC(w2683), .C(w2693) );
	vdp_slatch g2689 (.Q(w2687), .D(REG_BUS[2]), .nC(w2683), .C(w2693) );
	vdp_slatch g2690 (.Q(w2877), .D(REG_BUS[1]), .nC(w2683), .C(w2693) );
	vdp_slatch g2691 (.Q(w2685), .D(REG_BUS[0]), .nC(w2683), .C(w2693) );
	vdp_slatch g2692 (.Q(w2850), .D(REG_BUS[6]), .nC(w2683), .C(w2693) );
	vdp_aon2222 g2693 (.Z(w2827), .B2(w2766), .B1(w2771), .A2(w2900), .A1(w2766), .D2(w2762), .D1(w2771), .C2(w2771), .C1(HIGHLIGHT) );
	vdp_aon22 g2694 (.Z(w2792), .B2(w2762), .B1(w2776), .A2(w2901), .A1(w2767) );
	vdp_aon22 g2695 (.Z(w2797), .B2(w2762), .B1(w2772), .A2(w2900), .A1(w2767) );
	vdp_not g2696 (.nZ(w2780), .A(w2826) );
	vdp_not g2697 (.nZ(w2774), .A(w2775) );
	vdp_not g2698 (.nZ(w2779), .A(w2778) );
	vdp_not g2699 (.nZ(w2798), .A(w2827) );
	vdp_not g2700 (.nZ(w2791), .A(w2784) );
	vdp_comp_we g2701 (.Z(w2766), .A(w2670) );
	vdp_not g2702 (.nZ(w2861), .A(w2819) );
	vdp_not g2703 (.nZ(w2822), .A(w2820) );
	vdp_not g2704 (.nZ(w2823), .A(w2824) );
	vdp_not g2705 (.nZ(w2787), .A(HIGHLIGHT) );
	vdp_sr_bit g2706 (.Q(SHADOW), .D(w2643), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2707 (.Q(w2824), .D(w2641), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2708 (.Q(HIGHLIGHT), .D(w2642), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2709 (.Q(w2819), .D(w2821), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2710 (.Q(w2820), .D(w2666), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g2711 (.Z(w2896), .A(w2823), .B(w2861), .C(w2820) );
	vdp_and3 g2712 (.Z(w2898), .A(w2822), .B(w2824), .C(w2861) );
	vdp_and3 g2713 (.Z(w2897), .A(w2823), .B(w2861), .C(w2822) );
	vdp_and3 g2714 (.Z(w2785), .A(w2861), .B(w2820), .C(w2824) );
	vdp_and3 g2715 (.Z(w2783), .A(w2823), .B(w2819), .C(w2822) );
	vdp_and3 g2716 (.Z(w2781), .A(w2819), .B(w2820), .C(w2824) );
	vdp_and3 g2717 (.Z(w2899), .A(w2823), .B(w2820), .C(w2819) );
	vdp_and3 g2718 (.Z(w2782), .A(w2822), .B(w2824), .C(w2819) );
	vdp_sr_bit g2719 (.Q(w2778), .D(w2825), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2720 (.Q(w2775), .D(w2631), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2721 (.Q(w2826), .D(w2667), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g2722 (.Z(w2777), .A(w2779), .B(w2780), .C(w2774) );
	vdp_and3 g2723 (.Z(w2776), .A(w2774), .B(w2778), .C(w2780) );
	vdp_and3 g2724 (.Z(w2901), .A(w2779), .B(w2780), .C(w2775) );
	vdp_and3 g2725 (.Z(w2772), .A(w2780), .B(w2775), .C(w2778) );
	vdp_and3 g2726 (.Z(w2773), .A(w2774), .B(w2778), .C(w2826) );
	vdp_and3 g2727 (.Z(w2770), .A(w2779), .B(w2826), .C(w2774) );
	vdp_and3 g2728 (.Z(w2900), .A(w2779), .B(w2775), .C(w2826) );
	vdp_and3 g2729 (.Z(w2771), .A(w2826), .B(w2775), .C(w2778) );
	vdp_not g2730 (.nZ(w2860), .A(w2915) );
	vdp_not g2731 (.nZ(w2815), .A(w2817) );
	vdp_not g2732 (.nZ(w2816), .A(w2818) );
	vdp_sr_bit g2733 (.Q(w2817), .D(w2856), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2734 (.Q(w2818), .D(w2854), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2735 (.Q(w2915), .D(w2629), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g2736 (.Z(w2769), .A(w2816), .B(w2860), .C(w2815) );
	vdp_and3 g2737 (.Z(w2768), .A(w2815), .B(w2818), .C(w2860) );
	vdp_and3 g2738 (.A(w2816), .B(w2860), .C(w2817), .Z(w2765) );
	vdp_and3 g2739 (.Z(w2902), .A(w2860), .B(w2817), .C(w2818) );
	vdp_and3 g2740 (.Z(w2764), .A(w2816), .B(w2915), .C(w2815) );
	vdp_and3 g2741 (.Z(w2904), .A(w2815), .B(w2818), .C(w2915) );
	vdp_and3 g2742 (.Z(w2859), .A(w2915), .B(w2817), .C(w2818) );
	vdp_and3 g2743 (.Z(w2903), .A(w2816), .B(w2817), .C(w2915) );
	vdp_aon22 g2744 (.nZ(w2849), .B2(w2762), .B1(w2903), .A2(w2904), .A1(HIGHLIGHT) );
	vdp_aon22 g2745 (.nZ(w2814), .B2(w2762), .B1(w2764), .A2(w2768), .A1(HIGHLIGHT) );
	vdp_aon22 g2746 (.nZ(w2848), .B2(HIGHLIGHT), .B1(w2769), .A2(w2859), .A1(w2767) );
	vdp_and g2747 (.nZ(w2813), .B(HIGHLIGHT), .A(w2764) );
	vdp_and g2748 (.nZ(w2847), .B(HIGHLIGHT), .A(w2903) );
	vdp_and g2749 (.nZ(w2846), .B(HIGHLIGHT), .A(w2765) );
	vdp_aon22 g2750 (.nZ(w2845), .B2(w2766), .B1(w2904), .A2(w2764), .A1(w2766) );
	vdp_aon22 g2751 (.nZ(w2844), .B2(w2762), .B1(w2904), .A2(w2902), .A1(HIGHLIGHT) );
	vdp_aon2222 g2752 (.Z(w2828), .B2(w2766), .B1(w2859), .A2(w2903), .A1(w2766), .D2(w2762), .D1(w2859), .C2(w2859), .C1(HIGHLIGHT) );
	vdp_aon22 g2753 (.Z(w2811), .B2(w2762), .B1(w2768), .A2(w2765), .A1(w2767) );
	vdp_aon22 g2754 (.Z(w2808), .B2(w2762), .B1(w2902), .A2(w2903), .A1(w2767) );
	vdp_and g2755 (.Z(w2812), .B(w2904), .A(w2767) );
	vdp_and g2756 (.Z(w2807), .B(w2767), .A(w2902) );
	vdp_and g2757 (.Z(w2809), .B(w2768), .A(w2767) );
	vdp_aon22 g2758 (.Z(w2806), .B2(w2766), .B1(w2902), .A2(w2765), .A1(w2766) );
	vdp_aon22 g2759 (.Z(w2805), .B2(w2762), .B1(w2765), .A2(w2764), .A1(w2767) );
	vdp_aon2222 g2760 (.Z(w2843), .B2(w2766), .B1(w2768), .A2(w2769), .A1(w2766), .D2(w2762), .D1(w2769), .C2(w2769), .C1(w2767) );
	vdp_not g2761 (.nZ(w2810), .A(w2828) );
	vdp_aon22 g2762 (.nZ(w2842), .B2(w2762), .B1(w2900), .A2(w2773), .A1(HIGHLIGHT) );
	vdp_aon22 g2763 (.nZ(w2841), .B2(w2762), .B1(w2770), .A2(w2776), .A1(HIGHLIGHT) );
	vdp_aon22 g2764 (.nZ(w2804), .B2(HIGHLIGHT), .B1(w2777), .A2(w2771), .A1(w2767) );
	vdp_and g2765 (.nZ(w2803), .B(HIGHLIGHT), .A(w2770) );
	vdp_and g2766 (.nZ(w2802), .B(HIGHLIGHT), .A(w2900) );
	vdp_and g2767 (.nZ(w2801), .B(HIGHLIGHT), .A(w2901) );
	vdp_aon22 g2768 (.nZ(w2800), .B2(w2766), .B1(w2773), .A2(w2770), .A1(w2766) );
	vdp_aon22 g2769 (.nZ(w2799), .B2(w2762), .B1(w2773), .A2(w2772), .A1(HIGHLIGHT) );
	vdp_and g2770 (.Z(w2796), .B(w2773), .A(w2767) );
	vdp_and g2771 (.Z(w2893), .B(w2767), .A(w2772) );
	vdp_and g2772 (.Z(w2795), .B(w2776), .A(w2767) );
	vdp_aon22 g2773 (.Z(w2794), .B2(w2766), .B1(w2772), .A2(w2901), .A1(w2766) );
	vdp_aon22 g2774 (.Z(w2793), .B2(w2762), .B1(w2901), .A2(w2770), .A1(w2767) );
	vdp_aon2222 g2775 (.Z(w2894), .B2(w2766), .B1(w2776), .A2(w2777), .A1(w2766), .D2(w2762), .D1(w2777), .C2(w2777), .C1(w2767) );
	vdp_aon22 g2776 (.nZ(w2790), .B2(w2762), .B1(w2899), .A2(w2782), .A1(HIGHLIGHT) );
	vdp_aon22 g2777 (.nZ(w2840), .B2(w2762), .B1(w2783), .A2(w2898), .A1(HIGHLIGHT) );
	vdp_aon22 g2778 (.nZ(w2836), .B2(HIGHLIGHT), .B1(w2897), .A2(w2781), .A1(w2767) );
	vdp_and g2779 (.nZ(w2837), .B(HIGHLIGHT), .A(w2783) );
	vdp_and g2780 (.nZ(w2838), .B(HIGHLIGHT), .A(w2899) );
	vdp_and g2781 (.nZ(w2835), .B(HIGHLIGHT), .A(w2896) );
	vdp_aon22 g2782 (.nZ(w2839), .B2(w2766), .B1(w2782), .A2(w2783), .A1(w2766) );
	vdp_aon22 g2783 (.nZ(w2895), .B2(w2762), .B1(w2782), .A2(w2785), .A1(HIGHLIGHT) );
	vdp_aon2222 g2784 (.Z(w2784), .B2(w2766), .B1(w2781), .A2(w2899), .A1(w2766), .D2(w2762), .D1(w2781), .C2(w2781), .C1(HIGHLIGHT) );
	vdp_aon22 g2785 (.Z(w2788), .B2(w2762), .B1(w2898), .A2(w2896), .A1(w2767) );
	vdp_aon22 g2786 (.Z(w2789), .B2(w2766), .B1(w2785), .A2(w2896), .A1(w2766) );
	vdp_aon22 g2787 (.Z(w2834), .B2(w2762), .B1(w2785), .A2(w2899), .A1(w2767) );
	vdp_and g2788 (.Z(w2833), .B(w2767), .A(w2785) );
	vdp_and g2789 (.Z(w2832), .B(w2898), .A(w2767) );
	vdp_and g2790 (.Z(w2831), .B(w2767), .A(w2782) );
	vdp_aon22 g2791 (.Z(w2829), .B2(w2762), .B1(w2896), .A2(w2783), .A1(w2767) );
	vdp_aon2222 g2792 (.Z(w2830), .B2(w2766), .B1(w2898), .A2(w2897), .A1(w2766), .D2(w2762), .D1(w2897), .C2(w2897), .C1(w2767) );
	vdp_nor3 g2793 (.Z(w2762), .A(w2766), .B(SHADOW), .C(HIGHLIGHT) );
	vdp_and g2794 (.Z(w2767), .A(SHADOW), .B(w2787) );
	vdp_bufif0 g2795 (.A(w2685), .nE(w2692), .Z(COL[0]) );
	vdp_bufif0 g2796 (.A(w2877), .nE(w2692), .Z(COL[1]) );
	vdp_bufif0 g2797 (.A(w2687), .nE(w2692), .Z(COL[2]) );
	vdp_bufif0 g2798 (.A(w2691), .nE(w2692), .Z(COL[3]) );
	vdp_bufif0 g2799 (.A(w2705), .nE(w2692), .Z(COL[4]) );
	vdp_bufif0 g2800 (.A(w2876), .nE(w2692), .Z(COL[5]) );
	vdp_and g2801 (.Z(w2876), .A(M5), .B(w2703) );
	vdp_or g2802 (.Z(w2705), .A(w2675), .B(w2695) );
	vdp_not g2803 (.nZ(w2569), .A(M5) );
	vdp_not g2804 (.nZ(w2673), .A(w2875) );
	vdp_not g2805 (.nZ(w2674), .A(w2676) );
	vdp_not g2806 (.nZ(w2675), .A(M5) );
	vdp_not g2807 (.nZ(w2671), .A(w2677) );
	vdp_not g2808 (.nZ(w2692), .A(w2680) );
	vdp_comp_strong g2809 (.nZ(w2683), .Z(w2693), .A(w163) );
	vdp_not g2810 (.nZ(w2681), .A(w89) );
	vdp_not g2811 (.nZ(w2888), .A(w18) );
	vdp_aon222 g2812 (.Z(w2872), .B2(w2673), .A2(w2674), .A1(VRAMA[0]), .B1(VRAMA[1]), .C2(w2671), .C1(COL[0]) );
	vdp_aon222 g2813 (.Z(w2889), .B2(w2673), .A2(w2674), .A1(VRAMA[1]), .B1(VRAMA[2]), .C2(w2671), .C1(COL[1]) );
	vdp_aon222 g2814 (.Z(w2686), .B2(w2673), .A2(w2674), .A1(VRAMA[2]), .B1(VRAMA[3]), .C2(w2671), .C1(COL[2]) );
	vdp_aon222 g2815 (.Z(w2696), .B2(w2673), .A2(w2674), .A1(VRAMA[3]), .B1(VRAMA[4]), .C2(w2671), .C1(COL[3]) );
	vdp_aon222 g2816 (.Z(w2702), .B2(w2673), .A2(w2674), .A1(VRAMA[4]), .B1(VRAMA[5]), .C2(w2671), .C1(COL[4]) );
	vdp_aon222 g2817 (.Z(w2761), .B2(w2673), .A2(w2674), .A1(1'b0), .B1(VRAMA[6]), .C2(w2671), .C1(COL[5]) );
	vdp_nand g2818 (.Z(w2875), .A(w2677), .B(M5) );
	vdp_nand g2819 (.Z(w2676), .A(w2677), .B(w2675) );
	vdp_and g2820 (.Z(w2707), .A(w2708), .B(w2923) );
	vdp_aon222 g2821 (.Z(w2923), .B2(w2918), .A2(w2713), .A1(w2668), .B1(w2715), .C2(w2917), .C1(w2736) );
	vdp_not g2822 (.nZ(w2918), .A(w2871) );
	vdp_not g2823 (.nZ(w2917), .A(w2669) );
	vdp_not g2824 (.nZ(w2741), .A(w2726) );
	vdp_nor g2825 (.Z(w2715), .A(w2669), .B(w2864) );
	vdp_nor g2826 (.Z(w2871), .A(w2736), .B(w2735) );
	vdp_and g2827 (.Z(w2714), .A(w2709), .B(w2749) );
	vdp_and g2828 (.Z(w2713), .A(w2726), .B(w2740) );
	vdp_and g2829 (.Z(w2743), .A(w2740), .B(w2741) );
	vdp_or g2830 (.Z(w2864), .A(w2744), .B(w2743) );
	vdp_or g2831 (.Z(w2712), .A(w2668), .B(w2669) );
	vdp_and g2832 (.Z(w2682), .A(w2708), .B(w2681) );
	vdp_and g2833 (.Z(w2853), .A(w2709), .B(w2746) );
	vdp_and g2834 (.Z(w2863), .A(w2710), .B(w2748) );
	vdp_not g2835 (.nZ(w2754), .A(w89) );
	vdp_or g2836 (.Z(w2716), .A(w2747), .B(w2733) );
	vdp_not g2837 (.nZ(w2921), .A(w2710) );
	vdp_not g2838 (.nZ(w2851), .A(w2611) );
	vdp_not g2839 (.nZ(w2738), .A(w2727) );
	vdp_not g2840 (.nZ(w2737), .A(w2728) );
	vdp_not g2841 (.nZ(w2742), .A(w2612) );
	vdp_and g2842 (.Z(w2759), .A(w2710), .B(w2745) );
	vdp_and g2843 (.Z(w2739), .A(w2711), .B(w2751) );
	vdp_not g2844 (.nZ(w2862), .A(w86) );
	vdp_not g2845 (.nZ(w2869), .A(w87) );
	vdp_and g2846 (.Z(w2744), .A(w2869), .B(w86) );
	vdp_and g2847 (.Z(w2747), .A(w2862), .B(w87) );
	vdp_and g2848 (.Z(w2758), .A(w86), .B(w87) );
	vdp_or3 g2849 (.Z(w2677), .A(w96), .B(w172), .C(w173) );
	vdp_and3 g2850 (.Z(w2868), .A(w2711), .B(w2710), .C(w2748) );
	vdp_and3 g2851 (.Z(w2746), .A(w2737), .B(w2727), .C(w2612) );
	vdp_and3 g2852 (.Z(w2745), .A(w2738), .B(w2728), .C(w2742) );
	vdp_and3 g2853 (.Z(w2751), .A(w2737), .B(w2727), .C(w2742) );
	vdp_and3 g2854 (.Z(w2748), .A(w2727), .B(w2728), .C(w2742) );
	vdp_and g2855 (.Z(w2858), .A(M5), .B(S_TE) );
	vdp_or g2856 (.Z(w2709), .A(w2851), .B(w2726) );
	vdp_and3 g2857 (.Z(w2719), .A(w2713), .B(w2669), .C(w2871) );
	vdp_and3 g2858 (.Z(w2867), .A(w2711), .B(w2709), .C(w2746) );
	vdp_and3 g2859 (.Z(w2866), .A(w2711), .B(w2709), .C(w2751) );
	vdp_and3 g2860 (.Z(w2733), .A(w2732), .B(w2682), .C(w2921) );
	vdp_and3 g2861 (.Z(w2726), .A(w2712), .B(w2729), .C(w2858) );
	vdp_and3 g2862 (.Z(w2755), .A(w2710), .B(w2709), .C(w2749) );
	vdp_and3 g2863 (.Z(w2920), .A(w2710), .B(w2709), .C(w2745) );
	vdp_and3 g2864 (.Z(w2752), .A(w2711), .B(w2710), .C(w2709) );
	vdp_and3 g2865 (.Z(w2753), .A(w2682), .B(w2750), .C(w2919) );
	vdp_and g2866 (.Z(w2718), .A(w2852), .B(w2865) );
	vdp_not g2867 (.nZ(w2756), .A(w2682) );
	vdp_not g2868 (.nZ(w2919), .A(w2711) );
	vdp_or g2869 (.Z(w2717), .A(w2758), .B(w2753) );
	vdp_or g2870 (.Z(w2865), .A(w2756), .B(w2752) );
	vdp_not g2871 (.nZ(w2880), .A(M5) );
	vdp_notif0 g2872 (.A(w2913), .nE(w2650), .nZ(w321) );
	vdp_notif0 g2873 (.nZ(RD_DATA[2]), .A(w2912), .nE(w2650) );
	vdp_notif0 g2874 (.nZ(RD_DATA[1]), .A(w2911), .nE(w2650) );
	vdp_notif0 g2875 (.nZ(AD_DATA[7]), .A(w2910), .nE(w2650) );
	vdp_notif0 g2876 (.nZ(AD_DATA[6]), .A(w2909), .nE(w2650) );
	vdp_notif0 g2877 (.nZ(AD_DATA[5]), .A(w2908), .nE(w2650) );
	vdp_notif0 g2878 (.nZ(AD_DATA[3]), .A(w2907), .nE(w2650) );
	vdp_notif0 g2879 (.nZ(AD_DATA[2]), .A(w2906), .nE(w2650) );
	vdp_notif0 g2880 (.nZ(AD_DATA[1]), .A(w2905), .nE(w2650) );
	vdp_notif0 g2881 (.nZ(DB[1]), .A(w2643), .nE(w2634) );
	vdp_notif0 g2882 (.nZ(DB[0]), .A(w2642), .nE(w2634) );
	vdp_notif0 g2883 (.nZ(DB[2]), .A(w2854), .nE(w2634) );
	vdp_notif0 g2884 (.nZ(DB[5]), .A(w2825), .nE(w2634) );
	vdp_notif0 g2885 (.nZ(DB[8]), .A(w2641), .nE(w2634) );
	vdp_notif0 g2886 (.nZ(DB[10]), .A(w2821), .nE(w2634) );
	vdp_notif0 g2887 (.nZ(DB[9]), .A(w2666), .nE(w2634) );
	vdp_notif0 g2888 (.nZ(DB[7]), .A(w2667), .nE(w2634) );
	vdp_notif0 g2889 (.nZ(DB[6]), .A(w2631), .nE(w2634) );
	vdp_notif0 g2890 (.nZ(DB[4]), .A(w2629), .nE(w2634) );
	vdp_comp_we g2891 (.A(M5), .nZ(w2624), .Z(w2623) );
	vdp_notif0 g2892 (.nZ(DB[3]), .A(w2856), .nE(w2634) );
	vdp_not g2893 (.A(w76), .nZ(w2634) );
	vdp_and g2894 (.Z(w2625), .A(w2626), .B(w2621) );
	vdp_and3 g2895 (.Z(w2856), .A(w85), .B(w2626), .C(w2855) );
	vdp_and3 g2896 (.Z(w2629), .A(w85), .B(w2626), .C(w2891) );
	vdp_and3 g2897 (.Z(w2631), .A(w85), .B(w2626), .C(w2630) );
	vdp_and3 g2898 (.Z(w2667), .A(w85), .B(w2626), .C(w2633) );
	vdp_and3 g2899 (.Z(w2666), .A(w85), .B(w2626), .C(w2636) );
	vdp_and3 g2900 (.Z(w2821), .A(w85), .B(w2626), .C(w2639) );
	vdp_and3 g2901 (.Z(w2641), .A(M5), .B(w2626), .C(w2640) );
	vdp_and3 g2902 (.Z(w2825), .A(M5), .B(w2626), .C(w2647) );
	vdp_and3 g2903 (.Z(w2854), .A(M5), .B(w2626), .C(w2632) );
	vdp_comp_strong g2904 (.nZ(w2645), .A(w2644), .Z(w2648) );
	vdp_and g2905 (.Z(w2644), .A(w2646), .B(HCLK1) );
	vdp_not g2906 (.nZ(w2650), .A(w2914) );
	vdp_aon22 g2907 (.Z(w2879), .B2(FIFOo[5]), .A2(FIFOo[7]), .A1(w2698), .B1(w2697) );
	vdp_aon22 g2908 (.Z(w2661), .B2(FIFOo[4]), .A2(FIFOo[6]), .A1(w2698), .B1(w2697) );
	vdp_aon22 g2909 (.Z(w2658), .B2(FIFOo[3]), .A2(FIFOo[5]), .A1(w2698), .B1(w2697) );
	vdp_aon22 g2910 (.Z(w2657), .B2(FIFOo[2]), .A2(FIFOo[3]), .A1(w2698), .B1(w2697) );
	vdp_aon22 g2911 (.Z(w2656), .B2(FIFOo[1]), .A2(FIFOo[2]), .A1(w2698), .B1(w2697) );
	vdp_aon22 g2912 (.Z(w2660), .B2(FIFOo[0]), .A2(FIFOo[1]), .A1(w2698), .B1(w2697) );
	vdp_comp_we g2913 (.Z(w2698), .nZ(w2697), .A(M5) );
	vdp_aon22 g2914 (.Z(w2689), .B2(w2880), .A2(M5), .A1(w2857), .B1(w17) );
	vdp_aon22 g2915 (.Z(COL[7]), .B2(w2720), .A2(w2706), .A1(w89), .B1(w2754) );
	vdp_aon22 g2916 (.Z(w117), .B2(w2734), .A2(w2850), .A1(w89), .B1(w2754) );
	vdp_and3 g2917 (.Z(w2740), .A(w2682), .B(w2611), .C(w2922) );
	vdp_aon22 g2918 (.Z(w2749), .B2(w2737), .A2(w2728), .A1(w2612), .B1(w2738) );
	vdp_aon22 g2919 (.Z(w2633), .B2(w2647), .A2(w2637), .A1(w2623), .B1(w2624) );
	vdp_aon22 g2920 (.Z(w2630), .B2(w2627), .A2(w2628), .A1(w2623), .B1(w2624) );
	vdp_aon22 g2921 (.Z(w2855), .B2(w2632), .A2(w2622), .A1(w2623), .B1(w2624) );
	vdp_aon22 g2922 (.Z(w2891), .B2(w2622), .A2(w2627), .A1(w2623), .B1(w2624) );
	vdp_aon22 g2923 (.Z(w2636), .B2(w2628), .A2(w2635), .A1(w2623), .B1(w2624) );
	vdp_aon22 g2924 (.Z(w2639), .B2(w2637), .A2(w2638), .A1(w2623), .B1(w2624) );
	vdp_and4 g2925 (.Z(w2735), .A(w2738), .B(w2612), .C(w2858), .D(w2737) );
	vdp_or5 g2926 (.Z(w2732), .A(w2714), .B(w2745), .C(w2748), .D(w2867), .E(w2866) );
	vdp_or5 g2927 (.Z(w2750), .A(w2755), .B(w2751), .C(w2853), .D(w2863), .E(w2920) );
	vdp_or5 g2928 (.Z(w2922), .A(w2746), .B(w2749), .C(w2759), .D(w2739), .E(w2868) );
	vdp_nor4 g2929 (.Z(w2699), .A(COL[2]), .B(COL[3]), .C(COL[1]), .D(COL[0]) );
	vdp_nor g2930 (.Z(w2852), .A(w86), .B(w87) );
	vdp_nor g2931 (.Z(w2710), .A(w2870), .B(w2874) );
	vdp_nor g2932 (.Z(w2870), .A(w2611), .B(M5) );
	vdp_nand g2933 (.Z(w2711), .A(M5), .B(w2873) );
	vdp_nand g2934 (.Z(w2722), .A(SPR_PRIO), .B(w18) );
	vdp_and4 g2935 (.Z(w2736), .A(w2737), .B(w2858), .C(w2738), .D(w2742) );
	vdp_aoi21 g2936 (.Z(w2890), .B(w2625), .A2(w2888), .A1(w2672) );
	vdp_nor g2937 (.Z(w2760), .A(w20), .B(w19) );
	vdp_n_fet g2938 (.A(w2680), .Z(COL[6]) );
	vdp_slatch g2939 (.Q(w3999), .D(S[3]), .C(w3050), .nC(w3040) );
	vdp_slatch g2940 (.Q(w4001), .D(S[3]), .C(w3031), .nC(w3030) );
	vdp_slatch g2941 (.Q(w4003), .D(S[3]), .C(w3032), .nC(w3028) );
	vdp_slatch g2942 (.Q(w4005), .D(S[3]), .C(w3049), .nC(w3041) );
	vdp_slatch g2943 (.Q(w4007), .D(S[7]), .C(w3050), .nC(w3040) );
	vdp_slatch g2944 (.Q(w4010), .D(S[7]), .C(w3031), .nC(w3030) );
	vdp_slatch g2945 (.Q(w4009), .D(S[7]), .C(w3032), .nC(w3028) );
	vdp_slatch g2946 (.Q(w4014), .D(S[7]), .C(w3049), .nC(w3041) );
	vdp_slatch g2947 (.Q(w4013), .D(S[2]), .C(w3050), .nC(w3040) );
	vdp_slatch g2948 (.Q(w4020), .D(S[2]), .C(w3031), .nC(w3030) );
	vdp_slatch g2949 (.Q(w4019), .D(S[2]), .C(w3032), .nC(w3028) );
	vdp_slatch g2950 (.Q(w4022), .D(S[2]), .C(w3049), .nC(w3041) );
	vdp_slatch g2951 (.Q(w4021), .D(S[6]), .C(w3050), .nC(w3040) );
	vdp_slatch g2952 (.Q(w4026), .D(S[6]), .C(w3031), .nC(w3030) );
	vdp_slatch g2953 (.Q(w4025), .D(S[6]), .C(w3032), .nC(w3028) );
	vdp_slatch g2954 (.Q(w4030), .D(S[6]), .C(w3049), .nC(w3041) );
	vdp_slatch g2955 (.Q(w4029), .D(S[1]), .C(w3050), .nC(w3040) );
	vdp_slatch g2956 (.Q(w4034), .D(S[1]), .C(w3031), .nC(w3030) );
	vdp_slatch g2957 (.Q(w4033), .D(S[1]), .C(w3032), .nC(w3028) );
	vdp_slatch g2958 (.Q(w4038), .D(S[1]), .C(w3049), .nC(w3041) );
	vdp_slatch g2959 (.Q(w4037), .D(S[5]), .C(w3050), .nC(w3040) );
	vdp_slatch g2960 (.Q(w4042), .D(S[5]), .C(w3031), .nC(w3030) );
	vdp_slatch g2961 (.Q(w4041), .D(S[5]), .C(w3032), .nC(w3028) );
	vdp_slatch g2962 (.Q(w4046), .D(S[5]), .C(w3049), .nC(w3041) );
	vdp_slatch g2963 (.Q(w4045), .D(S[0]), .C(w3050), .nC(w3040) );
	vdp_slatch g2964 (.Q(w4050), .D(S[0]), .C(w3031), .nC(w3030) );
	vdp_slatch g2965 (.Q(w4049), .D(S[0]), .C(w3032), .nC(w3028) );
	vdp_slatch g2966 (.Q(w4054), .D(S[0]), .C(w3049), .nC(w3041) );
	vdp_slatch g2967 (.Q(w4053), .D(S[4]), .C(w3050), .nC(w3040) );
	vdp_slatch g2968 (.Q(w4058), .D(S[4]), .C(w3031), .nC(w3030) );
	vdp_slatch g2969 (.Q(w4057), .D(S[4]), .C(w3032), .nC(w3028) );
	vdp_slatch g2970 (.Q(w4061), .D(S[4]), .C(w3049), .nC(w3041) );
	vdp_slatch g2971 (.Q(w4000), .D(w3999), .C(w3019), .nC(w3037) );
	vdp_slatch g2972 (.Q(w4002), .D(w4001), .C(w3038), .nC(w3029) );
	vdp_slatch g2973 (.Q(w4004), .D(w4003), .C(w3039), .nC(w3027) );
	vdp_slatch g2974 (.Q(w4006), .D(w4005), .C(w3035), .nC(w3036) );
	vdp_slatch g2975 (.Q(w4008), .D(w4007), .C(w3019), .nC(w3037) );
	vdp_slatch g2976 (.Q(w4012), .D(w4010), .C(w3038), .nC(w3029) );
	vdp_slatch g2977 (.Q(w4011), .D(w4009), .C(w3039), .nC(w3027) );
	vdp_slatch g2978 (.Q(w4016), .D(w4014), .C(w3035), .nC(w3036) );
	vdp_slatch g2979 (.Q(w4015), .D(w4013), .C(w3019), .nC(w3037) );
	vdp_slatch g2980 (.Q(w4018), .D(w4020), .C(w3038), .nC(w3029) );
	vdp_slatch g2981 (.Q(w4017), .D(w4019), .C(w3039), .nC(w3027) );
	vdp_slatch g2982 (.Q(w4024), .D(w4022), .C(w3035), .nC(w3036) );
	vdp_slatch g2983 (.Q(w4023), .D(w4021), .C(w3019), .nC(w3037) );
	vdp_slatch g2984 (.Q(w4028), .D(w4026), .C(w3038), .nC(w3029) );
	vdp_slatch g2985 (.Q(w4027), .D(w4025), .C(w3039), .nC(w3027) );
	vdp_slatch g2986 (.Q(w4032), .D(w4030), .C(w3035), .nC(w3036) );
	vdp_slatch g2987 (.Q(w4031), .D(w4029), .C(w3019), .nC(w3037) );
	vdp_slatch g2988 (.Q(w4036), .D(w4034), .C(w3038), .nC(w3029) );
	vdp_slatch g2989 (.Q(w4035), .D(w4033), .C(w3039), .nC(w3027) );
	vdp_slatch g2990 (.Q(w4040), .D(w4038), .C(w3035), .nC(w3036) );
	vdp_slatch g2991 (.Q(w4039), .D(w4037), .C(w3019), .nC(w3037) );
	vdp_slatch g2992 (.Q(w4044), .D(w4042), .C(w3038), .nC(w3029) );
	vdp_slatch g2993 (.Q(w4043), .D(w4041), .C(w3039), .nC(w3027) );
	vdp_slatch g2994 (.Q(w4048), .D(w4046), .C(w3035), .nC(w3036) );
	vdp_slatch g2995 (.Q(w4047), .D(w4045), .C(w3019), .nC(w3037) );
	vdp_slatch g2996 (.Q(w4052), .D(w4050), .C(w3038), .nC(w3029) );
	vdp_slatch g2997 (.Q(w4051), .D(w4049), .C(w3039), .nC(w3027) );
	vdp_slatch g2998 (.Q(w4056), .D(w4054), .C(w3035), .nC(w3036) );
	vdp_slatch g2999 (.Q(w4055), .D(w4053), .C(w3019), .nC(w3037) );
	vdp_slatch g3000 (.Q(w4060), .D(w4058), .C(w3038), .nC(w3029) );
	vdp_slatch g3001 (.Q(w4059), .D(w4057), .C(w3039), .nC(w3027) );
	vdp_slatch g3002 (.Q(w4062), .D(w4061), .C(w3035), .nC(w3036) );
	vdp_slatch g3003 (.Q(w3077), .D(w4000), .C(w3042), .nC(w3068) );
	vdp_slatch g3004 (.Q(w3076), .D(w4002), .C(w3020), .nC(w3078) );
	vdp_slatch g3005 (.Q(w3075), .D(w4004), .C(w3033), .nC(w3079) );
	vdp_slatch g3006 (.Q(w3074), .D(w4006), .C(w3034), .nC(w3007) );
	vdp_slatch g3007 (.Q(w3073), .D(w4008), .C(w3042), .nC(w3068) );
	vdp_slatch g3008 (.Q(w3072), .D(w4012), .C(w3020), .nC(w3078) );
	vdp_slatch g3009 (.Q(w3071), .D(w4011), .C(w3033), .nC(w3079) );
	vdp_slatch g3010 (.Q(w3070), .D(w4016), .C(w3034), .nC(w3007) );
	vdp_slatch g3011 (.Q(w3069), .D(w4015), .C(w3042), .nC(w3068) );
	vdp_slatch g3012 (.Q(w3082), .D(w4018), .C(w3020), .nC(w3078) );
	vdp_slatch g3013 (.Q(w3086), .D(w4017), .C(w3033), .nC(w3079) );
	vdp_slatch g3014 (.Q(w3085), .D(w4024), .C(w3034), .nC(w3007) );
	vdp_slatch g3015 (.Q(w3084), .D(w4023), .C(w3042), .nC(w3068) );
	vdp_slatch g3016 (.Q(w3080), .D(w4028), .C(w3020), .nC(w3078) );
	vdp_slatch g3017 (.Q(w3081), .D(w4027), .C(w3033), .nC(w3079) );
	vdp_slatch g3018 (.D(w4032), .Q(w3083), .C(w3034), .nC(w3007) );
	vdp_slatch g3019 (.Q(w3087), .D(w4031), .C(w3042), .nC(w3068) );
	vdp_slatch g3020 (.Q(w3088), .D(w4036), .C(w3020), .nC(w3078) );
	vdp_slatch g3021 (.Q(w3090), .D(w4035), .C(w3033), .nC(w3079) );
	vdp_slatch g3022 (.Q(w3089), .D(w4040), .C(w3034), .nC(w3007) );
	vdp_slatch g3023 (.Q(w3131), .D(w4039), .C(w3042), .nC(w3068) );
	vdp_slatch g3024 (.Q(w3132), .D(w4044), .C(w3020), .nC(w3078) );
	vdp_slatch g3025 (.Q(w3128), .D(w4043), .C(w3033), .nC(w3079) );
	vdp_slatch g3026 (.Q(w3123), .D(w4048), .C(w3034), .nC(w3007) );
	vdp_slatch g3027 (.Q(w3135), .D(w4047), .C(w3042), .nC(w3068) );
	vdp_slatch g3028 (.Q(w3134), .D(w4052), .C(w3020), .nC(w3078) );
	vdp_slatch g3029 (.Q(w3133), .D(w4051), .C(w3033), .nC(w3079) );
	vdp_slatch g3030 (.Q(w3130), .D(w4056), .C(w3034), .nC(w3007) );
	vdp_slatch g3031 (.Q(w3116), .D(w4055), .C(w3042), .nC(w3068) );
	vdp_slatch g3032 (.Q(w3115), .D(w4060), .C(w3020), .nC(w3078) );
	vdp_slatch g3033 (.Q(w3117), .D(w4059), .C(w3033), .nC(w3079) );
	vdp_slatch g3034 (.Q(w3118), .D(w4062), .C(w3034), .nC(w3007) );
	vdp_slatch g3035 (.Q(w3195), .D(w4283), .C(w3191), .nC(w3193) );
	vdp_slatch g3036 (.Q(w3196), .D(w4284), .C(w3190), .nC(w3201) );
	vdp_slatch g3037 (.Q(w3197), .D(w4286), .C(w3189), .nC(w3202) );
	vdp_slatch g3038 (.Q(w3198), .D(w4285), .C(w3188), .nC(w3194) );
	vdp_slatch g3039 (.Q(w3199), .D(w4118), .C(w3191), .nC(w3193) );
	vdp_slatch g3040 (.Q(w3200), .D(w4117), .C(w3190), .nC(w3201) );
	vdp_slatch g3041 (.Q(w3206), .D(w4112), .C(w3189), .nC(w3202) );
	vdp_slatch g3042 (.Q(w3207), .D(w4111), .C(w3188), .nC(w3194) );
	vdp_slatch g3043 (.Q(w3208), .D(w4108), .C(w3191), .nC(w3193) );
	vdp_slatch g3044 (.Q(w3209), .D(w4107), .C(w3190), .nC(w3201) );
	vdp_slatch g3045 (.Q(w3210), .D(w4106), .C(w3189), .nC(w3202) );
	vdp_slatch g3046 (.Q(w3205), .D(w4103), .C(w3188), .nC(w3194) );
	vdp_slatch g3047 (.Q(w3211), .D(w4100), .C(w3191), .nC(w3193) );
	vdp_slatch g3048 (.Q(w3212), .D(w4101), .C(w3190), .nC(w3201) );
	vdp_slatch g3049 (.Q(w3213), .D(w4096), .C(w3189), .nC(w3202) );
	vdp_slatch g3050 (.Q(w3214), .D(w4097), .C(w3188), .nC(w3194) );
	vdp_slatch g3051 (.Q(w3139), .D(w4094), .C(w3191), .nC(w3193) );
	vdp_slatch g3052 (.Q(w3891), .D(w4093), .C(w3190), .nC(w3201) );
	vdp_slatch g3053 (.Q(w3141), .D(w4090), .C(w3189), .nC(w3202) );
	vdp_slatch g3054 (.Q(w3142), .D(w4089), .C(w3188), .nC(w3194) );
	vdp_slatch g3055 (.Q(w3215), .D(w4086), .C(w3191), .nC(w3193) );
	vdp_slatch g3056 (.Q(w3140), .D(w4085), .C(w3190), .nC(w3201) );
	vdp_slatch g3057 (.Q(w3120), .D(w4082), .C(w3189), .nC(w3202) );
	vdp_slatch g3058 (.Q(w3143), .D(w4081), .C(w3188), .nC(w3194) );
	vdp_slatch g3059 (.Q(w3146), .D(w4078), .C(w3191), .nC(w3193) );
	vdp_slatch g3060 (.Q(w3154), .D(w4077), .C(w3190), .nC(w3201) );
	vdp_slatch g3061 (.Q(w3153), .D(w4074), .C(w3189), .nC(w3202) );
	vdp_slatch g3062 (.Q(w3152), .D(w4073), .C(w3188), .nC(w3194) );
	vdp_slatch g3063 (.Q(w3150), .D(w4070), .C(w3191), .nC(w3193) );
	vdp_slatch g3064 (.Q(w3144), .D(w4069), .C(w3190), .nC(w3201) );
	vdp_slatch g3065 (.Q(w3151), .D(w4066), .C(w3189), .nC(w3202) );
	vdp_slatch g3066 (.Q(w3145), .D(w4065), .C(w3188), .nC(w3194) );
	vdp_slatch g3067 (.Q(w4283), .D(w4121), .C(w3192), .nC(w3179) );
	vdp_slatch g3068 (.Q(w4284), .D(w4122), .C(w2999), .nC(w3180) );
	vdp_slatch g3069 (.Q(w4286), .D(w4120), .C(w3186), .nC(w2987) );
	vdp_slatch g3070 (.Q(w4285), .D(w4119), .C(w3187), .nC(w2988) );
	vdp_slatch g3071 (.Q(w4118), .D(w4116), .C(w3192), .nC(w3179) );
	vdp_slatch g3072 (.Q(w4117), .D(w4115), .C(w2999), .nC(w3180) );
	vdp_slatch g3073 (.Q(w4112), .D(w4114), .C(w3186), .nC(w2987) );
	vdp_slatch g3074 (.Q(w4111), .D(w4113), .C(w3187), .nC(w2988) );
	vdp_slatch g3075 (.Q(w4108), .D(w4110), .C(w3192), .nC(w3179) );
	vdp_slatch g3076 (.Q(w4107), .D(w4109), .C(w2999), .nC(w3180) );
	vdp_slatch g3077 (.Q(w4106), .D(w4104), .C(w3186), .nC(w2987) );
	vdp_slatch g3078 (.Q(w4103), .D(w4105), .C(w3187), .nC(w2988) );
	vdp_slatch g3079 (.Q(w4100), .D(w4102), .C(w3192), .nC(w3179) );
	vdp_slatch g3080 (.Q(w4101), .D(w4099), .C(w2999), .nC(w3180) );
	vdp_slatch g3081 (.Q(w4096), .D(w4098), .C(w3186), .nC(w2987) );
	vdp_slatch g3082 (.Q(w4097), .D(w4095), .C(w3187), .nC(w2988) );
	vdp_slatch g3083 (.Q(w4094), .D(w4092), .C(w3192), .nC(w3179) );
	vdp_slatch g3084 (.Q(w4093), .D(w4091), .C(w2999), .nC(w3180) );
	vdp_slatch g3085 (.Q(w4090), .D(w4088), .C(w3186), .nC(w2987) );
	vdp_slatch g3086 (.Q(w4089), .D(w4087), .C(w3187), .nC(w2988) );
	vdp_slatch g3087 (.Q(w4086), .D(w4084), .C(w3192), .nC(w3179) );
	vdp_slatch g3088 (.Q(w4085), .D(w4083), .C(w2999), .nC(w3180) );
	vdp_slatch g3089 (.Q(w4082), .D(w4080), .C(w3186), .nC(w2987) );
	vdp_slatch g3090 (.Q(w4081), .D(w4079), .C(w3187), .nC(w2988) );
	vdp_slatch g3091 (.Q(w4078), .D(w4076), .C(w3192), .nC(w3179) );
	vdp_slatch g3092 (.Q(w4077), .D(w4075), .C(w2999), .nC(w3180) );
	vdp_slatch g3093 (.Q(w4074), .D(w4072), .C(w3186), .nC(w2987) );
	vdp_slatch g3094 (.Q(w4073), .D(w4071), .C(w3187), .nC(w2988) );
	vdp_slatch g3095 (.Q(w4070), .D(w4068), .C(w3192), .nC(w3179) );
	vdp_slatch g3096 (.Q(w4069), .D(w4067), .C(w2999), .nC(w3180) );
	vdp_slatch g3097 (.Q(w4066), .D(w4064), .C(w3186), .nC(w2987) );
	vdp_slatch g3098 (.Q(w4065), .D(w4063), .C(w3187), .nC(w2988) );
	vdp_slatch g3099 (.Q(w4121), .D(S[3]), .C(w2952), .nC(w2985) );
	vdp_slatch g3100 (.Q(w4122), .D(S[3]), .C(w2956), .nC(w2989) );
	vdp_slatch g3101 (.Q(w4120), .D(S[3]), .C(w2959), .nC(w2986) );
	vdp_slatch g3102 (.Q(w4119), .D(S[3]), .C(w2961), .nC(w2984) );
	vdp_slatch g3103 (.Q(w4116), .D(S[7]), .C(w2952), .nC(w2985) );
	vdp_slatch g3104 (.Q(w4115), .D(S[7]), .C(w2956), .nC(w2989) );
	vdp_slatch g3105 (.Q(w4114), .D(S[7]), .C(w2959), .nC(w2986) );
	vdp_slatch g3106 (.Q(w4113), .D(S[7]), .C(w2961), .nC(w2984) );
	vdp_slatch g3107 (.Q(w4110), .D(S[2]), .C(w2952), .nC(w2985) );
	vdp_slatch g3108 (.Q(w4109), .D(S[2]), .C(w2956), .nC(w2989) );
	vdp_slatch g3109 (.Q(w4104), .D(S[2]), .C(w2959), .nC(w2986) );
	vdp_slatch g3110 (.Q(w4105), .D(S[2]), .C(w2961), .nC(w2984) );
	vdp_slatch g3111 (.Q(w4102), .D(S[6]), .C(w2952), .nC(w2985) );
	vdp_slatch g3112 (.Q(w4099), .D(S[6]), .C(w2956), .nC(w2989) );
	vdp_slatch g3113 (.Q(w4098), .D(S[6]), .C(w2959), .nC(w2986) );
	vdp_slatch g3114 (.Q(w4095), .D(S[6]), .C(w2961), .nC(w2984) );
	vdp_slatch g3115 (.Q(w4092), .D(S[1]), .C(w2952), .nC(w2985) );
	vdp_slatch g3116 (.Q(w4091), .D(S[1]), .C(w2956), .nC(w2989) );
	vdp_slatch g3117 (.Q(w4088), .D(S[1]), .C(w2959), .nC(w2986) );
	vdp_slatch g3118 (.Q(w4087), .D(S[1]), .C(w2961), .nC(w2984) );
	vdp_slatch g3119 (.Q(w4084), .D(S[5]), .C(w2952), .nC(w2985) );
	vdp_slatch g3120 (.Q(w4083), .D(S[5]), .C(w2956), .nC(w2989) );
	vdp_slatch g3121 (.Q(w4080), .D(S[5]), .C(w2959), .nC(w2986) );
	vdp_slatch g3122 (.Q(w4079), .D(S[5]), .C(w2961), .nC(w2984) );
	vdp_slatch g3123 (.Q(w4076), .D(S[0]), .C(w2952), .nC(w2985) );
	vdp_slatch g3124 (.Q(w4075), .D(S[0]), .C(w2956), .nC(w2989) );
	vdp_slatch g3125 (.Q(w4072), .D(S[0]), .C(w2959), .nC(w2986) );
	vdp_slatch g3126 (.Q(w4071), .D(S[0]), .C(w2961), .nC(w2984) );
	vdp_slatch g3127 (.Q(w4068), .D(S[4]), .C(w2952), .nC(w2985) );
	vdp_slatch g3128 (.Q(w4067), .D(S[4]), .C(w2956), .nC(w2989) );
	vdp_slatch g3129 (.Q(w4064), .D(S[4]), .C(w2959), .nC(w2986) );
	vdp_slatch g3130 (.Q(w4063), .D(S[4]), .C(w2961), .nC(w2984) );
	vdp_slatch g3131 (.Q(w4126), .D(S[3]), .C(w2953), .nC(w2977) );
	vdp_slatch g3132 (.Q(w4125), .D(S[3]), .C(w2957), .nC(w2982) );
	vdp_slatch g3133 (.Q(w4130), .D(S[3]), .C(w2958), .nC(w2983) );
	vdp_slatch g3134 (.Q(w4129), .D(S[3]), .C(w2960), .nC(w2978) );
	vdp_slatch g3135 (.Q(w4134), .D(S[7]), .C(w2953), .nC(w2977) );
	vdp_slatch g3136 (.Q(w4133), .D(S[7]), .C(w2957), .nC(w2982) );
	vdp_slatch g3137 (.Q(w4138), .D(S[7]), .C(w2958), .nC(w2983) );
	vdp_slatch g3138 (.Q(w4137), .D(S[7]), .C(w2960), .nC(w2978) );
	vdp_slatch g3139 (.Q(w4142), .D(S[2]), .C(w2953), .nC(w2977) );
	vdp_slatch g3140 (.Q(w4141), .D(S[2]), .C(w2957), .nC(w2982) );
	vdp_slatch g3141 (.Q(w4146), .D(S[2]), .C(w2958), .nC(w2983) );
	vdp_slatch g3142 (.Q(w4145), .D(S[2]), .C(w2960), .nC(w2978) );
	vdp_slatch g3143 (.Q(w4148), .D(S[6]), .C(w2953), .nC(w2977) );
	vdp_slatch g3144 (.Q(w4149), .D(S[6]), .C(w2957), .nC(w2982) );
	vdp_slatch g3145 (.Q(w4185), .D(S[6]), .C(w2958), .nC(w2983) );
	vdp_slatch g3146 (.Q(w4184), .D(S[6]), .C(w2960), .nC(w2978) );
	vdp_slatch g3147 (.Q(w4181), .D(S[1]), .C(w2953), .nC(w2977) );
	vdp_slatch g3148 (.Q(w4180), .D(S[1]), .C(w2957), .nC(w2982) );
	vdp_slatch g3149 (.Q(w4177), .D(S[1]), .C(w2958), .nC(w2983) );
	vdp_slatch g3150 (.Q(w4176), .D(S[1]), .C(w2960), .nC(w2978) );
	vdp_slatch g3151 (.Q(w4173), .D(S[5]), .C(w2953), .nC(w2977) );
	vdp_slatch g3152 (.Q(w4172), .D(S[5]), .C(w2957), .nC(w2982) );
	vdp_slatch g3153 (.Q(w4169), .D(S[5]), .C(w2958), .nC(w2983) );
	vdp_slatch g3154 (.Q(w4168), .D(S[5]), .C(w2960), .nC(w2978) );
	vdp_slatch g3155 (.Q(w4165), .D(S[0]), .C(w2953), .nC(w2977) );
	vdp_slatch g3156 (.Q(w4164), .D(S[0]), .C(w2957), .nC(w2982) );
	vdp_slatch g3157 (.Q(w4161), .D(S[0]), .C(w2958), .nC(w2983) );
	vdp_slatch g3158 (.Q(w4160), .D(S[0]), .C(w2960), .nC(w2978) );
	vdp_slatch g3159 (.Q(w4157), .D(S[4]), .C(w2953), .nC(w2977) );
	vdp_slatch g3160 (.Q(w4156), .D(S[4]), .C(w2957), .nC(w2982) );
	vdp_slatch g3161 (.Q(w4153), .D(S[4]), .C(w2958), .nC(w2983) );
	vdp_slatch g3162 (.Q(w4152), .D(S[4]), .C(w2960), .nC(w2978) );
	vdp_slatch g3163 (.Q(w4124), .D(w4126), .C(w2940), .nC(w2979) );
	vdp_slatch g3164 (.Q(w4123), .D(w4125), .C(w2943), .nC(w2980) );
	vdp_slatch g3165 (.Q(w4128), .D(w4130), .C(w2948), .nC(w2981) );
	vdp_slatch g3166 (.Q(w4127), .D(w4129), .C(w2945), .nC(w2950) );
	vdp_slatch g3167 (.Q(w4132), .D(w4134), .C(w2940), .nC(w2979) );
	vdp_slatch g3168 (.Q(w4131), .D(w4133), .C(w2943), .nC(w2980) );
	vdp_slatch g3169 (.Q(w4136), .D(w4138), .C(w2948), .nC(w2981) );
	vdp_slatch g3170 (.Q(w4135), .D(w4137), .C(w2945), .nC(w2950) );
	vdp_slatch g3171 (.Q(w4140), .D(w4142), .C(w2940), .nC(w2979) );
	vdp_slatch g3172 (.Q(w4139), .D(w4141), .C(w2943), .nC(w2980) );
	vdp_slatch g3173 (.Q(w4250), .D(w4146), .C(w2948), .nC(w2981) );
	vdp_slatch g3174 (.Q(w4144), .D(w4145), .C(w2945), .nC(w2950) );
	vdp_slatch g3175 (.Q(w4143), .D(w4148), .C(w2940), .nC(w2979) );
	vdp_slatch g3176 (.Q(w4147), .D(w4149), .C(w2943), .nC(w2980) );
	vdp_slatch g3177 (.Q(w4183), .D(w4185), .C(w2948), .nC(w2981) );
	vdp_slatch g3178 (.Q(w4182), .D(w4184), .C(w2945), .nC(w2950) );
	vdp_slatch g3179 (.Q(w4179), .D(w4181), .C(w2940), .nC(w2979) );
	vdp_slatch g3180 (.Q(w4178), .D(w4180), .C(w2943), .nC(w2980) );
	vdp_slatch g3181 (.Q(w4175), .D(w4177), .C(w2948), .nC(w2981) );
	vdp_slatch g3182 (.Q(w4174), .D(w4176), .C(w2945), .nC(w2950) );
	vdp_slatch g3183 (.Q(w4171), .D(w4173), .C(w2940), .nC(w2979) );
	vdp_slatch g3184 (.Q(w4170), .D(w4172), .C(w2943), .nC(w2980) );
	vdp_slatch g3185 (.Q(w4167), .D(w4169), .C(w2948), .nC(w2981) );
	vdp_slatch g3186 (.Q(w4166), .D(w4168), .C(w2945), .nC(w2950) );
	vdp_slatch g3187 (.D(w4165), .Q(w4163), .C(w2940), .nC(w2979) );
	vdp_slatch g3188 (.Q(w4162), .D(w4164), .C(w2943), .nC(w2980) );
	vdp_slatch g3189 (.Q(w4159), .D(w4161), .C(w2948), .nC(w2981) );
	vdp_slatch g3190 (.Q(w4158), .D(w4160), .C(w2945), .nC(w2950) );
	vdp_slatch g3191 (.Q(w4155), .D(w4157), .C(w2940), .nC(w2979) );
	vdp_slatch g3192 (.Q(w4154), .D(w4156), .C(w2943), .nC(w2980) );
	vdp_slatch g3193 (.Q(w4151), .D(w4153), .C(w2948), .nC(w2981) );
	vdp_slatch g3194 (.Q(w4150), .D(w4152), .C(w2945), .nC(w2950) );
	vdp_slatch g3195 (.Q(w3261), .D(w4124), .C(w2941), .nC(w2942) );
	vdp_slatch g3196 (.Q(w3260), .D(w4123), .C(w2949), .nC(w2944) );
	vdp_slatch g3197 (.Q(w3248), .D(w4128), .C(w2946), .nC(w2947) );
	vdp_slatch g3198 (.Q(w3246), .D(w4127), .C(w2939), .nC(w2938) );
	vdp_slatch g3199 (.Q(w3259), .D(w4132), .C(w2941), .nC(w2942) );
	vdp_slatch g3200 (.Q(w3258), .D(w4131), .C(w2949), .nC(w2944) );
	vdp_slatch g3201 (.D(w4136), .C(w2946), .nC(w2947), .Q(w3257) );
	vdp_slatch g3202 (.Q(w3245), .D(w4135), .C(w2939), .nC(w2938) );
	vdp_slatch g3203 (.Q(w3256), .D(w4140), .C(w2941), .nC(w2942) );
	vdp_slatch g3204 (.Q(w3255), .D(w4139), .C(w2949), .nC(w2944) );
	vdp_slatch g3205 (.Q(w3254), .D(w4250), .C(w2946), .nC(w2947) );
	vdp_slatch g3206 (.Q(w3253), .D(w4144), .C(w2939), .nC(w2938) );
	vdp_slatch g3207 (.Q(w3252), .D(w4143), .C(w2941), .nC(w2942) );
	vdp_slatch g3208 (.Q(w3251), .D(w4147), .C(w2949), .nC(w2944) );
	vdp_slatch g3209 (.Q(w3250), .D(w4183), .C(w2946), .nC(w2947) );
	vdp_slatch g3210 (.Q(w3249), .D(w4182), .C(w2939), .nC(w2938) );
	vdp_slatch g3211 (.Q(w3241), .D(w4179), .C(w2941), .nC(w2942) );
	vdp_slatch g3212 (.Q(w3287), .D(w4178), .C(w2949), .nC(w2944) );
	vdp_slatch g3213 (.Q(w3242), .D(w4175), .C(w2946), .nC(w2947) );
	vdp_slatch g3214 (.Q(w3243), .D(w4174), .C(w2939), .nC(w2938) );
	vdp_slatch g3215 (.Q(w3291), .D(w4171), .C(w2941), .nC(w2942) );
	vdp_slatch g3216 (.Q(w3300), .D(w4170), .C(w2949), .nC(w2944) );
	vdp_slatch g3217 (.Q(w3292), .D(w4167), .C(w2946), .nC(w2947) );
	vdp_slatch g3218 (.Q(w3299), .D(w4166), .nC(w2938), .C(w2939) );
	vdp_slatch g3219 (.Q(w3298), .D(w4163), .C(w2941), .nC(w2942) );
	vdp_slatch g3220 (.Q(w3297), .D(w4162), .C(w2949), .nC(w2944) );
	vdp_slatch g3221 (.Q(w3293), .D(w4159), .C(w2946), .nC(w2947) );
	vdp_slatch g3222 (.Q(w3296), .D(w4158), .C(w2939), .nC(w2938) );
	vdp_slatch g3223 (.Q(w3295), .D(w4155), .C(w2941), .nC(w2942) );
	vdp_slatch g3224 (.Q(w3294), .D(w4154), .C(w2949), .nC(w2944) );
	vdp_slatch g3225 (.Q(w3247), .D(w4151), .C(w2946), .nC(w2947) );
	vdp_slatch g3226 (.Q(w3244), .D(w4150), .C(w2939), .nC(w2938) );
	vdp_slatch g3227 (.Q(w3279), .D(w4189), .nC(w3341), .C(w3340) );
	vdp_slatch g3228 (.Q(w3388), .D(w4188), .nC(w3344), .C(w3345) );
	vdp_slatch g3229 (.Q(w3281), .D(w4193), .nC(w3343), .C(w3342) );
	vdp_slatch g3230 (.Q(w3280), .D(w4192), .nC(w3347), .C(w3346) );
	vdp_slatch g3231 (.Q(w3387), .D(w4197), .nC(w3341), .C(w3340) );
	vdp_slatch g3232 (.Q(w3391), .D(w4196), .nC(w3344), .C(w3345) );
	vdp_slatch g3233 (.Q(w3390), .D(w4201), .nC(w3343), .C(w3342) );
	vdp_slatch g3234 (.Q(w3389), .D(w4200), .nC(w3347), .C(w3346) );
	vdp_slatch g3235 (.Q(w3282), .D(w4205), .nC(w3341), .C(w3340) );
	vdp_slatch g3236 (.Q(w3392), .D(w4204), .nC(w3344), .C(w3345) );
	vdp_slatch g3237 (.Q(w3386), .D(w4209), .nC(w3343), .C(w3342) );
	vdp_slatch g3238 (.Q(w3393), .D(w4208), .nC(w3347), .C(w3346) );
	vdp_slatch g3239 (.Q(w3394), .D(w4213), .nC(w3341), .C(w3340) );
	vdp_slatch g3240 (.Q(w3395), .D(w4212), .nC(w3344), .C(w3345) );
	vdp_slatch g3241 (.Q(w3283), .D(w4217), .nC(w3343), .C(w3342) );
	vdp_slatch g3242 (.Q(w3284), .D(w4216), .nC(w3347), .C(w3346) );
	vdp_slatch g3243 (.Q(w3378), .D(w4221), .nC(w3341), .C(w3340) );
	vdp_slatch g3244 (.Q(w3379), .D(w4220), .nC(w3344), .C(w3345) );
	vdp_slatch g3245 (.Q(w3380), .D(w4225), .nC(w3343), .C(w3342) );
	vdp_slatch g3246 (.Q(w3381), .D(w4224), .nC(w3347), .C(w3346) );
	vdp_slatch g3247 (.Q(w3382), .D(w4229), .nC(w3341), .C(w3340) );
	vdp_slatch g3248 (.Q(w3383), .D(w4228), .nC(w3344), .C(w3345) );
	vdp_slatch g3249 (.Q(w3384), .D(w4233), .nC(w3343), .C(w3342) );
	vdp_slatch g3250 (.Q(w3385), .D(w4232), .nC(w3347), .C(w3346) );
	vdp_slatch g3251 (.Q(w3377), .D(w4237), .nC(w3341), .C(w3340) );
	vdp_slatch g3252 (.Q(w3376), .D(w4236), .nC(w3344), .C(w3345) );
	vdp_slatch g3253 (.Q(w3375), .D(w4241), .nC(w3343), .C(w3342) );
	vdp_slatch g3254 (.Q(w3374), .D(w4240), .nC(w3347), .C(w3346) );
	vdp_slatch g3255 (.Q(w3373), .D(w4245), .nC(w3341), .C(w3340) );
	vdp_slatch g3256 (.Q(w3372), .D(w4244), .nC(w3344), .C(w3345) );
	vdp_slatch g3257 (.Q(w3370), .D(w4249), .nC(w3343), .C(w3342) );
	vdp_slatch g3258 (.Q(w3371), .D(w4248), .nC(w3347), .C(w3346) );
	vdp_slatch g3259 (.Q(w4189), .D(w4187), .C(w3305), .nC(w3339) );
	vdp_slatch g3260 (.Q(w4188), .D(w4186), .C(w3331), .nC(w3333) );
	vdp_slatch g3261 (.Q(w4193), .D(w4191), .C(w3306), .nC(w3334) );
	vdp_slatch g3262 (.Q(w4192), .D(w4190), .C(w3338), .nC(w3337) );
	vdp_slatch g3263 (.Q(w4197), .D(w4195), .C(w3305), .nC(w3339) );
	vdp_slatch g3264 (.Q(w4196), .D(w4194), .C(w3331), .nC(w3333) );
	vdp_slatch g3265 (.Q(w4201), .D(w4199), .C(w3306), .nC(w3334) );
	vdp_slatch g3266 (.Q(w4200), .D(w4198), .C(w3338), .nC(w3337) );
	vdp_slatch g3267 (.Q(w4205), .D(w4203), .C(w3305), .nC(w3339) );
	vdp_slatch g3268 (.Q(w4204), .D(w4202), .C(w3331), .nC(w3333) );
	vdp_slatch g3269 (.Q(w4209), .D(w4207), .C(w3306), .nC(w3334) );
	vdp_slatch g3270 (.Q(w4208), .D(w4206), .C(w3338), .nC(w3337) );
	vdp_slatch g3271 (.Q(w4213), .D(w4211), .C(w3305), .nC(w3339) );
	vdp_slatch g3272 (.Q(w4212), .D(w4210), .C(w3331), .nC(w3333) );
	vdp_slatch g3273 (.Q(w4217), .D(w4215), .C(w3306), .nC(w3334) );
	vdp_slatch g3274 (.Q(w4216), .D(w4214), .C(w3338), .nC(w3337) );
	vdp_slatch g3275 (.Q(w4221), .D(w4219), .C(w3305), .nC(w3339) );
	vdp_slatch g3276 (.Q(w4220), .D(w4218), .C(w3331), .nC(w3333) );
	vdp_slatch g3277 (.Q(w4225), .D(w4223), .C(w3306), .nC(w3334) );
	vdp_slatch g3278 (.Q(w4224), .D(w4222), .C(w3338), .nC(w3337) );
	vdp_slatch g3279 (.Q(w4229), .D(w4227), .C(w3305), .nC(w3339) );
	vdp_slatch g3280 (.Q(w4228), .D(w4226), .C(w3331), .nC(w3333) );
	vdp_slatch g3281 (.Q(w4233), .D(w4231), .C(w3306), .nC(w3334) );
	vdp_slatch g3282 (.Q(w4232), .D(w4230), .C(w3338), .nC(w3337) );
	vdp_slatch g3283 (.Q(w4237), .D(w4235), .C(w3305), .nC(w3339) );
	vdp_slatch g3284 (.Q(w4236), .D(w4234), .C(w3331), .nC(w3333) );
	vdp_slatch g3285 (.Q(w4241), .D(w4239), .C(w3306), .nC(w3334) );
	vdp_slatch g3286 (.Q(w4240), .D(w4238), .C(w3338), .nC(w3337) );
	vdp_slatch g3287 (.Q(w4245), .D(w4243), .C(w3305), .nC(w3339) );
	vdp_slatch g3288 (.Q(w4244), .D(w4242), .C(w3331), .nC(w3333) );
	vdp_slatch g3289 (.Q(w4249), .D(w4247), .C(w3306), .nC(w3334) );
	vdp_slatch g3290 (.Q(w4248), .D(w4246), .C(w3338), .nC(w3337) );
	vdp_slatch g3291 (.Q(w4187), .D(S[3]), .nC(w3332), .C(w3360) );
	vdp_slatch g3292 (.Q(w4186), .D(S[3]), .nC(w3348), .C(w3361) );
	vdp_slatch g3293 (.Q(w4191), .D(S[3]), .nC(w3335), .C(w3359) );
	vdp_slatch g3294 (.Q(w4190), .D(S[3]), .nC(w3336), .C(w3358) );
	vdp_slatch g3295 (.Q(w4195), .D(S[7]), .nC(w3332), .C(w3360) );
	vdp_slatch g3296 (.Q(w4194), .D(S[7]), .nC(w3348), .C(w3361) );
	vdp_slatch g3297 (.Q(w4199), .D(S[7]), .nC(w3335), .C(w3359) );
	vdp_slatch g3298 (.Q(w4198), .D(S[7]), .nC(w3336), .C(w3358) );
	vdp_slatch g3299 (.Q(w4203), .D(S[2]), .nC(w3332), .C(w3360) );
	vdp_slatch g3300 (.Q(w4202), .D(S[2]), .nC(w3348), .C(w3361) );
	vdp_slatch g3301 (.Q(w4207), .D(S[2]), .nC(w3335), .C(w3359) );
	vdp_slatch g3302 (.Q(w4206), .D(S[2]), .nC(w3336), .C(w3358) );
	vdp_slatch g3303 (.Q(w4211), .D(S[6]), .nC(w3332), .C(w3360) );
	vdp_slatch g3304 (.Q(w4210), .D(S[6]), .nC(w3348), .C(w3361) );
	vdp_slatch g3305 (.Q(w4215), .D(S[6]), .nC(w3335), .C(w3359) );
	vdp_slatch g3306 (.Q(w4214), .D(S[6]), .nC(w3336), .C(w3358) );
	vdp_slatch g3307 (.Q(w4219), .D(S[1]), .nC(w3332), .C(w3360) );
	vdp_slatch g3308 (.Q(w4218), .D(S[1]), .nC(w3348), .C(w3361) );
	vdp_slatch g3309 (.Q(w4223), .D(S[1]), .nC(w3335), .C(w3359) );
	vdp_slatch g3310 (.Q(w4222), .D(S[1]), .nC(w3336), .C(w3358) );
	vdp_slatch g3311 (.Q(w4227), .D(S[5]), .nC(w3332), .C(w3360) );
	vdp_slatch g3312 (.Q(w4226), .D(S[5]), .nC(w3348), .C(w3361) );
	vdp_slatch g3313 (.Q(w4231), .D(S[5]), .nC(w3335), .C(w3359) );
	vdp_slatch g3314 (.Q(w4230), .D(S[5]), .nC(w3336), .C(w3358) );
	vdp_slatch g3315 (.Q(w4235), .D(S[0]), .nC(w3332), .C(w3360) );
	vdp_slatch g3316 (.Q(w4234), .D(S[0]), .nC(w3348), .C(w3361) );
	vdp_slatch g3317 (.Q(w4239), .D(S[0]), .nC(w3335), .C(w3359) );
	vdp_slatch g3318 (.Q(w4238), .D(S[0]), .nC(w3336), .C(w3358) );
	vdp_slatch g3319 (.Q(w4243), .D(S[4]), .nC(w3332), .C(w3360) );
	vdp_slatch g3320 (.Q(w4242), .D(S[4]), .nC(w3348), .C(w3361) );
	vdp_slatch g3321 (.Q(w4247), .D(S[4]), .nC(w3335), .C(w3359) );
	vdp_slatch g3322 (.Q(w4246), .D(S[4]), .nC(w3336), .C(w3358) );
	vdp_aon2x8 g3323 (.Z(w3890), .A1(w3077), .B1(w3076), .C1(w3075), .D2(w3074), .A2(w3121), .B2(w3122), .C2(w3127), .D1(w3126), .E2(w3124), .F1(w3125), .E1(w3073), .F2(w3072), .G1(w3071), .H2(w3070), .G2(w3129), .H1(w3119) );
	vdp_aon2x8 g3324 (.Z(w3101), .A1(w3195), .B1(w3122), .C1(w3197), .D2(w3126), .A2(w3121), .B2(w3196), .C2(w3127), .D1(w3198), .E2(w3124), .F1(w3125), .E1(w3199), .F2(w3200), .G1(w3206), .H2(w3207), .G2(w3129), .H1(w3119) );
	vdp_aon2x8 g3325 (.Z(w3104), .A1(w3069), .B1(w3082), .C1(w3086), .D2(w3085), .A2(w3121), .B2(w3122), .C2(w3127), .D1(w3126), .E2(w3124), .F1(w3125), .E1(w3084), .F2(w3080), .G1(w3081), .H2(w3083), .G2(w3129), .H1(w3119) );
	vdp_aon2x8 g3326 (.Z(w3105), .A1(w3208), .B1(w3122), .C1(w3210), .D2(w3126), .A2(w3121), .B2(w3209), .C2(w3127), .D1(w3205), .E2(w3124), .F1(w3125), .E1(w3211), .F2(w3212), .G1(w3213), .H2(w3214), .G2(w3129), .H1(w3119) );
	vdp_aon2x8 g3327 (.Z(w3103), .A1(w3139), .B1(w3122), .C1(w3141), .D2(w3142), .A2(w3121), .B2(w3891), .C2(w3127), .D1(w3126), .E2(w3124), .F1(w3125), .E1(w3215), .F2(w3140), .G1(w3120), .H2(w3143), .G2(w3129), .H1(w3119) );
	vdp_aon2x8 g3328 (.Z(w3106), .A1(w3146), .B1(w3122), .C1(w3153), .D2(w3152), .A2(w3121), .B2(w3154), .C2(w3127), .D1(w3126), .E2(w3124), .F1(w3125), .E1(w3150), .F2(w3144), .G1(w3151), .G2(w3129), .H1(w3119), .H2(w3145) );
	vdp_aon2x8 g3329 (.Z(w3102), .A1(w3087), .B1(w3088), .C1(w3090), .D2(w3089), .A2(w3121), .B2(w3122), .C2(w3127), .D1(w3126), .E2(w3124), .F1(w3125), .E1(w3131), .F2(w3132), .G1(w3128), .H2(w3123), .G2(w3129), .H1(w3119) );
	vdp_aon2x8 g3330 (.Z(w3107), .A1(w3135), .B1(w3134), .C1(w3133), .D2(w3130), .A2(w3121), .B2(w3122), .C2(w3127), .D1(w3126), .E2(w3124), .F1(w3125), .E1(w3116), .F2(w3115), .G1(w3117), .H2(w3118), .G2(w3129), .H1(w3119) );
	vdp_aon2x8 g3331 (.A1(w3261), .B1(w3260), .C1(w3248), .D2(w3246), .A2(w3278), .B2(w3277), .C2(w3276), .D1(w3275), .E2(w3274), .F1(w3273), .E1(w3259), .F2(w3258), .G1(w3257), .H2(w3245), .G2(w3271), .H1(w3272), .Z(w3290) );
	vdp_aon2x8 g3332 (.Z(w3318), .A1(w3256), .B1(w3255), .C1(w3254), .D2(w3253), .A2(w3278), .B2(w3277), .C2(w3276), .D1(w3275), .E2(w3274), .F1(w3273), .E1(w3252), .F2(w3251), .G1(w3250), .H2(w3249), .G2(w3271), .H1(w3272) );
	vdp_aon2x8 g3333 (.Z(w3289), .A1(w3248), .B1(w3257), .C1(w3254), .D2(w3250), .A2(w3273), .B2(w3272), .C2(w3277), .D1(w3275), .E2(w3274), .F1(w3271), .E1(w3242), .F2(w3292), .G1(w3293), .H2(w3247), .G2(w3278), .H1(w3276) );
	vdp_aon2x8 g3334 (.Z(w3321), .A1(w3241), .B1(w3287), .C1(w3242), .D2(w3243), .A2(w3278), .B2(w3277), .C2(w3276), .D1(w3275), .E2(w3274), .F1(w3273), .E1(w3291), .F2(w3300), .G1(w3292), .H2(w3299), .G2(w3271), .H1(w3272) );
	vdp_aon2x8 g3335 (.Z(w3288), .A1(w3298), .B1(w3297), .C1(w3293), .D2(w3296), .A2(w3278), .B2(w3277), .C2(w3276), .D1(w3275), .E2(w3274), .F1(w3273), .E1(w3295), .F2(w3294), .G1(w3247), .H2(w3244), .G2(w3271), .H1(w3272) );
	vdp_aon2x8 g3336 (.Z(w3323), .A1(w3377), .B1(w3277), .C1(w3375), .D2(w3275), .A2(w3278), .B2(w3376), .C2(w3276), .D1(w3374), .E2(w3274), .F1(w3273), .E1(w3373), .F2(w3372), .G1(w3370), .H2(w3371), .G2(w3271), .H1(w3272) );
	vdp_aon2x8 g3337 (.Z(w3324), .A1(w3378), .B1(w3277), .C1(w3380), .D2(w3275), .A2(w3278), .B2(w3379), .C2(w3276), .D1(w3381), .E2(w3274), .F1(w3273), .E1(w3382), .F2(w3383), .G1(w3384), .H2(w3385), .G2(w3271), .H1(w3272) );
	vdp_aon2x8 g3338 (.Z(w3322), .A1(w3246), .B1(w3245), .C1(w3253), .D2(w3249), .A2(w3273), .B2(w3272), .C2(w3277), .D1(w3275), .E2(w3274), .F1(w3271), .E1(w3243), .F2(w3299), .G1(w3296), .H2(w3244), .G2(w3278), .H1(w3276) );
	vdp_aon2x8 g3339 (.Z(w3317), .A1(w3280), .B1(w3272), .C1(w3393), .D2(w3275), .A2(w3273), .B2(w3389), .C2(w3277), .D1(w3284), .E2(w3274), .F1(w3271), .E1(w3381), .F2(w3385), .G1(w3374), .H2(w3371), .G2(w3278), .H1(w3276) );
	vdp_aon2x8 g3340 (.Z(w3320), .A1(w3281), .B1(w3272), .C1(w3386), .D2(w3275), .A2(w3273), .B2(w3390), .C2(w3277), .D1(w3283), .E2(w3274), .F1(w3271), .E1(w3380), .F2(w3384), .G1(w3375), .H2(w3370), .G2(w3278), .H1(w3276) );
	vdp_aon2x8 g3341 (.Z(w3319), .A1(w3282), .B1(w3277), .C1(w3386), .D2(w3275), .A2(w3278), .B2(w3392), .C2(w3276), .D1(w3393), .E2(w3274), .F1(w3273), .E1(w3394), .F2(w3395), .G1(w3283), .H2(w3284), .G2(w3271), .H1(w3272) );
	vdp_aon2x8 g3342 (.A1(w3279), .B1(w3277), .C1(w3281), .D2(w3275), .A2(w3278), .B2(w3388), .C2(w3276), .D1(w3280), .E2(w3274), .F1(w3273), .E1(w3387), .F2(w3391), .G1(w3390), .H2(w3389), .G2(w3271), .H1(w3272), .Z(w3325) );
	vdp_sr_bit g3343 (.Q(w3268), .D(w3411), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3344 (.Q(w3411), .D(w3327), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3345 (.Q(w3328), .D(w3412), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3346 (.Q(w3412), .D(w3330), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3347 (.Q(w3329), .D(w3304), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3348 (.Q(w3918), .D(w3329), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3349 (.Q(w3396), .D(w3326), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3350 (.Q(w3303), .D(w3396), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3351 (.Q(w3920), .D(w3313), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3352 (.Q(w3302), .D(w3920), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3353 (.Q(w3301), .D(w3269), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3354 (.Q(w3269), .D(w3312), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3355 (.Q(w2728), .D(w3314), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3356 (.Q(w3397), .D(w2728), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3357 (.Q(w3093), .D(w3111), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3358 (.Q(w3095), .D(w3093), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3359 (.Q(w3098), .D(w3094), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3360 (.Q(w3094), .D(w3110), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3361 (.Q(w3109), .D(w3091), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3362 (.Q(w3091), .D(w3112), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3363 (.Q(w3092), .D(w3108), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3364 (.Q(w3100), .D(w3092), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3365 (.Q(w3178), .D(w2727), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3366 (.Q(w2727), .D(w3177), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3367 (.Q(w3901), .D(w3113), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3368 (.Q(w3099), .D(w3901), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3369 (.Q(w3900), .D(w3176), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3370 (.Q(w3097), .D(w3900), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3371 (.Q(w3025), .D(VRAMA[1]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3372 (.Q(w3057), .D(VRAMA[2]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3373 (.Q(w3059), .D(VRAMA[3]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3374 (.Q(w3060), .D(VRAMA[4]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3375 (.Q(w3061), .D(VRAMA[5]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3376 (.Q(w3062), .D(VRAMA[6]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3377 (.Q(w3898), .D(w3048), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3378 (.Q(w3398), .D(w3898), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3379 (.Q(w3047), .D(w3399), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3380 (.Q(w3399), .D(w3398), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_dlatch_inv g3381 (.nQ(w3048), .D(w3012), .C(DCLK1), .nC(nDCLK1) );
	vdp_slatch g3382 (.Q(w3170), .D(w4251), .C(w3163), .nC(w2926) );
	vdp_slatch g3383 (.Q(w3169), .D(w4252), .C(w3163), .nC(w2926) );
	vdp_slatch g3384 (.Q(w3168), .D(w4253), .C(w3163), .nC(w2926) );
	vdp_slatch g3385 (.Q(w3167), .D(w4254), .C(w3163), .nC(w2926) );
	vdp_slatch g3386 (.Q(w3166), .D(w4255), .C(w3163), .nC(w2926) );
	vdp_slatch g3387 (.Q(w3165), .D(w4256), .C(w3163), .nC(w2926) );
	vdp_slatch g3388 (.Q(w3164), .D(w4258), .C(w3163), .nC(w2926) );
	vdp_slatch g3389 (.Q(w2927), .D(w4257), .C(w3163), .nC(w2926) );
	vdp_slatch g3390 (.Q(w4251), .D(w2993), .C(w3185), .nC(w3217) );
	vdp_slatch g3391 (.Q(w4252), .D(w2968), .C(w3185), .nC(w3217) );
	vdp_slatch g3392 (.Q(w4253), .D(w2970), .C(w3185), .nC(w3217) );
	vdp_slatch g3393 (.Q(w4254), .D(w2971), .C(w3185), .nC(w3217) );
	vdp_slatch g3394 (.Q(w4255), .D(w2972), .C(w3185), .nC(w3217) );
	vdp_slatch g3395 (.Q(w4256), .D(w2994), .C(w3185), .nC(w3217) );
	vdp_slatch g3396 (.Q(w4258), .D(w2998), .C(w3185), .nC(w3217) );
	vdp_slatch g3397 (.Q(w4257), .D(w2997), .C(w3185), .nC(w3217) );
	vdp_slatch g3398 (.Q(w4259), .D(w2934), .C(w2936), .nC(w2935) );
	vdp_slatch g3399 (.Q(w4260), .D(w2967), .C(w2936), .nC(w2935) );
	vdp_slatch g3400 (.Q(w4261), .D(w2933), .C(w2936), .nC(w2935) );
	vdp_slatch g3401 (.Q(w4262), .D(w3950), .C(w2936), .nC(w2935) );
	vdp_slatch g3402 (.Q(w4263), .D(w3407), .C(w2936), .nC(w2935) );
	vdp_slatch g3403 (.Q(w4264), .D(w2974), .C(w2936), .nC(w2935) );
	vdp_slatch g3404 (.Q(w4265), .D(w2930), .C(w2936), .nC(w2935) );
	vdp_slatch g3405 (.Q(w4266), .D(w2975), .C(w2936), .nC(w2935) );
	vdp_slatch g3406 (.Q(w3226), .D(w4259), .C(w2937), .nC(w3219) );
	vdp_slatch g3407 (.Q(w3225), .D(w4260), .C(w2937), .nC(w3219) );
	vdp_slatch g3408 (.Q(w3224), .D(w4261), .C(w2937), .nC(w3219) );
	vdp_slatch g3409 (.Q(w3223), .D(w4262), .C(w2937), .nC(w3219) );
	vdp_slatch g3410 (.Q(w3222), .D(w4263), .C(w2937), .nC(w3219) );
	vdp_slatch g3411 (.Q(w3221), .D(w4264), .C(w2937), .nC(w3219) );
	vdp_slatch g3412 (.Q(w3220), .D(w4265), .C(w2937), .nC(w3219) );
	vdp_slatch g3413 (.Q(w4288), .D(w4266), .C(w2937), .nC(w3219) );
	vdp_slatch g3414 (.Q(w3362), .D(w3356), .C(w3045), .nC(w3353) );
	vdp_slatch g3415 (.Q(w3355), .D(w3052), .C(w3045), .nC(w3353) );
	vdp_slatch g3416 (.Q(w3737), .D(w3354), .C(w3045), .nC(w3353) );
	vdp_slatch g3417 (.Q(w3349), .D(w3352), .C(w3045), .nC(w3353) );
	vdp_slatch g3418 (.Q(w2934), .D(w2993), .C(w2996), .nC(w2995) );
	vdp_slatch g3419 (.Q(w2967), .D(w2968), .C(w2996), .nC(w2995) );
	vdp_slatch g3420 (.Q(w2933), .D(w2970), .C(w2996), .nC(w2995) );
	vdp_slatch g3421 (.Q(w3950), .D(w2971), .C(w2996), .nC(w2995) );
	vdp_slatch g3422 (.Q(w3407), .D(w2972), .C(w2996), .nC(w2995) );
	vdp_slatch g3423 (.Q(w2974), .D(w2994), .C(w2996), .nC(w2995) );
	vdp_slatch g3424 (.Q(w2930), .D(w2998), .C(w2996), .nC(w2995) );
	vdp_slatch g3425 (.Q(w2975), .D(w2997), .C(w2996), .nC(w2995) );
	vdp_cnt_bit_load g3426 (.D(w3354), .nL(w3016), .L(w3013), .R(1'b0), .Q(w3015), .CI(w3403), .CO(w3404), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3427 (.D(w3052), .nL(w3016), .L(w3013), .R(1'b0), .Q(w3889), .CI(w3404), .CO(w3405), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3428 (.D(w3017), .nL(w3016), .L(w3013), .R(1'b0), .Q(w3001), .CI(w3405), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3429 (.CO(w3403), .CI(1'b1), .D(w3352), .nL(w3016), .L(w3013), .R(1'b0), .Q(w3011), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3430 (.CO(w3402), .CI(1'b1), .D(w3349), .nL(w3351), .L(w3044), .R(1'b0), .Q(w3369), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3431 (.CO(w3401), .CI(w3402), .D(w3737), .nL(w3351), .L(w3044), .R(1'b0), .Q(w3315), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3432 (.CO(w3400), .CI(w3401), .D(w3355), .nL(w3351), .L(w3044), .R(1'b0), .Q(w3357), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3433 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .CI(w3400), .D(w3362), .nL(w3351), .L(w3044), .R(1'b0), .Q(w3267) );
	vdp_xor g3434 (.Z(w3155), .B(w3889), .A(w3010) );
	vdp_xor g3435 (.B(w3015), .A(w3010), .Z(w3002) );
	vdp_xor g3436 (.Z(w3158), .B(w3011), .A(w3010) );
	vdp_sr_bit g3437 (.Q(w3009), .D(w3896), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3438 (.Q(w3895), .D(w3009), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3439 (.Q(w3175), .D(w3895), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3440 (.Q(w3904), .D(w3406), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3441 (.Q(w3406), .D(w3905), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3442 (.Q(w3905), .D(w3906), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3443 (.Q(w2932), .D(w2931), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3444 (.Q(w2931), .D(w2929), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3445 (.Q(w2929), .D(w2928), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3446 (.Q(w3908), .D(w3909), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3447 (.Q(w3877), .D(w3908), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3448 (.Q(w3907), .D(w3877), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3449 (.Q(w3912), .D(w3911), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3450 (.Q(w3913), .D(w3912), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3451 (.Q(w3910), .D(w3913), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3452 (.Q(w3023), .D(w3910), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3453 (.Q(w3991), .D(w3992), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3454 (.Q(w3992), .D(w3914), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_xor g3455 (.Z(w3229), .A(w3311), .B(w3357) );
	vdp_xor g3456 (.Z(w3234), .A(w3311), .B(w3368) );
	vdp_xor g3457 (.Z(w3228), .A(w3311), .B(w3369) );
	vdp_dlatch_inv g3458 (.nQ(w3894), .D(w3893), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g3459 (.nQ(w2928), .D(w2973), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g3460 (.nQ(w3909), .D(w2924), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g3461 (.nQ(w3367), .D(w3915), .nC(nHCLK1), .C(HCLK1) );
	vdp_xor g3462 (.Z(w3368), .A(w3315), .B(M5) );
	vdp_sr_bit g3463 (.Q(w3409), .D(w3316), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_dlatch_inv g3464 (.nQ(w3911), .D(w3021), .nC(nDCLK1), .C(DCLK1) );
	vdp_comp_strong g3465 (.Z(w2941), .nZ(w2942), .A(w3218) );
	vdp_comp_strong g3466 (.Z(w2949), .nZ(w2944), .A(w3218) );
	vdp_comp_strong g3467 (.Z(w2946), .nZ(w2947), .A(w3218) );
	vdp_comp_strong g3468 (.Z(w2939), .nZ(w2938), .A(w3218) );
	vdp_comp_strong g3469 (.Z(w2940), .nZ(w2979), .A(w3024) );
	vdp_comp_strong g3470 (.Z(w2943), .nZ(w2980), .A(w3024) );
	vdp_comp_strong g3471 (.Z(w2948), .nZ(w2981), .A(w3024) );
	vdp_comp_strong g3472 (.Z(w2945), .nZ(w2950), .A(w3024) );
	vdp_comp_strong g3473 (.Z(w2953), .nZ(w2977), .A(w2976) );
	vdp_comp_strong g3474 (.Z(w2957), .nZ(w2982), .A(w3286) );
	vdp_comp_strong g3475 (.Z(w2958), .nZ(w2983), .A(w3285) );
	vdp_comp_strong g3476 (.Z(w2960), .nZ(w2978), .A(w2969) );
	vdp_comp_strong g3477 (.Z(w2952), .nZ(w2985), .A(w3903) );
	vdp_comp_strong g3478 (.Z(w2956), .nZ(w2989), .A(w2990) );
	vdp_comp_strong g3479 (.Z(w2959), .nZ(w2986), .A(w2992) );
	vdp_comp_strong g3480 (.Z(w2961), .nZ(w2984), .A(w2991) );
	vdp_comp_strong g3481 (.Z(w3192), .nZ(w3179), .A(w2925) );
	vdp_comp_strong g3482 (.Z(w2999), .nZ(w3180), .A(w2925) );
	vdp_comp_strong g3483 (.Z(w3186), .nZ(w2987), .A(w2925) );
	vdp_comp_strong g3484 (.Z(w3187), .nZ(w2988), .A(w2925) );
	vdp_comp_strong g3485 (.Z(w3191), .nZ(w3193), .A(w3000) );
	vdp_comp_strong g3486 (.Z(w3190), .nZ(w3201), .A(w3000) );
	vdp_comp_strong g3487 (.Z(w3189), .nZ(w3202), .A(w3000) );
	vdp_comp_strong g3488 (.Z(w3188), .nZ(w3194), .A(w3000) );
	vdp_comp_strong g3489 (.Z(w3042), .nZ(w3068), .A(w3000) );
	vdp_comp_strong g3490 (.Z(w3020), .nZ(w3078), .A(w3000) );
	vdp_comp_strong g3491 (.Z(w3033), .nZ(w3079), .A(w3000) );
	vdp_comp_strong g3492 (.Z(w3034), .nZ(w3007), .A(w3000) );
	vdp_comp_strong g3493 (.Z(w3019), .nZ(w3037), .A(w2925) );
	vdp_comp_strong g3494 (.Z(w3038), .nZ(w3029), .A(w2925) );
	vdp_comp_strong g3495 (.Z(w3039), .nZ(w3027), .A(w2925) );
	vdp_comp_strong g3496 (.Z(w3035), .nZ(w3036), .A(w2925) );
	vdp_comp_strong g3497 (.Z(w3050), .nZ(w3040), .A(w3051) );
	vdp_comp_strong g3498 (.Z(w3031), .nZ(w3030), .A(w3053) );
	vdp_comp_strong g3499 (.Z(w3032), .nZ(w3028), .A(w3054) );
	vdp_comp_strong g3500 (.Z(w3049), .nZ(w3041), .A(w3055) );
	vdp_comp_strong g3501 (.Z(w3360), .nZ(w3332), .A(w3173) );
	vdp_comp_strong g3502 (.Z(w3361), .nZ(w3348), .A(w3363) );
	vdp_comp_strong g3503 (.Z(w3359), .nZ(w3335), .A(w3364) );
	vdp_comp_strong g3504 (.Z(w3358), .nZ(w3336), .A(w3365) );
	vdp_comp_strong g3505 (.Z(w3305), .nZ(w3339), .A(w3024) );
	vdp_comp_strong g3506 (.Z(w3331), .nZ(w3333), .A(w3024) );
	vdp_comp_strong g3507 (.Z(w3306), .nZ(w3334), .A(w3024) );
	vdp_comp_strong g3508 (.Z(w3338), .nZ(w3337), .A(w3024) );
	vdp_comp_strong g3509 (.Z(w3340), .nZ(w3341), .A(w3218) );
	vdp_comp_strong g3510 (.Z(w3345), .nZ(w3344), .A(w3218) );
	vdp_comp_strong g3511 (.Z(w3342), .nZ(w3343), .A(w3218) );
	vdp_comp_strong g3512 (.Z(w3346), .nZ(w3347), .A(w3218) );
	vdp_not g3513 (.nZ(w3017), .A(w3356) );
	vdp_not g3514 (.nZ(w3896), .A(w3136) );
	vdp_not g3515 (.nZ(w3138), .A(w91) );
	vdp_not g3516 (.nZ(w3137), .A(w428) );
	vdp_not g3517 (.nZ(w3003), .A(w3137) );
	vdp_comp_strong g3518 (.Z(w3163), .nZ(w2926), .A(w3000) );
	vdp_comp_strong g3519 (.Z(w3185), .nZ(w3217), .A(w2925) );
	vdp_comp_strong g3520 (.Z(w2996), .nZ(w2995), .A(w3173) );
	vdp_comp_strong g3521 (.Z(w2937), .nZ(w3219), .A(w3218) );
	vdp_comp_strong g3522 (.Z(w2936), .nZ(w2935), .A(w3024) );
	vdp_comp_strong g3523 (.Z(w3045), .nZ(w3353), .A(w3409) );
	vdp_not g3524 (.nZ(w3235), .A(w3228) );
	vdp_not g3525 (.nZ(w3227), .A(w3234) );
	vdp_not g3526 (.nZ(w3238), .A(w3229) );
	vdp_nand3 g3527 (.Z(w3232), .A(w3238), .B(w3234), .C(w3228) );
	vdp_not g3528 (.nZ(w3277), .A(w3231) );
	vdp_nand3 g3529 (.Z(w3231), .A(w3229), .B(w3227), .C(w3228) );
	vdp_nand3 g3530 (.Z(w3230), .A(w3229), .B(w3234), .C(w3228) );
	vdp_nand3 g3531 (.Z(w3236), .A(w3229), .B(w3234), .C(w3235) );
	vdp_nand3 g3532 (.Z(w3233), .A(w3238), .B(w3227), .C(w3228) );
	vdp_nand3 g3533 (.Z(w3239), .A(w3238), .B(w3234), .C(w3235) );
	vdp_nand3 g3534 (.Z(w3237), .A(w3229), .B(w3227), .C(w3235) );
	vdp_nand3 g3535 (.Z(w3240), .A(w3235), .B(w3238), .C(w3227) );
	vdp_not g3536 (.nZ(w3278), .A(w3230) );
	vdp_not g3537 (.nZ(w3276), .A(w3232) );
	vdp_not g3538 (.nZ(w3275), .A(w3233) );
	vdp_not g3539 (.nZ(w3273), .A(w3237) );
	vdp_not g3540 (.nZ(w3274), .A(w3236) );
	vdp_not g3541 (.nZ(w3272), .A(w3240) );
	vdp_not g3542 (.nZ(w3271), .A(w3239) );
	vdp_not g3543 (.nZ(w3148), .A(w3158) );
	vdp_not g3544 (.nZ(w3156), .A(w3008) );
	vdp_not g3545 (.nZ(w3147), .A(w3155) );
	vdp_nand3 g3546 (.Z(w3160), .A(w3147), .B(w3008), .C(w3158) );
	vdp_not g3547 (.nZ(w3122), .A(w3162) );
	vdp_nand3 g3548 (.Z(w3162), .A(w3155), .B(w3156), .C(w3158) );
	vdp_nand3 g3549 (.Z(w3161), .A(w3155), .B(w3008), .C(w3158) );
	vdp_nand3 g3550 (.Z(w3902), .A(w3155), .B(w3008), .C(w3148) );
	vdp_nand3 g3551 (.Z(w3159), .A(w3147), .B(w3156), .C(w3158) );
	vdp_nand3 g3552 (.Z(w3157), .A(w3155), .B(w3156), .C(w3148) );
	vdp_not g3553 (.nZ(w3121), .A(w3161) );
	vdp_not g3554 (.nZ(w3127), .A(w3160) );
	vdp_not g3555 (.nZ(w3126), .A(w3159) );
	vdp_not g3556 (.nZ(w3125), .A(w3157) );
	vdp_not g3557 (.nZ(w3124), .A(w3902) );
	vdp_aon22 g3558 (.Z(w3177), .A1(w3164), .B1(w3171), .A2(w3172), .B2(w2927) );
	vdp_aon22 g3559 (.Z(w3176), .A1(w3166), .B1(w3171), .A2(w3172), .B2(w3165) );
	vdp_aon22 g3560 (.Z(w3113), .A1(w3168), .B1(w3171), .A2(w3172), .B2(w3167) );
	vdp_aon22 g3561 (.Z(w3010), .A1(w3170), .B1(w3171), .A2(w3172), .B2(w3169) );
	vdp_sr_bit g3562 (.Q(w3006), .D(w3897), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3563 (.Q(w3897), .D(w3005), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_xor g3564 (.Z(w3008), .A(w3002), .B(1'b1) );
	vdp_xor g3565 (.A(HPOS[3]), .B(w3026), .Z(w3949) );
	vdp_aon22 g3566 (.Z(w3064), .A1(w3057), .B1(w3058), .A2(w3056), .B2(w3948) );
	vdp_aon22 g3567 (.Z(w3065), .A1(w3059), .B1(w3058), .A2(w3056), .B2(w3947) );
	vdp_aon22 g3568 (.Z(w3067), .A1(w3060), .B1(w3058), .A2(w3056), .B2(w3946) );
	vdp_aon22 g3569 (.Z(w3066), .A1(w3061), .B1(w3058), .A2(w3056), .B2(w3945) );
	vdp_aon22 g3570 (.Z(w3490), .A1(w3062), .B1(w3058), .A2(w3056), .B2(w3944) );
	vdp_aon22 g3571 (.Z(w3108), .A1(w3204), .B1(w3890), .A2(w3101), .B2(w3203) );
	vdp_aon22 g3572 (.Z(w3112), .A1(w3204), .B1(w3102), .A2(w3103), .B2(w3203) );
	vdp_aon22 g3573 (.Z(w3110), .A1(w3204), .B1(w3107), .A2(w3106), .B2(w3203) );
	vdp_aon22 g3574 (.Z(w3111), .A1(w3204), .B1(w3104), .A2(w3105), .B2(w3203) );
	vdp_aon222 g3575 (.Z(w3327), .A1(w3319), .B1(w3318), .C1(w3317), .A2(w3265), .B2(w3266), .C2(w3264) );
	vdp_aon222 g3576 (.Z(w3330), .A1(w3323), .B1(w3288), .C1(w3322), .A2(w3265), .B2(w3266), .C2(w3264) );
	vdp_aon222 g3577 (.Z(w3304), .A1(w3324), .B1(w3321), .C1(w3289), .A2(w3265), .B2(w3266), .C2(w3264) );
	vdp_aon222 g3578 (.A1(w3325), .B1(w3290), .C1(w3320), .A2(w3265), .B2(w3266), .C2(w3264), .Z(w3326) );
	vdp_and5 g3579 (.Z(w3366), .A(w3316), .B(w3362), .C(w3355), .D(w3737), .E(w3349) );
	vdp_aon22 g3580 (.Z(w3313), .A1(w3222), .B1(w3410), .A2(w3043), .B2(w3221) );
	vdp_aon22 g3581 (.Z(w3312), .A1(w3224), .B1(w3410), .A2(w3043), .B2(w3223) );
	vdp_aon22 g3582 (.Z(w3311), .A1(w3226), .B1(w3410), .A2(w3043), .B2(w3225) );
	vdp_aon22 g3583 (.Z(w3314), .A1(w3220), .B1(w3410), .A2(w3043), .B2(w4288) );
	vdp_aon22 g3584 (.Z(w3022), .A1(w3308), .B1(w3047), .A2(w3023), .B2(M5) );
	vdp_and4 g3585 (.Z(w3309), .A(w3369), .B(w3315), .C(w3357), .D(w3310) );
	vdp_comp_we g3586 (.Z(w3043), .nZ(w3410), .A(w3307) );
	vdp_comp_we g3587 (.Z(w3203), .nZ(w3204), .A(w3001) );
	vdp_comp_we g3588 (.Z(w3172), .nZ(w3171), .A(w3001) );
	vdp_comp_we g3589 (.Z(w3013), .nZ(w3016), .A(w3096) );
	vdp_comp_we g3590 (.Z(w3056), .nZ(w3058), .A(w3577) );
	vdp_comp_we g3591 (.Z(w3044), .nZ(w3351), .A(w3316) );
	vdp_not g3592 (.nZ(w3916), .A(M5) );
	vdp_dlatch_inv g3593 (.nQ(w3906), .D(w3018), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g3594 (.Z(w3183), .A(DCLK2), .B(w2929) );
	vdp_and g3595 (.Z(w3184), .A(DCLK2), .B(w2928) );
	vdp_and g3596 (.Z(w3182), .A(DCLK2), .B(w2931) );
	vdp_and g3597 (.Z(w3181), .A(DCLK2), .B(w2932) );
	vdp_and g3598 (.Z(w2991), .A(w3906), .B(DCLK2) );
	vdp_and g3599 (.Z(w2992), .A(w3905), .B(DCLK2) );
	vdp_and g3600 (.Z(w2990), .A(w3406), .B(DCLK2) );
	vdp_and g3601 (.Z(w3903), .A(w3904), .B(DCLK2) );
	vdp_and g3602 (.Z(w2976), .A(DCLK2), .B(w3907) );
	vdp_and g3603 (.Z(w3286), .A(DCLK2), .B(w3877) );
	vdp_and g3604 (.Z(w3285), .A(DCLK2), .B(w3908) );
	vdp_and g3605 (.Z(w2969), .A(DCLK2), .B(w3909) );
	vdp_and g3606 (.Z(w3000), .A(w3894), .B(HCLK2) );
	vdp_and g3607 (.Z(w3174), .A(w3138), .B(w3009) );
	vdp_and g3608 (.Z(w3218), .A(w3367), .B(HCLK2) );
	vdp_or g3609 (.Z(w3310), .A(w3916), .B(w3267) );
	vdp_and g3610 (.Z(w3024), .A(w3022), .B(DCLK2) );
	vdp_and g3611 (.Z(w3365), .A(DCLK2), .B(w3911) );
	vdp_and g3612 (.Z(w3364), .A(DCLK2), .B(w3912) );
	vdp_and g3613 (.Z(w3363), .A(DCLK2), .B(w3913) );
	vdp_and g3614 (.Z(w3173), .A(DCLK2), .B(w3910) );
	vdp_and g3615 (.Z(w3307), .A(M5), .B(w3267) );
	vdp_and g3616 (.Z(w3945), .A(VSCR), .B(HPOS[7]) );
	vdp_and g3617 (.Z(w3944), .A(VSCR), .B(HPOS[8]) );
	vdp_and g3618 (.Z(w3055), .A(DCLK2), .B(w3048) );
	vdp_and g3619 (.Z(w3946), .A(VSCR), .B(HPOS[6]) );
	vdp_and g3620 (.Z(w3054), .A(DCLK2), .B(w3898) );
	vdp_and g3621 (.Z(w3053), .A(DCLK2), .B(w3398) );
	vdp_and g3622 (.Z(w3051), .A(DCLK2), .B(w3399) );
	vdp_and g3623 (.Z(w3947), .A(VSCR), .B(HPOS[5]) );
	vdp_and g3624 (.Z(w2925), .A(DCLK2), .B(w3047) );
	vdp_and g3625 (.Z(w3948), .A(VSCR), .B(HPOS[4]) );
	vdp_aon22 g3626 (.Z(w3063), .A1(w3025), .B1(w3058), .A2(w3056), .B2(w3949) );
	vdp_and g3627 (.nZ(w3026), .A(VSCR), .B(M5) );
	vdp_or4 g3628 (.Z(w2873), .D(w3091), .C(w3092), .B(w3093), .A(w3094) );
	vdp_or g3629 (.Z(w3096), .A(w80), .B(w14) );
	vdp_or g3630 (.Z(w3316), .A(w9), .B(w78) );
	vdp_or4 g3631 (.Z(w2874), .A(w3412), .B(w3411), .C(w3396), .D(w3329) );
	vdp_not g3632 (.nZ(w3914), .A(w3270) );
	vdp_not g3633 (.nZ(w3005), .A(w3114) );
	vdp_not g3634 (.nZ(w3308), .A(M5) );
	vdp_aoi21 g3635 (.Z(w3270), .A1(w93), .A2(w3003), .B(w16) );
	vdp_aoi21 g3636 (.Z(w3114), .A1(w94), .A2(w3003), .B(w10) );
	vdp_aoi21 g3637 (.Z(w3136), .A1(w91), .A2(w3003), .B(w11) );
	vdp_nand4 g3638 (.D(w3001), .C(w3011), .Z(w3893), .A(w3889), .B(w3015) );
	vdp_nand3 g3639 (.Z(w3149), .A(w3147), .B(w3008), .C(w3148) );
	vdp_not g3640 (.nZ(w3129), .A(w3149) );
	vdp_nand3 g3641 (.Z(w3216), .A(w3148), .B(w3147), .C(w3156) );
	vdp_not g3642 (.nZ(w3119), .A(w3216) );
	vdp_not g3643 (.nZ(w3266), .A(w3262) );
	vdp_not g3644 (.nZ(w3265), .A(w3263) );
	vdp_not g3645 (.nZ(w3892), .A(w3267) );
	vdp_not g3646 (.nZ(w3264), .A(M5) );
	vdp_not g3647 (.nZ(w3919), .A(PLANE_A_PRIO) );
	vdp_not g3648 (.nZ(w3899), .A(PLANE_B_PRIO) );
	vdp_bufif0 g3649 (.Z(COL[5]), .A(w3097), .nE(w3899) );
	vdp_bufif0 g3650 (.Z(COL[6]), .A(w3178), .nE(w3899) );
	vdp_bufif0 g3651 (.Z(COL[4]), .A(w3099), .nE(w3899) );
	vdp_bufif0 g3652 (.Z(COL[3]), .A(w3100), .nE(w3899) );
	vdp_bufif0 g3653 (.Z(COL[2]), .A(w3095), .nE(w3899) );
	vdp_bufif0 g3654 (.Z(COL[1]), .A(w3109), .nE(w3899) );
	vdp_bufif0 g3655 (.Z(COL[0]), .A(w3098), .nE(w3899) );
	vdp_bufif0 g3656 (.Z(COL[5]), .A(w3302), .nE(w3919) );
	vdp_bufif0 g3657 (.Z(COL[6]), .A(w3397), .nE(w3919) );
	vdp_bufif0 g3658 (.Z(COL[4]), .A(w3301), .nE(w3919) );
	vdp_bufif0 g3659 (.Z(COL[3]), .A(w3303), .nE(w3919) );
	vdp_bufif0 g3660 (.Z(COL[2]), .A(w3268), .nE(w3919) );
	vdp_bufif0 g3661 (.Z(COL[1]), .A(w3918), .nE(w3919) );
	vdp_bufif0 g3662 (.Z(COL[0]), .A(w3328), .nE(w3919) );
	vdp_nand g3663 (.Z(w3012), .B(HCLK1), .A(w3006) );
	vdp_nand g3664 (.Z(w3018), .B(HCLK1), .A(w3005) );
	vdp_nand g3665 (.Z(w2973), .A(w3507), .B(HCLK1) );
	vdp_nand g3666 (.Z(w2924), .A(w3914), .B(HCLK1) );
	vdp_nor g3667 (.Z(w3915), .A(w3309), .B(w3366) );
	vdp_nand g3668 (.Z(w3021), .A(w3991), .B(HCLK1) );
	vdp_nand g3669 (.Z(w3263), .A(M5), .B(w3267) );
	vdp_nand g3670 (.Z(w3262), .A(M5), .B(w3892) );
	vdp_xor g3671 (.Z(w3427), .A(w3426), .B(w3425) );
	vdp_aon22 g3672 (.Z(w3425), .A1(w3423), .B1(w3502), .A2(VPOS[3]), .B2(w3424) );
	vdp_xnor g3673 (.Z(w3429), .A(w3426), .B(w3503) );
	vdp_aon22 g3674 (.Z(w3503), .A1(w3423), .B1(w3502), .A2(VPOS[2]), .B2(w3428) );
	vdp_xnor g3675 (.Z(w3431), .A(w3426), .B(w3501) );
	vdp_aon22 g3676 (.Z(w3501), .A1(w3423), .B1(w3502), .A2(VPOS[1]), .B2(w3430) );
	vdp_notif0 g3677 (.nZ(VRAMA[4]), .A(w3429), .nE(w3480) );
	vdp_notif0 g3678 (.nZ(VRAMA[3]), .A(w3431), .nE(w3480) );
	vdp_xnor g3679 (.Z(w3499), .A(w3426), .B(w3500) );
	vdp_aon22 g3680 (.Z(w3500), .A1(w3423), .B1(w3502), .A2(VPOS[0]), .B2(w3432) );
	vdp_notif0 g3681 (.nZ(VRAMA[2]), .A(w3499), .nE(w3480) );
	vdp_notif0 g3682 (.nZ(VRAMA[1]), .A(w3498), .nE(w3480) );
	vdp_notif0 g3683 (.nZ(VRAMA[0]), .A(1'b1), .nE(w3480) );
	vdp_not g3684 (.nZ(w3495), .A(w3506) );
	vdp_not g3685 (.nZ(w3480), .A(w3505) );
	vdp_comp_we g3686 (.Z(w3423), .nZ(w3502), .A(w3985) );
	vdp_comp_we g3687 (.Z(w3433), .nZ(w3497), .A(w1) );
	vdp_notif0 g3688 (.nZ(VRAMA[5]), .A(w3435), .nE(w3495) );
	vdp_aoi22 g3689 (.Z(w3435), .A1(w3427), .B1(w3434), .A2(w3433), .B2(w3497) );
	vdp_notif0 g3690 (.nZ(VRAMA[6]), .A(w3436), .nE(w3495) );
	vdp_aoi22 g3691 (.Z(w3436), .A1(w3434), .B1(w3437), .A2(w3433), .B2(w3497) );
	vdp_notif0 g3692 (.nZ(VRAMA[7]), .A(w3438), .nE(w3495) );
	vdp_aoi22 g3693 (.Z(w3438), .A1(w3437), .B1(w3439), .A2(w3433), .B2(w3497) );
	vdp_notif0 g3694 (.nZ(VRAMA[8]), .A(w3440), .nE(w3495) );
	vdp_aoi22 g3695 (.Z(w3440), .A1(w3439), .B1(w3441), .A2(w3433), .B2(w3497) );
	vdp_notif0 g3696 (.nZ(VRAMA[9]), .A(w3922), .nE(w3495) );
	vdp_aoi22 g3697 (.Z(w3922), .A1(w3441), .B1(w3443), .A2(w3433), .B2(w3497) );
	vdp_notif0 g3698 (.nZ(VRAMA[10]), .A(w3442), .nE(w3495) );
	vdp_aoi22 g3699 (.Z(w3442), .A1(w3443), .B1(w3444), .A2(w3433), .B2(w3497) );
	vdp_notif0 g3700 (.nZ(VRAMA[11]), .A(w3921), .nE(w3495) );
	vdp_aoi22 g3701 (.Z(w3921), .A1(w3444), .B1(w3446), .A2(w3433), .B2(w3497) );
	vdp_notif0 g3702 (.nZ(VRAMA[12]), .A(w3447), .nE(w3495) );
	vdp_aoi22 g3703 (.Z(w3447), .A1(w3446), .B1(w3445), .A2(w3433), .B2(w3497) );
	vdp_notif0 g3704 (.nZ(VRAMA[13]), .A(w3449), .nE(w3495) );
	vdp_aoi22 g3705 (.Z(w3449), .A1(w3445), .B1(w3448), .A2(w3433), .B2(w3497) );
	vdp_not g3706 (.nZ(w3496), .A(w3942) );
	vdp_notif0 g3707 (.nZ(VRAMA[14]), .A(w3451), .nE(w3496) );
	vdp_aoi22 g3708 (.Z(w3451), .A1(w3448), .B1(w3450), .A2(w3433), .B2(w3497) );
	vdp_notif0 g3709 (.nZ(VRAMA[15]), .A(w3453), .nE(w3496) );
	vdp_aoi22 g3710 (.Z(w3453), .A1(w3450), .B1(w3452), .A2(w3433), .B2(w3497) );
	vdp_notif0 g3711 (.nZ(VRAMA[16]), .A(w3455), .nE(w3496) );
	vdp_aoi22 g3712 (.Z(w3455), .A1(w3452), .B1(w3454), .A2(w3433), .B2(w3497) );
	vdp_notif0 g3713 (.nZ(VRAMA[5]), .A(w3458), .nE(w3494) );
	vdp_aoi22 g3714 (.Z(w3458), .A1(w3456), .B1(w3427), .A2(w3457), .B2(w3493) );
	vdp_notif0 g3715 (.nZ(VRAMA[6]), .A(w3460), .nE(w3494) );
	vdp_aoi22 g3716 (.Z(w3460), .A1(w3456), .B1(w3457), .A2(w3459), .B2(w3493) );
	vdp_notif0 g3717 (.nZ(VRAMA[7]), .A(w3461), .nE(w3494) );
	vdp_aoi22 g3718 (.Z(w3461), .A1(w3456), .B1(w3459), .A2(w3479), .B2(w3493) );
	vdp_notif0 g3719 (.nZ(VRAMA[8]), .A(w3462), .nE(w3494) );
	vdp_aoi22 g3720 (.Z(w3462), .A1(w3456), .B1(w3479), .A2(w3463), .B2(w3493) );
	vdp_notif0 g3721 (.nZ(VRAMA[9]), .A(w3464), .nE(w3494) );
	vdp_aoi22 g3722 (.Z(w3464), .A1(w3456), .B1(w3463), .A2(w3465), .B2(w3493) );
	vdp_notif0 g3723 (.nZ(VRAMA[10]), .A(w3467), .nE(w3494) );
	vdp_aoi22 g3724 (.Z(w3467), .A1(w3456), .B1(w3465), .A2(w3466), .B2(w3493) );
	vdp_notif0 g3725 (.nZ(VRAMA[11]), .A(w3469), .nE(w3492) );
	vdp_aoi22 g3726 (.Z(w3469), .A1(w3456), .B1(w3466), .A2(w3468), .B2(w3493) );
	vdp_notif0 g3727 (.nZ(VRAMA[12]), .A(w3471), .nE(w3492) );
	vdp_aoi22 g3728 (.Z(w3471), .A1(w3456), .B1(w3468), .A2(w3470), .B2(w3493) );
	vdp_notif0 g3729 (.nZ(VRAMA[14]), .A(w3474), .nE(w3492) );
	vdp_aoi22 g3730 (.Z(w3474), .A1(w3456), .B1(w3472), .A2(w3475), .B2(w3493) );
	vdp_notif0 g3731 (.nZ(VRAMA[15]), .A(w3477), .nE(w3492) );
	vdp_aoi22 g3732 (.Z(w3477), .A1(w3456), .B1(w3475), .A2(w3476), .B2(w3493) );
	vdp_notif0 g3733 (.nZ(VRAMA[16]), .A(w3478), .nE(w3492) );
	vdp_aoi22 g3734 (.Z(w3478), .A1(w3456), .B1(w3476), .A2(w3454), .B2(w3493) );
	vdp_notif0 g3735 (.nZ(VRAMA[13]), .A(w3473), .nE(w3492) );
	vdp_aoi22 g3736 (.Z(w3473), .A1(w3456), .B1(w3470), .A2(w3472), .B2(w3493) );
	vdp_not g3737 (.nZ(w3494), .A(w3422) );
	vdp_comp_we g3738 (.Z(w3493), .nZ(w3456), .A(w1) );
	vdp_aon22 g3739 (.Z(w3454), .A1(w3417), .B1(w3416), .A2(w3418), .B2(w3489) );
	vdp_not g3740 (.nZ(w3492), .A(w3422) );
	vdp_not g3741 (.nZ(w3418), .A(w3489) );
	vdp_sr_bit g3742 (.Q(w3505), .D(w3520), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3743 (.Q(w3489), .D(HPOS[3]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3744 (.Q(w3498), .D(w3556), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3745 (.Q(w3506), .D(w3993), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3746 (.Q(w3504), .D(w3984), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3747 (.Q(w3524), .D(w3983), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3748 (.Q(w3491), .D(w3982), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3749 (.Q(w3958), .D(w3959), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3750 (.Q(w3960), .D(w3958), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3751 (.Q(w3507), .D(w3960), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3752 (.Q(w3538), .D(w97), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3753 (.Q(w3517), .D(w35), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3754 (.Q(w3961), .D(w36), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3755 (.Q(w3578), .D(w3961), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3756 (.Q(w3579), .D(w3517), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3757 (.Q(w3576), .D(w3538), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3758 (.Q(w3580), .D(w3490), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3759 (.Q(w3581), .D(w3066), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3760 (.Q(w3582), .D(w3067), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3761 (.Q(w3583), .D(w3065), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3762 (.Q(w3611), .D(w3064), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3763 (.Q(w3612), .D(w3063), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3764 (.Q(w3515), .D(w3513), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3765 (.Q(w3516), .D(w3515), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3766 (.Q(w3962), .D(w3516), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_aon22 g3767 (.Z(w3529), .A1(H40), .B1(HPOS[8]), .A2(w3527), .B2(w3526) );
	vdp_aon22 g3768 (.Z(w3608), .A1(w3509), .B1(HPOS[8]), .A2(w3529), .B2(w3519) );
	vdp_aon22 g3769 (.Z(w3571), .A1(w3514), .B1(w3527), .A2(w3529), .B2(w3519) );
	vdp_or3 g3770 (.Z(w3577), .A(w3538), .B(w3517), .C(w3961) );
	vdp_or g3771 (.Z(w3530), .A(M5), .B(w3356) );
	vdp_bufif0 g3772 (.Z(VRAMA[1]), .A(w3957), .nE(w3518) );
	vdp_or g3773 (.Z(w3604), .A(w3529), .B(HPOS[4]) );
	vdp_bufif0 g3774 (.Z(VRAMA[2]), .A(w3532), .nE(w3518) );
	vdp_or g3775 (.Z(w3605), .A(w3529), .B(HPOS[5]) );
	vdp_bufif0 g3776 (.Z(VRAMA[3]), .A(w3533), .nE(w3518) );
	vdp_or g3777 (.Z(w3609), .A(w3529), .B(HPOS[6]) );
	vdp_bufif0 g3778 (.Z(VRAMA[4]), .A(w3534), .nE(w3518) );
	vdp_or g3779 (.Z(w3607), .A(w3529), .B(HPOS[7]) );
	vdp_bufif0 g3780 (.Z(VRAMA[5]), .A(w3535), .nE(w3518) );
	vdp_bufif0 g3781 (.Z(VRAMA[5]), .A(w3508), .nE(w3518) );
	vdp_not g3782 (.nZ(w3523), .A(w3415) );
	vdp_not g3783 (.nZ(w3963), .A(HPOS[3]) );
	vdp_dlatch_inv g3784 (.nQ(w3513), .D(w3512), .C(DCLK1), .nC(nDCLK1) );
	vdp_not g3785 (.nZ(w3527), .A(w3941) );
	vdp_not g3786 (.nZ(w3519), .A(w3529) );
	vdp_not g3787 (.nZ(w3526), .A(H40) );
	vdp_not g3788 (.nZ(w3518), .A(w3525) );
	vdp_bufif0 g3789 (.Z(VRAMA[0]), .A(1'b0), .nE(w3518) );
	vdp_or g3790 (.Z(w3525), .A(w3504), .B(w3524) );
	vdp_or g3791 (.Z(w3959), .A(w3522), .B(w6) );
	vdp_nand3 g3792 (.Z(w3575), .A(M5), .B(w3523), .C(HPOS[3]) );
	vdp_nand3 g3793 (.Z(w3536), .A(M5), .B(w3523), .C(w3963) );
	vdp_and g3794 (.Z(w3537), .A(DCLK2), .B(w3962) );
	vdp_and g3795 (.Z(w3511), .A(w3516), .B(DCLK2) );
	vdp_and g3796 (.Z(w3574), .A(w3515), .B(DCLK2) );
	vdp_and g3797 (.Z(w3510), .A(w3513), .B(DCLK2) );
	vdp_and g3798 (.Z(w3942), .A(M5), .B(w3506) );
	vdp_and g3799 (.Z(w3564), .A(HPOS[3]), .B(w3528) );
	vdp_and g3800 (.Z(w3982), .A(w3415), .B(w6) );
	vdp_and g3801 (.Z(w3983), .A(w3523), .B(w6) );
	vdp_and3 g3802 (.Z(w3984), .A(w3522), .B(M5), .C(w3521) );
	vdp_nor g3803 (.Z(w3528), .A(M5), .B(w3529) );
	vdp_nand g3804 (.Z(w3512), .A(w3175), .B(HCLK1) );
	vdp_oai21 g3805 (.A1(HPOS[6]), .A2(HPOS[7]), .B(HPOS[8]), .Z(w3941) );
	vdp_slatch g3806 (.Q(w3553), .D(REG_BUS[0]), .C(w3599), .nC(w3598) );
	vdp_slatch g3807 (.Q(w3549), .D(S[0]), .C(w3594), .nC(w3593) );
	vdp_slatch g3808 (.Q(w3550), .D(S[0]), .C(w3595), .nC(w3592) );
	vdp_slatch g3809 (.Q(w3551), .D(REG_BUS[1]), .C(w3599), .nC(w3598) );
	vdp_slatch g3810 (.Q(w3547), .D(S[1]), .C(w3594), .nC(w3593) );
	vdp_slatch g3811 (.Q(w3620), .D(S[1]), .C(w3595), .nC(w3592) );
	vdp_slatch g3812 (.Q(w3621), .D(REG_BUS[2]), .C(w3599), .nC(w3598) );
	vdp_slatch g3813 (.Q(w3541), .D(S[2]), .C(w3594), .nC(w3593) );
	vdp_slatch g3814 (.Q(w3622), .D(S[2]), .C(w3595), .nC(w3592) );
	vdp_slatch g3815 (.Q(w3618), .D(REG_BUS[3]), .C(w3599), .nC(w3598) );
	vdp_slatch g3816 (.Q(w3617), .D(S[3]), .C(w3594), .nC(w3593) );
	vdp_slatch g3817 (.Q(w4280), .D(S[3]), .C(w3595), .nC(w3592) );
	vdp_slatch g3818 (.Q(w3563), .D(REG_BUS[4]), .C(w3599), .nC(w3598) );
	vdp_slatch g3819 (.Q(w3616), .D(S[4]), .C(w3594), .nC(w3593) );
	vdp_slatch g3820 (.Q(w3615), .D(S[4]), .C(w3595), .nC(w3592) );
	vdp_slatch g3821 (.Q(w3614), .D(REG_BUS[5]), .C(w3599), .nC(w3598) );
	vdp_slatch g3822 (.Q(w3602), .D(S[5]), .C(w3594), .nC(w3593) );
	vdp_slatch g3823 (.Q(w3601), .D(S[5]), .C(w3595), .nC(w3592) );
	vdp_slatch g3824 (.Q(w3600), .D(REG_BUS[6]), .C(w3599), .nC(w3598) );
	vdp_slatch g3825 (.Q(w3596), .D(S[6]), .C(w3594), .nC(w3593) );
	vdp_slatch g3826 (.Q(w3597), .D(S[6]), .C(w3595), .nC(w3592) );
	vdp_slatch g3827 (.Q(w3591), .D(REG_BUS[7]), .C(w3599), .nC(w3598) );
	vdp_slatch g3828 (.Q(w3590), .D(S[7]), .C(w3594), .nC(w3593) );
	vdp_slatch g3829 (.Q(w3589), .D(S[7]), .C(w3595), .nC(w3592) );
	vdp_slatch g3830 (.Q(w3587), .D(S[0]), .C(w3567), .nC(w3584) );
	vdp_slatch g3831 (.Q(w3569), .D(S[0]), .C(w3568), .nC(w3588) );
	vdp_slatch g3832 (.Q(w3573), .D(S[1]), .C(w3568), .nC(w3588) );
	vdp_slatch g3833 (.Q(w3572), .D(S[1]), .C(w3567), .nC(w3584) );
	vdp_slatch g3834 (.Q(w3565), .D(w3591), .C(w3546), .nC(w3545) );
	vdp_slatch g3835 (.Q(w3559), .D(w3600), .C(w3546), .nC(w3545) );
	vdp_slatch g3836 (.Q(w3562), .D(w3614), .C(w3546), .nC(w3545) );
	vdp_slatch g3837 (.Q(w3624), .D(w3563), .C(w3546), .nC(w3545) );
	vdp_slatch g3838 (.Q(w3539), .D(w3618), .C(w3546), .nC(w3545) );
	vdp_slatch g3839 (.Q(w3540), .D(w3621), .C(w3546), .nC(w3545) );
	vdp_slatch g3840 (.Q(w3548), .D(w3551), .C(w3546), .nC(w3545) );
	vdp_slatch g3841 (.Q(w3552), .D(w3553), .C(w3546), .nC(w3545) );
	vdp_fa g3842 (.CI(w3939), .SUM(w3888), .B(w3571), .A(w3586) );
	vdp_fa g3843 (.CO(w3939), .CI(w3570), .SUM(w3764), .B(w3608), .A(w3613) );
	vdp_fa g3844 (.CO(w3613), .CI(w3566), .SUM(w3535), .B(w3607), .A(w3938) );
	vdp_fa g3845 (.CO(w3938), .CI(w3560), .SUM(w3534), .B(w3609), .A(w3610) );
	vdp_fa g3846 (.CO(w3610), .CI(w3561), .SUM(w3533), .B(w3605), .A(w3606) );
	vdp_fa g3847 (.CO(w3606), .CI(w3663), .SUM(w3532), .B(w3604), .A(w3603) );
	vdp_fa g3848 (.CO(w3603), .CI(w3530), .SUM(w3957), .B(w3564), .A(1'b1) );
	vdp_aon222 g3849 (.A1(w3543), .B1(w3531), .C1(w3542), .A2(w3572), .B2(w3573), .C2(1'b0), .Z(w3586) );
	vdp_aon222 g3850 (.A1(w3543), .B1(w3531), .C1(w3542), .A2(w3587), .B2(w3569), .C2(1'b0), .Z(w3570) );
	vdp_aon222 g3851 (.A1(w3543), .B1(w3531), .C1(w3542), .A2(w3589), .B2(w3590), .C2(w3565), .Z(w3566) );
	vdp_aon222 g3852 (.A1(w3543), .B1(w3531), .C1(w3542), .A2(w3597), .B2(w3596), .C2(w3559), .Z(w3560) );
	vdp_aon222 g3853 (.A1(w3543), .B1(w3531), .C1(w3542), .A2(w3601), .B2(w3602), .C2(w3562), .Z(w3561) );
	vdp_aon222 g3854 (.A1(w3543), .B1(w3531), .C1(w3542), .A2(w3615), .B2(w3616), .C2(w3624), .Z(w3663) );
	vdp_aon222 g3855 (.A1(w3543), .B1(w3531), .C1(w3542), .A2(w4280), .B2(w3617), .C2(w3539), .Z(w3356) );
	vdp_aon222 g3856 (.A1(w3543), .B1(w3531), .C1(w3542), .A2(w3622), .B2(w3541), .C2(w3540), .Z(w3052) );
	vdp_aon222 g3857 (.A1(w3543), .B1(w3531), .A2(w3620), .B2(w3547), .C2(w3548), .Z(w3354), .C1(w3542) );
	vdp_aon222 g3858 (.A1(w3543), .B1(w3531), .C1(w3542), .A2(w3550), .B2(w3549), .C2(w3552), .Z(w3352) );
	vdp_comp_strong g3859 (.Z(w3567), .nZ(w3584), .A(w3537) );
	vdp_comp_strong g3860 (.Z(w3568), .nZ(w3588), .A(w3574) );
	vdp_not g3861 (.nZ(w3531), .A(w3536) );
	vdp_not g3862 (.nZ(w3543), .A(w3575) );
	vdp_not g3863 (.nZ(w3542), .A(w3619) );
	vdp_not g3864 (.nZ(w3554), .A(w84) );
	vdp_not g3865 (.nZ(w3521), .A(w92) );
	vdp_not g3866 (.nZ(w3555), .A(w3556) );
	vdp_not g3867 (.nZ(w3522), .A(w3557) );
	vdp_not g3868 (.nZ(w3558), .A(M5) );
	vdp_comp_strong g3869 (.Z(w3594), .nZ(w3593), .A(w3510) );
	vdp_comp_strong g3870 (.Z(w3595), .nZ(w3592), .A(w3511) );
	vdp_comp_strong g3871 (.Z(w3599), .nZ(w3598), .A(w170) );
	vdp_comp_strong g3872 (.Z(w3546), .nZ(w3545), .A(w3623) );
	vdp_or g3873 (.Z(w3619), .A(w3943), .B(M5) );
	vdp_or g3874 (.Z(w3993), .A(w12), .B(w3555) );
	vdp_or g3875 (.Z(w3520), .A(w12), .B(w13) );
	vdp_or g3876 (.Z(w3623), .A(w4), .B(w91) );
	vdp_or5 g3877 (.E(w3554), .C(VPOS[6]), .D(VPOS[5]), .Z(w3943), .A(VPOS[7]), .B(VPOS[4]) );
	vdp_aoi21 g3878 (.Z(w3557), .A1(w92), .A2(w3003), .B(w7) );
	vdp_nand g3879 (.Z(w3556), .A(w13), .B(w3558) );
	vdp_slatch g3880 (.Q(w3658), .D(w4271), .C(w3627), .nC(w3628) );
	vdp_slatch g3881 (.Q(w3633), .D(w4272), .C(w3627), .nC(w3628) );
	vdp_slatch g3882 (.Q(w3634), .D(w4273), .C(w3627), .nC(w3628) );
	vdp_slatch g3883 (.Q(w3635), .D(w4270), .C(w3627), .nC(w3628) );
	vdp_slatch g3884 (.Q(w3637), .D(w4269), .C(w3627), .nC(w3628) );
	vdp_slatch g3885 (.Q(w3636), .D(w4268), .C(w3627), .nC(w3628) );
	vdp_slatch g3886 (.nQ(w3642), .D(w4276), .C(w3629), .nC(w3630) );
	vdp_slatch g3887 (.Q(w3653), .D(w4277), .C(w3629), .nC(w3630) );
	vdp_slatch g3888 (.Q(w3641), .D(w4278), .C(w3629), .nC(w3630) );
	vdp_slatch g3889 (.Q(w3640), .D(w4279), .C(w3629), .nC(w3630) );
	vdp_slatch g3890 (.Q(w3639), .D(w4275), .C(w3629), .nC(w3630) );
	vdp_slatch g3891 (.Q(w3638), .D(w4274), .C(w3629), .nC(w3630) );
	vdp_comp_strong g3892 (.Z(w3627), .nZ(w3628), .A(w3647) );
	vdp_comp_strong g3893 (.Z(w3629), .nZ(w3630), .A(w3964) );
	vdp_cgi2a g3894 (.Z(w3887), .A(w3638), .B(HPOS[4]), .C(1'b1) );
	vdp_cgi2a g3895 (.Z(w3882), .A(w3639), .B(HPOS[5]), .C(w3887) );
	vdp_cgi2a g3896 (.Z(w3881), .A(w3640), .B(HPOS[6]), .C(w3882) );
	vdp_cgi2a g3897 (.Z(w3883), .A(w3641), .B(HPOS[7]), .C(w3881) );
	vdp_cgi2a g3898 (.Z(w3643), .A(w3653), .B(HPOS[8]), .C(w3883) );
	vdp_cgi2a g3899 (.Z(w3648), .A(w3645), .B(w3633), .C(w3966) );
	vdp_cgi2a g3900 (.Z(w3966), .A(w3646), .B(w3634), .C(w3884) );
	vdp_cgi2a g3901 (.Z(w3884), .A(w3649), .B(w3635), .C(w3885) );
	vdp_cgi2a g3902 (.Z(w3885), .A(w3652), .B(w3637), .C(w3886) );
	vdp_cgi2a g3903 (.Z(w3886), .A(w3651), .B(w3636), .C(1'b0) );
	vdp_slatch g3904 (.Q(w4271), .D(REG_BUS[7]), .C(w3655), .nC(w3632) );
	vdp_slatch g3905 (.Q(w4272), .D(REG_BUS[4]), .C(w3655), .nC(w3632) );
	vdp_slatch g3906 (.Q(w4273), .D(REG_BUS[3]), .C(w3655), .nC(w3632) );
	vdp_slatch g3907 (.Q(w4270), .D(REG_BUS[2]), .C(w3655), .nC(w3632) );
	vdp_slatch g3908 (.Q(w4269), .D(REG_BUS[1]), .C(w3655), .nC(w3632) );
	vdp_slatch g3909 (.Q(w4268), .D(REG_BUS[0]), .C(w3655), .nC(w3632) );
	vdp_comp_strong g3910 (.Z(w3655), .nZ(w3632), .A(w162) );
	vdp_slatch g3911 (.Q(w4276), .D(REG_BUS[7]), .C(w3656), .nC(w3654) );
	vdp_slatch g3912 (.Q(w4277), .D(REG_BUS[4]), .C(w3656), .nC(w3654) );
	vdp_slatch g3913 (.Q(w4278), .D(REG_BUS[3]), .C(w3656), .nC(w3654) );
	vdp_slatch g3914 (.Q(w4279), .D(REG_BUS[2]), .C(w3656), .nC(w3654) );
	vdp_slatch g3915 (.Q(w4275), .D(REG_BUS[1]), .C(w3656), .nC(w3654) );
	vdp_slatch g3916 (.Q(w4274), .D(REG_BUS[0]), .C(w3656), .nC(w3654) );
	vdp_comp_strong g3917 (.Z(w3656), .nZ(w3654), .A(w161) );
	vdp_xor g3918 (.Z(w3657), .A(w3658), .B(w3648) );
	vdp_xor g3919 (.Z(w3644), .A(w3642), .B(w3643) );
	vdp_aon22 g3920 (.Z(w3645), .A1(w3650), .B1(w3661), .A2(VPOS[8]), .B2(VPOS[7]) );
	vdp_aon22 g3921 (.Z(w3646), .A1(w3650), .B1(w3661), .A2(VPOS[7]), .B2(VPOS[6]) );
	vdp_aon22 g3922 (.Z(w3649), .A1(w3650), .B1(w3661), .A2(VPOS[6]), .B2(VPOS[5]) );
	vdp_aon22 g3923 (.Z(w3652), .A1(w3650), .B1(w3661), .A2(VPOS[5]), .B2(VPOS[4]) );
	vdp_aon22 g3924 (.Z(w3651), .A1(w3650), .B1(w3661), .A2(VPOS[4]), .B2(VPOS[3]) );
	vdp_aon22 g3925 (.Z(w3668), .A1(w3650), .B1(w3661), .A2(VPOS[3]), .B2(VPOS[2]) );
	vdp_aon22 g3926 (.Z(w3667), .A1(w3650), .B1(w3661), .A2(VPOS[2]), .B2(VPOS[1]) );
	vdp_aon22 g3927 (.Z(w3666), .A1(w3650), .B1(w3661), .A2(VPOS[1]), .B2(VPOS[0]) );
	vdp_comp_we g3928 (.Z(w3650), .nZ(w3661), .A(w1) );
	vdp_not g3929 (.nZ(w3415), .A(w3965) );
	vdp_not g3930 (.nZ(w3660), .A(HPOS[3]) );
	vdp_not g3931 (.nZ(w3968), .A(w3967) );
	vdp_or g3932 (.Z(w3964), .A(w91), .B(w4) );
	vdp_or g3933 (.Z(w3647), .A(w91), .B(w3968) );
	vdp_oai21 g3934 (.Z(w3967), .A1(w5), .A2(M5), .B(w4) );
	vdp_and g3935 (.Z(w3659), .A(w3644), .B(w3662) );
	vdp_oai211 g3936 (.Z(w3965), .A1(w3660), .A2(M5), .B(w3659), .C(w3657) );
	vdp_slatch g3937 (.nQ(w3701), .D(REG_BUS[4]), .C(w3673), .nC(w3674) );
	vdp_slatch g3938 (.nQ(w3703), .D(REG_BUS[4]), .C(w3671), .nC(w3672) );
	vdp_slatch g3939 (.nQ(w3702), .D(REG_BUS[5]), .C(w3673), .nC(w3674) );
	vdp_slatch g3940 (.nQ(w3704), .D(REG_BUS[5]), .C(w3671), .nC(w3672) );
	vdp_slatch g3941 (.nQ(w3677), .D(REG_BUS[6]), .C(w3673), .nC(w3674) );
	vdp_slatch g3942 (.nQ(w3678), .D(REG_BUS[6]), .C(w3671), .nC(w3672) );
	vdp_slatch g3943 (.nQ(w4267), .D(REG_BUS[1]), .C(w3671), .nC(w3672) );
	vdp_slatch g3944 (.nQ(w3697), .D(REG_BUS[2]), .C(w3673), .nC(w3674) );
	vdp_slatch g3945 (.nQ(w3698), .D(REG_BUS[2]), .C(w3671), .nC(w3672) );
	vdp_slatch g3946 (.nQ(w3699), .D(REG_BUS[3]), .C(w3673), .nC(w3674) );
	vdp_slatch g3947 (.nQ(w3700), .D(REG_BUS[3]), .C(w3671), .nC(w3672) );
	vdp_slatch g3948 (.nQ(w3705), .D(REG_BUS[0]), .C(w3671), .nC(w3672) );
	vdp_slatch g3949 (.nQ(w3675), .D(REG_BUS[1]), .C(w3673), .nC(w3674) );
	vdp_slatch g3950 (.Q(w3417), .D(REG_BUS[0]), .C(w3664), .nC(w3665) );
	vdp_slatch g3951 (.Q(w3416), .D(REG_BUS[4]), .C(w3664), .nC(w3665) );
	vdp_not g3952 (.nZ(w3970), .A(w3675) );
	vdp_aoi22 g3953 (.Z(w3694), .A1(HPOS[8]), .B1(w3651), .A2(w3670), .B2(w3669) );
	vdp_aoi22 g3954 (.Z(w3695), .A1(w3651), .B1(w3652), .A2(w3670), .B2(w3669) );
	vdp_aoi22 g3955 (.Z(w3682), .A1(w3652), .B1(w3649), .A2(w3670), .B2(w3669) );
	vdp_aoi22 g3956 (.Z(w3707), .A1(w3646), .B1(w3645), .A2(w3670), .B2(w3669) );
	vdp_aoi22 g3957 (.Z(w3696), .A1(w3649), .B1(w3646), .A2(w3670), .B2(w3669) );
	vdp_comp_strong g3958 (.Z(w3664), .nZ(w3665), .A(w169) );
	vdp_comp_strong g3959 (.Z(w3673), .nZ(w3674), .A(w165) );
	vdp_comp_strong g3960 (.Z(w3671), .nZ(w3672), .A(w168) );
	vdp_aoi22 g3961 (.Z(w3706), .A1(w3645), .B1(w3669), .A2(w3670), .B2(w3970) );
	vdp_nand g3962 (.Z(w3708), .A(w3645), .B(HSCR) );
	vdp_nand g3963 (.Z(w3681), .A(w3646), .B(HSCR) );
	vdp_nand g3964 (.Z(w3709), .A(w3652), .B(HSCR) );
	vdp_nand g3965 (.Z(w3683), .A(w3649), .B(HSCR) );
	vdp_nand g3966 (.Z(w3693), .A(w3651), .B(HSCR) );
	vdp_nand g3967 (.Z(w3969), .A(w3668), .B(LSCR) );
	vdp_nand g3968 (.Z(w3994), .A(w3667), .B(LSCR) );
	vdp_nand g3969 (.Z(w3689), .A(w3666), .B(LSCR) );
	vdp_nand g3970 (.Z(w3662), .A(HPOS[7]), .B(HPOS[8]) );
	vdp_comp_we g3971 (.Z(w3670), .nZ(w3669), .A(H40) );
	vdp_notif0 g3972 (.nZ(VRAMA[16]), .A(w3678), .nE(w3676) );
	vdp_notif0 g3973 (.nZ(VRAMA[16]), .A(w3677), .nE(w3680) );
	vdp_notif0 g3974 (.nZ(VRAMA[15]), .A(w3704), .nE(w3676) );
	vdp_notif0 g3975 (.nZ(VRAMA[15]), .A(w3702), .nE(w3680) );
	vdp_notif0 g3976 (.nZ(VRAMA[14]), .A(w3703), .nE(w3676) );
	vdp_notif0 g3977 (.nZ(VRAMA[14]), .A(w3701), .nE(w3680) );
	vdp_notif0 g3978 (.nZ(VRAMA[13]), .A(w3700), .nE(w3676) );
	vdp_notif0 g3979 (.nZ(VRAMA[13]), .A(w3699), .nE(w3680) );
	vdp_notif0 g3980 (.nZ(VRAMA[12]), .A(w3698), .nE(w3676) );
	vdp_notif0 g3981 (.nZ(VRAMA[12]), .A(w3697), .nE(w3680) );
	vdp_notif0 g3982 (.nZ(VRAMA[11]), .A(w4267), .nE(w3676) );
	vdp_notif0 g3983 (.nZ(VRAMA[11]), .A(w3706), .nE(w3680) );
	vdp_notif0 g3984 (.nZ(VRAMA[10]), .A(w3705), .nE(w3676) );
	vdp_notif0 g3985 (.nZ(VRAMA[10]), .A(w3707), .nE(w3680) );
	vdp_notif0 g3986 (.nZ(VRAMA[9]), .A(w3708), .nE(w3679) );
	vdp_notif0 g3987 (.nZ(VRAMA[9]), .A(w3696), .nE(w3680) );
	vdp_notif0 g3988 (.nZ(VRAMA[6]), .A(w3709), .nE(w3679) );
	vdp_notif0 g3989 (.nZ(VRAMA[6]), .A(w3694), .nE(w3684) );
	vdp_notif0 g3990 (.nZ(VRAMA[5]), .A(w3693), .nE(w3679) );
	vdp_notif0 g3991 (.nZ(VRAMA[5]), .A(w3692), .nE(w3684) );
	vdp_notif0 g3992 (.nZ(VRAMA[4]), .A(w3969), .nE(w3679) );
	vdp_notif0 g3993 (.nZ(VRAMA[4]), .A(w3691), .nE(w3684) );
	vdp_notif0 g3994 (.nZ(VRAMA[3]), .A(w3994), .nE(w3679) );
	vdp_notif0 g3995 (.nZ(VRAMA[3]), .A(w3690), .nE(w3684) );
	vdp_notif0 g3996 (.nZ(VRAMA[2]), .A(w3689), .nE(w3679) );
	vdp_notif0 g3997 (.nZ(VRAMA[2]), .A(w3688), .nE(w3684) );
	vdp_notif0 g3998 (.nZ(VRAMA[1]), .A(1'b1), .nE(w3679) );
	vdp_notif0 g3999 (.nZ(VRAMA[1]), .A(1'b1), .nE(w3684) );
	vdp_notif0 g4000 (.nZ(VRAMA[0]), .A(w3686), .nE(w3679) );
	vdp_notif0 g4001 (.nZ(VRAMA[0]), .A(w3686), .nE(w3684) );
	vdp_notif0 g4002 (.nZ(VRAMA[8]), .A(w3681), .nE(w3679) );
	vdp_notif0 g4003 (.nZ(VRAMA[8]), .A(w3682), .nE(w3684) );
	vdp_notif0 g4004 (.nZ(VRAMA[7]), .A(w3683), .nE(w3679) );
	vdp_notif0 g4005 (.nZ(VRAMA[7]), .A(w3695), .nE(w3684) );
	vdp_not g4006 (.nZ(w3686), .A(1'b0) );
	vdp_not g4007 (.nZ(w3688), .A(HPOS[4]) );
	vdp_not g4008 (.nZ(w3690), .A(HPOS[5]) );
	vdp_not g4009 (.nZ(w3691), .A(HPOS[6]) );
	vdp_not g4010 (.nZ(w3692), .A(HPOS[7]) );
	vdp_not g4011 (.nZ(w3679), .A(w3174) );
	vdp_not g4012 (.nZ(w3676), .A(w3174) );
	vdp_not g4013 (.nZ(w3684), .A(w3491) );
	vdp_not g4014 (.nZ(w3680), .A(w3491) );
	vdp_not g4015 (.nZ(w3716), .A(w3880) );
	vdp_comp_strong g4016 (.Z(w3710), .nZ(w3711), .A(w166) );
	vdp_comp_we g4017 (.Z(w3715), .nZ(w3714), .A(w3504) );
	vdp_comp_strong g4018 (.Z(w3713), .nZ(w3712), .A(w164) );
	vdp_slatch g4019 (.Q(w3736), .D(REG_BUS[6]), .C(w3710), .nC(w3711) );
	vdp_slatch g4020 (.Q(w3979), .D(REG_BUS[3]), .C(w3713), .nC(w3712) );
	vdp_slatch g4021 (.Q(w3735), .D(REG_BUS[5]), .C(w3710), .nC(w3711) );
	vdp_slatch g4022 (.Q(w3733), .D(REG_BUS[2]), .C(w3713), .nC(w3712) );
	vdp_slatch g4023 (.Q(w3719), .D(REG_BUS[4]), .C(w3710), .nC(w3711) );
	vdp_slatch g4024 (.Q(w4281), .D(REG_BUS[1]), .C(w3713), .nC(w3712) );
	vdp_slatch g4025 (.Q(w3722), .D(REG_BUS[3]), .C(w3710), .nC(w3711) );
	vdp_slatch g4026 (.Q(w3980), .D(REG_BUS[0]), .C(w3713), .nC(w3712) );
	vdp_slatch g4027 (.Q(w3730), .D(REG_BUS[1]), .C(w3710), .nC(w3711) );
	vdp_slatch g4028 (.Q(w3727), .D(REG_BUS[2]), .C(w3710), .nC(w3711) );
	vdp_bufif0 g4029 (.Z(VRAMA[11]), .A(w3729), .nE(w3718) );
	vdp_bufif0 g4030 (.Z(VRAMA[10]), .A(w3723), .nE(w3718) );
	vdp_bufif0 g4031 (.Z(VRAMA[13]), .A(w3731), .nE(w3718) );
	vdp_bufif0 g4032 (.Z(VRAMA[9]), .A(w3721), .nE(w3718) );
	vdp_bufif0 g4033 (.Z(VRAMA[8]), .A(w3720), .nE(w3718) );
	vdp_bufif0 g4034 (.Z(VRAMA[14]), .A(w3732), .nE(w3716) );
	vdp_bufif0 g4035 (.Z(VRAMA[7]), .A(w3717), .nE(w3718) );
	vdp_bufif0 g4036 (.Z(VRAMA[15]), .A(w3940), .nE(w3716) );
	vdp_bufif0 g4037 (.Z(VRAMA[16]), .A(w3734), .nE(w3716) );
	vdp_aon22 g4038 (.Z(w3734), .A1(w3714), .B1(w3715), .A2(w3736), .B2(w3979) );
	vdp_aon22 g4039 (.Z(w3940), .A1(w3714), .B1(w3715), .A2(w3735), .B2(w3733) );
	vdp_aon22 g4040 (.Z(w3732), .A1(w3714), .B1(w3715), .A2(w3719), .B2(w4281) );
	vdp_aon22 g4041 (.Z(w3731), .A1(w3714), .B1(w3715), .A2(w3722), .B2(w3980) );
	vdp_aon22 g4042 (.Z(w3729), .A1(w3725), .B1(w3728), .A2(w3730), .B2(w3726) );
	vdp_aon22 g4043 (.Z(w3724), .A1(w3725), .B1(w3738), .A2(w3727), .B2(w3726) );
	vdp_bufif0 g4044 (.Z(VRAMA[12]), .A(w3724), .nE(w3718) );
	vdp_not g4045 (.nZ(w3718), .A(w3525) );
	vdp_and g4046 (.Z(w3880), .A(w3525), .B(M5) );
	vdp_comp_we g4047 (.Z(w3726), .nZ(w3725), .A(M5) );
	vdp_fa g4048 (.CO(w3753), .CI(w3929), .SUM(w3773), .B(VPOS[6]), .A(w3928) );
	vdp_fa g4049 (.CO(w3928), .CI(w3931), .SUM(w3754), .B(VPOS[5]), .A(w3930) );
	vdp_fa g4050 (.CO(w3930), .CI(w3933), .SUM(w3755), .B(VPOS[4]), .A(w3932) );
	vdp_fa g4051 (.CO(w3932), .CI(w3821), .SUM(w3424), .B(VPOS[3]), .A(w3934) );
	vdp_fa g4052 (.CO(w3934), .CI(w3936), .SUM(w3428), .B(VPOS[2]), .A(w3935) );
	vdp_fa g4053 (.CO(w3935), .CI(w3875), .SUM(w3430), .B(VPOS[1]), .A(w3937) );
	vdp_fa g4054 (.CO(w3937), .CI(w3834), .SUM(w3432), .B(VPOS[0]), .A(1'b0) );
	vdp_fa g4055 (.CO(w3772), .CI(w3927), .SUM(w3770), .B(VPOS[7]), .A(w3753) );
	vdp_fa g4056 (.CO(w3752), .CI(w3807), .SUM(w3781), .B(VPOS[8]), .A(w3772) );
	vdp_fa g4057 (.CO(w3780), .CI(w3808), .SUM(w3747), .B(1'b0), .A(w3752) );
	vdp_fa g4058 (.CI(w3792), .SUM(w3748), .B(1'b0), .A(w3780) );
	vdp_aon22 g4059 (.Z(w3792), .A1(w3790), .B1(w3791), .A2(w3751), .B2(w3750) );
	vdp_aon22 g4060 (.Z(w3808), .A1(w3878), .B1(w3795), .A2(w3751), .B2(w3750) );
	vdp_aon22 g4061 (.Z(w3807), .A1(w3796), .B1(w3797), .A2(w3751), .B2(w3750) );
	vdp_aon22 g4062 (.Z(w3927), .A1(w3799), .B1(w3800), .A2(w3751), .B2(w3750) );
	vdp_aon22 g4063 (.Z(w3929), .A1(w3806), .B1(w3803), .A2(w3751), .B2(w3750) );
	vdp_aon22 g4064 (.Z(w3931), .A1(w3811), .B1(w3810), .A2(w3751), .B2(w3750) );
	vdp_aon22 g4065 (.Z(w3933), .A1(w3815), .B1(w3816), .A2(w3751), .B2(w3750) );
	vdp_aon22 g4066 (.Z(w3821), .A1(w3820), .B1(w3819), .A2(w3751), .B2(w3750) );
	vdp_aon22 g4067 (.Z(w3936), .A1(w3822), .B1(w3823), .A2(w3751), .B2(w3750) );
	vdp_aon22 g4068 (.Z(w3875), .A1(w3826), .B1(w3879), .A2(w3751), .B2(w3750) );
	vdp_aon22 g4069 (.Z(w3834), .A1(w3828), .B1(w3827), .A2(w3751), .B2(w3750) );
	vdp_comp_we g4070 (.Z(w3751), .nZ(w3750), .A(w3759) );
	vdp_comp_strong g4071 (.Z(w3761), .nZ(w3756), .A(w167) );
	vdp_sr_bit g4072 (.Q(w3782), .D(RD_DATA[1]), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4073 (.Q(w3757), .D(RD_DATA[2]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4074 (.Q(w3831), .D(w3782), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4075 (.Q(w3845), .D(w3757), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4076 (.Q(w3830), .D(HPOS[3]), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4077 (.Q(w3509), .D(REG_BUS[0]), .C(w3761), .nC(w3756) );
	vdp_slatch g4078 (.Q(w3514), .D(REG_BUS[1]), .C(w3761), .nC(w3756) );
	vdp_slatch g4079 (.Q(w3777), .D(REG_BUS[5]), .C(w3761), .nC(w3756) );
	vdp_slatch g4080 (.Q(w3776), .D(REG_BUS[4]), .C(w3761), .nC(w3756) );
	vdp_slatch g4081 (.Q(w3828), .D(w3832), .C(w3783), .nC(w3787) );
	vdp_slatch g4082 (.Q(w3990), .D(w3833), .C(w3789), .nC(w3784) );
	vdp_slatch g4083 (.Q(w3826), .D(w3825), .C(w3783), .nC(w3787) );
	vdp_slatch g4084 (.Q(w3989), .D(w3824), .C(w3789), .nC(w3784) );
	vdp_slatch g4085 (.Q(w3822), .D(w3847), .C(w3783), .nC(w3787) );
	vdp_slatch g4086 (.Q(w3988), .D(w3818), .C(w3789), .nC(w3784) );
	vdp_slatch g4087 (.Q(w3820), .D(w3817), .C(w3783), .nC(w3787) );
	vdp_slatch g4088 (.Q(w3987), .D(w3814), .C(w3789), .nC(w3784) );
	vdp_slatch g4089 (.Q(w3815), .D(w3813), .C(w3783), .nC(w3787) );
	vdp_slatch g4090 (.Q(w3986), .D(w3812), .C(w3789), .nC(w3784) );
	vdp_slatch g4091 (.Q(w3811), .D(w3805), .C(w3783), .nC(w3787) );
	vdp_slatch g4092 (.Q(w3997), .D(w3804), .C(w3789), .nC(w3784) );
	vdp_slatch g4093 (.Q(w3806), .D(w3801), .C(w3783), .nC(w3787) );
	vdp_slatch g4094 (.Q(w3998), .D(w3802), .C(w3789), .nC(w3784) );
	vdp_slatch g4095 (.Q(w3799), .D(w3798), .C(w3783), .nC(w3787) );
	vdp_slatch g4096 (.Q(w3797), .D(w3809), .C(w3789), .nC(w3784) );
	vdp_slatch g4097 (.Q(w3796), .D(w3852), .C(w3783), .nC(w3787) );
	vdp_slatch g4098 (.Q(w3795), .D(w3794), .C(w3789), .nC(w3784) );
	vdp_slatch g4099 (.Q(w3878), .D(w3793), .C(w3783), .nC(w3787) );
	vdp_slatch g4100 (.Q(w3791), .D(w3867), .C(w3789), .nC(w3784) );
	vdp_slatch g4101 (.Q(w3790), .D(w3788), .C(w3783), .nC(w3787) );
	vdp_slatch g4102 (.Q(w3973), .D(REG_BUS[0]), .C(w3836), .nC(w3835) );
	vdp_aon22 g4103 (.Z(w3829), .A1(w3832), .B1(w3844), .A2(w3846), .B2(w3973) );
	vdp_slatch g4104 (.Q(w3848), .D(REG_BUS[1]), .C(w3836), .nC(w3835) );
	vdp_aon22 g4105 (.Z(w3833), .A1(w3825), .B1(w3844), .A2(w3846), .B2(w3848) );
	vdp_slatch g4106 (.Q(w3972), .D(REG_BUS[2]), .C(w3836), .nC(w3835) );
	vdp_aon22 g4107 (.Z(w3824), .A1(w3847), .B1(w3844), .A2(w3846), .B2(w3972) );
	vdp_slatch g4108 (.Q(w3849), .D(REG_BUS[3]), .C(w3836), .nC(w3835) );
	vdp_aon22 g4109 (.Z(w3818), .A1(w3817), .B1(w3844), .A2(w3846), .B2(w3849) );
	vdp_slatch g4110 (.Q(w3850), .D(REG_BUS[4]), .C(w3836), .nC(w3835) );
	vdp_aon22 g4111 (.Z(w3814), .A1(w3813), .B1(w3844), .A2(w3846), .B2(w3850) );
	vdp_slatch g4112 (.Q(w3876), .D(REG_BUS[5]), .C(w3836), .nC(w3835) );
	vdp_aon22 g4113 (.Z(w3812), .A1(w3805), .B1(w3844), .A2(w3846), .B2(w3876) );
	vdp_slatch g4114 (.Q(w3971), .D(REG_BUS[6]), .C(w3836), .nC(w3835) );
	vdp_aon22 g4115 (.Z(w3804), .A1(w3801), .B1(w3844), .A2(w3846), .B2(w3971) );
	vdp_slatch g4116 (.Q(w3851), .D(REG_BUS[7]), .C(w3836), .nC(w3835) );
	vdp_aon22 g4117 (.Z(w3802), .A1(w3798), .B1(w3844), .A2(w3846), .B2(w3851) );
	vdp_aon22 g4118 (.Z(w3809), .A1(w3852), .B1(w3844), .A2(w3846), .B2(1'b0) );
	vdp_aon22 g4119 (.Z(w3794), .A1(w3793), .B1(w3844), .A2(w3846), .B2(1'b0) );
	vdp_aon22 g4120 (.Z(w3867), .A1(w3788), .B1(w3844), .A2(w3846), .B2(1'b0) );
	vdp_notif0 g4121 (.nZ(RD_DATA[2]), .A(w3868), .nE(w3840) );
	vdp_slatch g4122 (.nQ(w3868), .D(w3788), .C(w3839), .nC(w3838) );
	vdp_notif0 g4123 (.nZ(RD_DATA[1]), .A(w3853), .nE(w3840) );
	vdp_slatch g4124 (.nQ(w3853), .D(w3793), .C(w3839), .nC(w3838) );
	vdp_notif0 g4125 (.nZ(RD_DATA[0]), .A(w3996), .nE(w3840) );
	vdp_slatch g4126 (.nQ(w3996), .D(w3852), .C(w3839), .nC(w3838) );
	vdp_notif0 g4127 (.nZ(AD_DATA[7]), .A(w4287), .nE(w3840) );
	vdp_slatch g4128 (.nQ(w4287), .D(w3798), .C(w3839), .nC(w3838) );
	vdp_notif0 g4129 (.nZ(AD_DATA[6]), .A(w3854), .nE(w3840) );
	vdp_slatch g4130 (.nQ(w3854), .D(w3801), .C(w3839), .nC(w3838) );
	vdp_notif0 g4131 (.nZ(AD_DATA[5]), .A(w3855), .nE(w3840) );
	vdp_slatch g4132 (.nQ(w3855), .D(w3805), .C(w3839), .nC(w3838) );
	vdp_notif0 g4133 (.nZ(AD_DATA[4]), .A(w3856), .nE(w3840) );
	vdp_slatch g4134 (.nQ(w3856), .D(w3813), .C(w3839), .nC(w3838) );
	vdp_notif0 g4135 (.nZ(AD_DATA[3]), .A(w3865), .nE(w3840) );
	vdp_slatch g4136 (.nQ(w3865), .D(w3817), .C(w3839), .nC(w3838) );
	vdp_notif0 g4137 (.nZ(AD_DATA[2]), .A(w3863), .nE(w3840) );
	vdp_slatch g4138 (.nQ(w3863), .D(w3847), .C(w3839), .nC(w3838) );
	vdp_notif0 g4139 (.nZ(AD_DATA[1]), .A(w3858), .nE(w3840) );
	vdp_slatch g4140 (.nQ(w3858), .D(w3825), .C(w3839), .nC(w3838) );
	vdp_notif0 g4141 (.nZ(AD_DATA[0]), .A(w3862), .nE(w3840) );
	vdp_slatch g4142 (.nQ(w3862), .D(w3832), .C(w3839), .nC(w3838) );
	vdp_sr_bit g4143 (.Q(w3861), .D(w3576), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4144 (.Q(w3869), .D(w3873), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4145 (.Q(w3873), .D(RD_DATA[0]), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4146 (.Q(w3995), .D(w3829), .C(w3789), .nC(w3784) );
	vdp_comp_strong g4147 (.Z(w3789), .nZ(w3784), .A(w3843) );
	vdp_comp_strong g4148 (.Z(w3783), .nZ(w3787), .A(w3841) );
	vdp_comp_strong g4149 (.Z(w3836), .nZ(w3835), .A(w171) );
	vdp_sr_bit g4150 (.Q(w3785), .D(w3976), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_comp_strong g4151 (.Z(w3839), .nZ(w3838), .A(w3860) );
	vdp_not g4152 (.nZ(w3840), .A(w3861) );
	vdp_and g4153 (.Z(w3860), .A(w3576), .B(HCLK1) );
	vdp_and g4154 (.Z(w3800), .A(w3998), .B(w3785) );
	vdp_and g4155 (.Z(w3803), .A(w3997), .B(w3785) );
	vdp_and g4156 (.Z(w3810), .A(w3986), .B(w3785) );
	vdp_and g4157 (.Z(w3816), .A(w3987), .B(w3785) );
	vdp_and g4158 (.Z(w3819), .A(w3988), .B(w3785) );
	vdp_and g4159 (.Z(w3823), .A(w3989), .B(w3785) );
	vdp_and g4160 (.Z(w3879), .A(w3990), .B(w3785) );
	vdp_and g4161 (.Z(w3827), .A(w3995), .B(w3785) );
	vdp_not g4162 (.nZ(w3975), .A(w3974) );
	vdp_not g4163 (.nZ(w3841), .A(w3842) );
	vdp_not g4164 (.nZ(w3759), .A(w3758) );
	vdp_not g4165 (.nZ(w3763), .A(w3509) );
	vdp_not g4166 (.nZ(w3762), .A(w3514) );
	vdp_not g4167 (.nZ(w3740), .A(w3977) );
	vdp_not g4168 (.nZ(w3739), .A(w3978) );
	vdp_not g4169 (.nZ(w3741), .A(w3981) );
	vdp_not g4170 (.nZ(w3926), .A(M5) );
	vdp_not g4171 (.nZ(w3779), .A(w3925) );
	vdp_aon22 g4172 (.Z(w3767), .A1(w3746), .B1(w3754), .A2(w3773), .B2(w3749) );
	vdp_aon22 g4173 (.Z(w3771), .A1(w3746), .B1(w3773), .A2(w3770), .B2(w3749) );
	vdp_ha g4174 (.CO(w3775), .SUM(w3745), .B(w3774), .A(w3771) );
	vdp_aon222 g4175 (.A1(w3741), .B1(w3739), .C1(w3740), .A2(w3769), .B2(w3768), .C2(w3745), .Z(w3721) );
	vdp_aon22 g4176 (.Z(w3924), .A1(w3746), .B1(w3770), .A2(w3781), .B2(w3749) );
	vdp_ha g4177 (.SUM(w3744), .B(w3775), .A(w3924) );
	vdp_aon222 g4178 (.A1(w3741), .B1(w3739), .C1(w3740), .A2(w3768), .B2(w3745), .C2(w3744), .Z(w3723) );
	vdp_ha g4179 (.CO(w3774), .SUM(w3768), .B(w3767), .A(w3778) );
	vdp_aon222 g4180 (.A1(w3741), .B1(w3739), .C1(w3740), .A2(w3765), .B2(w3769), .C2(w3768), .Z(w3720) );
	vdp_aon22 g4181 (.Z(w3769), .A1(w3746), .B1(w3755), .A2(w3754), .B2(w3749) );
	vdp_aon222 g4182 (.A1(w3741), .B1(w3739), .C1(w3740), .A2(w3888), .B2(w3765), .C2(w3769), .Z(w3717) );
	vdp_aon222 g4183 (.A1(w3741), .B1(w3739), .C1(w3740), .A2(w3764), .B2(w3764), .C2(w3765), .Z(w3508) );
	vdp_aon22 g4184 (.Z(w3765), .A1(w3746), .B1(w3424), .A2(w3755), .B2(w3749) );
	vdp_comp_we g4185 (.Z(w3846), .nZ(w3844), .A(M5) );
	vdp_comp_we g4186 (.Z(w3746), .nZ(w3749), .A(w1) );
	vdp_and g4187 (.Z(w3778), .A(w3779), .B(w3926) );
	vdp_aon222 g4188 (.A1(w3741), .B1(w3739), .C1(w3740), .A2(w3745), .B2(w3744), .C2(w3742), .Z(w3728) );
	vdp_aon222 g4189 (.A1(w3741), .B1(w3739), .C1(w3740), .A2(w3744), .B2(w3742), .C2(w3923), .Z(w3738) );
	vdp_aon22 g4190 (.Z(w3743), .A1(w3746), .B1(w3747), .A2(w3748), .B2(w3749) );
	vdp_aon22 g4191 (.Z(w3766), .A1(w3746), .B1(w3781), .A2(w3747), .B2(w3749) );
	vdp_and g4192 (.Z(w3742), .B(w3766), .A(w3776) );
	vdp_and g4193 (.Z(w3923), .B(w3743), .A(w3777) );
	vdp_oai21 g4194 (.Z(w3758), .A1(VSCR), .A2(w3830), .B(M5) );
	vdp_aoi21 g4195 (.Z(w3842), .A1(HCLK1), .A2(w15), .B(w91) );
	vdp_oai211 g4196 (.Z(w3974), .A1(HCLK1), .A2(w4), .B(w5), .C(M5) );
	vdp_or g4197 (.Z(w3843), .A(w91), .B(w3975) );
	vdp_nand3 g4198 (.Z(w3976), .A(w83), .B(HPOS[6]), .C(HPOS[7]) );
	vdp_nand g4199 (.Z(w3981), .A(w3514), .B(w3509) );
	vdp_nand g4200 (.Z(w3978), .A(w3509), .B(w3762) );
	vdp_nand g4201 (.Z(w3977), .A(w3762), .B(w3763) );
	vdp_aoi31 g4202 (.Z(w3925), .B3(w3924), .B2(w3771), .B1(w3767), .A(w3766) );
	vdp_slatch g4203 (.Q(w3457), .D(S[0]), .C(w3419), .nC(w3046) );
	vdp_slatch g4204 (.Q(w3459), .D(S[1]), .C(w3419), .nC(w3046) );
	vdp_slatch g4205 (.Q(w3479), .D(S[2]), .C(w3419), .nC(w3046) );
	vdp_slatch g4206 (.Q(w3463), .D(S[3]), .C(w3419), .nC(w3046) );
	vdp_slatch g4207 (.Q(w3465), .D(S[4]), .C(w3419), .nC(w3046) );
	vdp_slatch g4208 (.Q(w3466), .D(S[5]), .C(w3419), .nC(w3046) );
	vdp_slatch g4209 (.Q(w3468), .D(S[6]), .C(w3419), .nC(w3046) );
	vdp_slatch g4210 (.Q(w3470), .D(S[7]), .C(w3419), .nC(w3046) );
	vdp_slatch g4211 (.Q(w3472), .D(S[0]), .C(w3414), .nC(w3413) );
	vdp_slatch g4212 (.Q(w3475), .D(S[1]), .C(w3414), .nC(w3413) );
	vdp_slatch g4213 (.Q(w3476), .D(S[2]), .C(w3414), .nC(w3413) );
	vdp_slatch g4214 (.Q(w2993), .D(S[3]), .C(w3414), .nC(w3413) );
	vdp_slatch g4215 (.Q(w3483), .D(S[4]), .C(w3414), .nC(w3413) );
	vdp_slatch g4216 (.Q(w2970), .D(S[5]), .C(w3414), .nC(w3413) );
	vdp_slatch g4217 (.Q(w2972), .D(S[6]), .C(w3414), .nC(w3413) );
	vdp_slatch g4218 (.Q(w2998), .D(S[7]), .C(w3414), .nC(w3413) );
	vdp_comp_strong g4219 (.Z(w3414), .nZ(w3413), .A(w3181) );
	vdp_comp_strong g4220 (.Z(w3419), .nZ(w3046), .A(w3182) );
	vdp_comp_strong g4221 (.Z(w3420), .nZ(w3481), .A(w3183) );
	vdp_slatch g4222 (.Q(w3956), .D(S[7]), .C(w3420), .nC(w3481) );
	vdp_slatch g4223 (.Q(w3955), .D(S[6]), .C(w3420), .nC(w3481) );
	vdp_slatch g4224 (.Q(w3954), .D(S[5]), .C(w3420), .nC(w3481) );
	vdp_slatch g4225 (.Q(w3486), .D(S[4]), .C(w3420), .nC(w3481) );
	vdp_slatch g4226 (.Q(w3487), .D(S[3]), .C(w3420), .nC(w3481) );
	vdp_slatch g4227 (.Q(w3452), .D(S[2]), .C(w3420), .nC(w3481) );
	vdp_slatch g4228 (.Q(w3450), .D(S[1]), .C(w3420), .nC(w3481) );
	vdp_slatch g4229 (.Q(w3448), .D(S[0]), .C(w3420), .nC(w3481) );
	vdp_slatch g4230 (.Q(w3445), .D(S[7]), .C(w3421), .nC(w3482) );
	vdp_slatch g4231 (.Q(w3446), .D(S[6]), .C(w3421), .nC(w3482) );
	vdp_slatch g4232 (.Q(w3444), .D(S[5]), .C(w3421), .nC(w3482) );
	vdp_slatch g4233 (.Q(w3443), .D(S[4]), .C(w3421), .nC(w3482) );
	vdp_slatch g4234 (.Q(w3441), .D(S[3]), .C(w3421), .nC(w3482) );
	vdp_slatch g4235 (.Q(w3439), .D(S[2]), .C(w3421), .nC(w3482) );
	vdp_slatch g4236 (.Q(w3437), .D(S[1]), .C(w3421), .nC(w3482) );
	vdp_slatch g4237 (.Q(w3434), .D(S[0]), .C(w3421), .nC(w3482) );
	vdp_sr_bit g4238 (.Q(w3985), .D(w3415), .C1(HCLK2), .C2(HCLK1), .nC2(nHCLK1), .nC1(nHCLK2) );
	vdp_sr_bit g4239 (.Q(w3422), .D(w3953), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and g4240 (.Z(w3953), .A(w13), .B(M5) );
	vdp_not g4241 (.nZ(w3952), .A(w3422) );
	vdp_aon22 g4242 (.Z(w2997), .A1(w3956), .B1(w3486), .A2(w3485), .B2(w3917) );
	vdp_aon22 g4243 (.Z(w2994), .A1(w3955), .B1(1'b0), .A2(w3485), .B2(w3917) );
	vdp_aon22 g4244 (.Z(w3484), .A1(w3486), .B1(w3452), .A2(w3485), .B2(w3917) );
	vdp_aon22 g4245 (.Z(w2968), .A1(w3487), .B1(w3450), .A2(w3485), .B2(w3917) );
	vdp_aon22 g4246 (.Z(w2971), .A1(w3954), .B1(w3487), .A2(w3485), .B2(w3917) );
	vdp_comp_strong g4247 (.Z(w3421), .nZ(w3482), .A(w3184) );
	vdp_comp_we g4248 (.Z(w3485), .nZ(w3917), .A(M5) );
	vdp_aon22 g4249 (.Z(w3426), .A1(w3483), .B1(w3484), .A2(w3422), .B2(w3952) );
	vdp_sr_bit g4250 (.Q(w3870), .D(FIFOo[0]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4251 (.Q(w3874), .D(FIFOo[1]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4252 (.Q(w3872), .D(FIFOo[2]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4253 (.Q(w3871), .D(FIFOo[3]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4254 (.Q(w3859), .D(FIFOo[4]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4255 (.Q(w3857), .D(FIFOo[5]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4256 (.Q(w3864), .D(FIFOo[6]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4257 (.Q(w3866), .D(FIFOo[7]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_aon22 g4258 (.Z(w1357), .B1(w4328), .A1(w1384), .B2(w4346), .A2(w43) );
	vdp_not g4259 (.nZ(w4346), .A(w43) );
	vdp_not g4260 (.nZ(w4318), .A(w4307) );
	vdp_not g4261 (.nZ(w4317), .A(w4318) );
	vdp_not g4262 (.nZ(w4316), .A(w4317) );
	vdp_not g4263 (.nZ(w4315), .A(w4316) );
	vdp_and g4264 (.Z(w4328), .B(w4319), .A(w4323) );
	vdp_not g4265 (.nZ(w4319), .A(w4322) );
	vdp_not g4266 (.nZ(w4322), .A(w4321) );
	vdp_not g4267 (.nZ(w4321), .A(w4320) );
	vdp_not g4268 (.nZ(w4320), .A(w4323) );
	vdp_or g4269 (.Z(w4323), .B(w4305), .A(w4304) );
	vdp_dff g4270 (.Q(w4305), .R(w4294), .D(w4304), .C(w4303) );
	vdp_not g4271 (.nZ(w4303), .A(w4324) );
	vdp_nor g4272 (.Z(w4302), .B(w4325), .A(w4304) );
	vdp_dff g4273 (.Q(w4304), .R(w4294), .D(w4325), .C(w4324) );
	vdp_dff g4274 (.Q(w4325), .R(w4294), .D(w4302), .C(w4324) );
	vdp_not g4275 (.nZ(w4324), .A(w4313) );
	vdp_not g4276 (.nZ(w4300), .A(w4313) );
	vdp_dff g4277 (.Q(w4297), .R(w4294), .D(w4326), .C(w4296) );
	vdp_dff g4278 (.Q(w4326), .R(w4294), .D(w4295), .C(w4293) );
	vdp_not g4279 (.nZ(w4293), .A(w4334) );
	vdp_dff g4280 (.Q(w4295), .R(w4294), .D(w4314), .C(w4293) );
	vdp_not g4281 (.nZ(w4296), .A(w4293) );
	vdp_nor g4282 (.Z(w4353), .B(w4329), .A(w4330) );
	vdp_nor g4283 (.Z(w4331), .B(w4329), .A(H40) );
	vdp_not g4284 (.nZ(w4330), .A(H40) );
	vdp_not g4285 (.nZ(w4308), .A(PAL) );
	vdp_AOI222 g4286 (.Z(w4301), .B1(w4333), .A1(w4332), .B2(w4353), .A2(w4329), .C1(w4300), .C2(w4331) );
	vdp_not g4287 (.nZ(EDCLK_O), .A(w4301) );
	vdp_or g4288 (.Z(w4327), .B(w4297), .A(w4326) );
	vdp_nor g4289 (.Z(w4314), .B(w4295), .A(w4326) );
	vdp_not g4290 (.nZ(w4290), .A(w4352) );
	vdp_nand g4291 (.Z(w4309), .B(w4290), .A(w4289) );
	vdp_sr_bit g4292 (.Q(w4352), .D(w4289), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_not g4293 (.nZ(w4351), .A(w4337) );
	vdp_not g4294 (.nZ(w1128), .A(w4350) );
	vdp_not g4295 (.nZ(SYSRES), .A(w4351) );
	vdp_comp_dff g4296 (.Q(w4289), .D(w4337), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_not g4297 (.nZ(w4347), .A(w4348) );
	vdp_not g4298 (.nZ(w4294), .A(w4349) );
	vdp_not g4299 (.nZ(w4336), .A(w4335) );
	vdp_nand g4300 (.Z(w4349), .B(w4336), .A(w4292) );
	vdp_not g4301 (.nZ(w4334), .A(w4338) );
	vdp_nand g4302 (.Z(w4341), .B(w4340), .A(w4339) );
	vdp_not g4303 (.nZ(w4313), .A(w4298) );
	vdp_nand g4304 (.Z(w4344), .B(w4343), .A(w4342) );
	vdp_not g4305 (.nZ(w4307), .A(w4312) );
	vdp_not g4306 (.nZ(RES), .A(w4309) );
	vdp_dff g4307 (.Q(w4292), .R(1'b0), .D(w4337), .C(w4310) );
	vdp_dff g4308 (.Q(w4335), .R(1'b0), .D(w4292), .C(w4310) );
	vdp_dff g4309 (.Q(w4348), .R(w4294), .D(w4338), .C(w4310) );
	vdp_dff g4310 (.Q(w4338), .R(w4294), .D(w4347), .C(w4310) );
	vdp_dff g4311 (.Q(w4339), .R(w4294), .D(w4298), .C(w4310) );
	vdp_dff g4312 (.Q(w4340), .R(w4294), .D(w4339), .C(w4310) );
	vdp_dff g4313 (.Q(w4298), .R(w4294), .D(w4341), .C(w4310) );
	vdp_dff g4314 (.Q(w4342), .R(w4294), .D(w4312), .C(w4310) );
	vdp_dff g4315 (.Q(w4343), .R(w4294), .D(w4342), .C(w4310) );
	vdp_dff g4316 (.Q(w4345), .R(w4294), .D(w4344), .C(w4310) );
	vdp_dff g4317 (.Q(w4312), .R(w4294), .D(w4345), .C(w4310) );
	vdp_not g4318 (.nZ(w4333), .A(w4334) );
	vdp_nand g4319 (.Z(w4337), .B(w1385), .A(w4350) );
	vdp_not g4320 (.nZ(M68K_CPU_CLOCK), .A(w4306) );
	vdp_or g4321 (.Z(w4329), .B(w43), .A(RS0) );
	vdp_aon22 g4322 (.Z(w4299), .B1(w4327), .A1(w4328), .B2(PAL), .A2(w4308) );
	vdp_or g4323 (.Z(w4306), .B(w4315), .A(w4307) );
	vdp_comp_we g4324 (.A(w2546), .nZ(nHCLK2), .Z(HCLK2) );
	vdp_comp_we g4325 (.A(w2545), .nZ(nHCLK1), .Z(HCLK1) );
	vdp_comp_we g4326 (.A(w4360), .nZ(nDCLK2), .Z(DCLK2) );
	vdp_comp_we g4327 (.A(EDCLK_O), .nZ(nDCLK1), .Z(DCLK1) );
	vdp_not g4328 (.nZ(w4360), .A(EDCLK_O) );
	vdp_sr_bit g4329 (.Q(w4455), .D(w4454), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4330 (.Q(w4473), .D(w4450), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4331 (.Q(w4450), .D(w4435), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4332 (.Q(w4435), .D(w4427), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4333 (.Q(w4430), .D(w6288), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4334 (.Q(w6288), .D(w6289), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4335 (.Q(w6289), .D(w6291), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4336 (.Q(w6291), .D(w6290), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4337 (.Q(w6290), .D(w6292), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4338 (.Q(w6292), .D(w6293), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4339 (.Q(w6293), .D(w6295), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4340 (.Q(w6295), .D(w6294), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4341 (.Q(w6294), .D(w6168), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4342 (.Q(w6168), .D(w4375), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4343 (.Q(w4411), .D(w4412), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4344 (.Q(w4412), .D(w23), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4345 (.Q(w4669), .D(w6296), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4346 (.Q(w4380), .D(w4703), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4347 (.Q(w4379), .D(w6284), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4348 (.Q(w6031), .D(w4457), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4349 (.Q(w4456), .D(w6297), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4350 (.Q(w4458), .D(w4448), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4351 (.Q(w6286), .D(w4), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4352 (.Q(w4399), .D(w4420), .nC(w4423), .C(w4424) );
	vdp_slatch g4353 (.Q(w4404), .D(w4421), .nC(w4423), .C(w4424) );
	vdp_slatch g4354 (.Q(w4391), .D(w4422), .nC(w4423), .C(w4424) );
	vdp_slatch g4355 (.Q(w4383), .D(w4428), .nC(w4423), .C(w4424) );
	vdp_slatch g4356 (.Q(w4382), .D(w4419), .nC(w4423), .C(w4424) );
	vdp_slatch g4357 (.Q(w4381), .D(w4418), .nC(w4423), .C(w4424) );
	vdp_slatch g4358 (.Q(w4432), .D(w4417), .nC(w4423), .C(w4424) );
	vdp_slatch g4359 (.Q(w4384), .D(w4415), .nC(w4423), .C(w4424) );
	vdp_slatch g4360 (.Q(w4387), .D(w4416), .nC(w4423), .C(w4424) );
	vdp_slatch g4361 (.Q(w4388), .D(w4414), .nC(w4423), .C(w4424) );
	vdp_comp_str g4362 (.nZ(w4423), .A(w4429), .Z(w4424) );
	vdp_sr_bit g4363 (.Q(w4451), .D(w4474), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4364 (.Q(w6017), .D(w38), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_xor g4365 (.Z(w4397), .B(w4389), .A(w4400) );
	vdp_xor g4366 (.Z(w4392), .B(w4390), .A(w4398) );
	vdp_xor g4367 (.Z(w4394), .B(w4377), .A(w4391) );
	vdp_xor g4368 (.Z(w6120), .B(w4377), .A(w4383) );
	vdp_xor g4369 (.Z(w6121), .B(w4377), .A(w4382) );
	vdp_xor g4370 (.Z(w6116), .B(w4377), .A(w4381) );
	vdp_aon22 g4371 (.Z(w6117), .B2(w4405), .B1(w4399), .A1(w4397), .A2(w4393) );
	vdp_aon22 g4372 (.Z(w6118), .B2(w4405), .B1(w4397), .A1(w4392), .A2(w4393) );
	vdp_aon22 g4373 (.Z(w6119), .B2(w4405), .B1(w4392), .A1(w4394), .A2(w4393) );
	vdp_aon22 g4374 (.Z(w4395), .B2(w4386), .B1(w4391), .A1(w4404), .A2(w4396) );
	vdp_aon22 g4375 (.Z(w4401), .B2(w4386), .B1(w4404), .A1(w4399), .A2(w4396) );
	vdp_aon22 g4376 (.Z(w4466), .B2(w4459), .B1(w4462), .A1(w4463), .A2(w72) );
	vdp_aon22 g4377 (.Z(w4467), .B2(w4461), .B1(w4462), .A1(w4463), .A2(w71) );
	vdp_aon22 g4378 (.Z(w4468), .B2(w4460), .B1(w4462), .A1(w4463), .A2(w70) );
	vdp_aon22 g4379 (.Z(w4469), .B2(w4464), .B1(w4462), .A1(w4463), .A2(w69) );
	vdp_aon22 g4380 (.Z(w4470), .B2(w4465), .B1(w4462), .A1(w4463), .A2(w68) );
	vdp_not g4381 (.nZ(w4436), .A(w4375) );
	vdp_not g4382 (.nZ(w4408), .A(w4440) );
	vdp_not g4383 (.nZ(w4439), .A(w107) );
	vdp_not g4384 (.nZ(w4444), .A(w4442) );
	vdp_not g4385 (.nZ(w4431), .A(M5) );
	vdp_not g4386 (.nZ(w4472), .A(w73) );
	vdp_not g4387 (.nZ(w4471), .A(w74) );
	vdp_not g4388 (.nZ(w4446), .A(1'b0) );
	vdp_not g4389 (.nZ(w4447), .A(M5) );
	vdp_not g4390 (.nZ(w4374), .A(w4375) );
	vdp_not g4391 (.nZ(w4378), .A(w4409) );
	vdp_not g4392 (.nZ(w4385), .A(w4388) );
	vdp_not g4393 (.nZ(w4390), .A(w4426) );
	vdp_and g4394 (.Z(w4427), .B(w4436), .A(w4437) );
	vdp_and g4395 (.Z(w4441), .B(w4439), .A(w4450) );
	vdp_or g4396 (.Z(w4438), .B(w4441), .A(w4453) );
	vdp_or g4397 (.Z(w4434), .B(w4476), .A(w4441) );
	vdp_and g4398 (.Z(w4452), .B(w4445), .A(1'b0) );
	vdp_and g4399 (.Z(w4475), .B(w4445), .A(w4446) );
	vdp_or g4400 (.Z(w4474), .B(w38), .A(w37) );
	vdp_and g4401 (.Z(SPRITE_OVF), .B(w6429), .A(w4) );
	vdp_and g4402 (.Z(w6284), .B(w4374), .A(w4376) );
	vdp_or g4403 (.Z(w4425), .B(w4380), .A(w4379) );
	vdp_and g4404 (.Z(w4389), .B(w4384), .A(w4377) );
	vdp_comp_we g4405 (.nZ(w4386), .A(w1), .Z(w4396) );
	vdp_comp_we g4406 (.nZ(w4405), .A(w1), .Z(w4393) );
	vdp_comp_we g4407 (.nZ(w4462), .A(w107), .Z(w4463) );
	vdp_not g4408 (.nZ(w4477), .A(w4454) );
	vdp_rs_ff g4409 (.Q(w6285), .R(w6286), .S(w4425) );
	vdp_rs_ff g4410 (.Q(w6429), .R(w6286), .S(w4379) );
	vdp_ha g4411 (.SUM(w4400), .B(w4401), .A(w4402) );
	vdp_ha g4412 (.SUM(w4398), .B(w4395), .A(w4403), .CO(w4402) );
	vdp_not g4413 (.nZ(w4410), .A(w4373) );
	vdp_and g4414 (.Z(w4413), .B(w4375), .A(w4376) );
	vdp_and3 g4415 (.Z(w4403), .B(w4384), .A(w4377), .C(w4385) );
	vdp_and3 g4416 (.Z(w4457), .B(w4455), .A(M5), .C(w4477) );
	vdp_and3 g4417 (.Z(w6297), .B(w4460), .A(w4459), .C(w4458) );
	vdp_and3 g4418 (.Z(w4476), .B(w74), .A(w4472), .C(w111) );
	vdp_and3 g4419 (.Z(w6287), .B(w73), .A(w4471), .C(w111) );
	vdp_and3 g4420 (.Z(w4453), .B(w4472), .A(w4471), .C(w111) );
	vdp_or3 g4421 (.Z(w4433), .B(w6287), .A(w4441), .C(w4444) );
	vdp_and3 g4422 (.Z(w4429), .B(HCLK1), .A(w4411), .C(DCLK1) );
	vdp_or3 g4423 (.Z(w4445), .B(w4448), .A(w4473), .C(w4447) );
	vdp_oai21 g4424 (.Z(w4426), .B(w4377), .A1(w4384), .A2(w4388) );
	vdp_nor g4425 (.Z(w4373), .B(w4413), .A(w4412) );
	vdp_nor g4426 (.Z(w6296), .B(w4378), .A(w6285) );
	vdp_nand g4427 (.Z(w4449), .B(w4431), .A(w4430) );
	vdp_nand g4428 (.Z(w4407), .B(w4472), .A(w4471) );
	vdp_nand g4429 (.Z(w4440), .B(w73), .A(w4471) );
	vdp_nand g4430 (.Z(w4406), .B(w74), .A(w4472) );
	vdp_nor g4431 (.Z(w4454), .B(w4456), .A(w4371) );
	vdp_cnt_bit_rev g4432 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4459), .CI(w4481), .B(w4451), .A(w4452) );
	vdp_cnt_bit_rev g4433 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4461), .CI(w4480), .B(w4451), .A(w4452), .CO(w4481) );
	vdp_cnt_bit_rev g4434 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4460), .CI(w4479), .B(w4451), .A(w4452), .CO(w4480) );
	vdp_cnt_bit_rev g4435 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4464), .CI(w4478), .B(w4451), .A(w4452), .CO(w4479) );
	vdp_cnt_bit_rev g4436 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4465), .CI(w4475), .B(w4451), .A(w4452), .CO(w4478) );
	vdp_cnt_bit_load g4437 (.Q(w4488), .D(w4528), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4490), .CI(w6332), .L(w4529), .nL(w4494) );
	vdp_cnt_bit_load g4438 (.Q(w4491), .D(w4533), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4490), .CI(w6331), .L(w4529), .nL(w4494), .CO(w6332) );
	vdp_cnt_bit_load g4439 (.Q(w4493), .D(w4534), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4490), .CI(w6330), .L(w4529), .nL(w4494), .CO(w6331) );
	vdp_cnt_bit_load g4440 (.Q(w4495), .D(w4558), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4490), .CI(w6329), .L(w4529), .nL(w4494), .CO(w6330) );
	vdp_cnt_bit_load g4441 (.Q(w4499), .D(w4559), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4490), .CI(w6328), .L(w4529), .nL(w4494), .CO(w6329) );
	vdp_cnt_bit_load g4442 (.Q(w4496), .D(w4560), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4490), .CI(w6327), .L(w4529), .nL(w4494), .CO(w6328) );
	vdp_cnt_bit_load g4443 (.Q(w4492), .D(w4561), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4490), .CI(w4489), .L(w4529), .nL(w4494), .CO(w6327) );
	vdp_fa g4444 (.SUM(w4636), .CO(w6342), .CI(1'b1), .A(w4691), .B(w4639) );
	vdp_fa g4445 (.SUM(w4638), .CO(w6343), .CI(w6342), .A(w4690), .B(w4643) );
	vdp_fa g4446 (.SUM(w4644), .CO(w6344), .CI(w6343), .A(w4689), .B(w4647) );
	vdp_fa g4447 (.SUM(w4646), .CO(w6345), .CI(w6344), .A(w4688), .B(w4649) );
	vdp_fa g4448 (.SUM(w4651), .CO(w6346), .CI(w6345), .A(w4687), .B(w4653) );
	vdp_fa g4449 (.SUM(w4657), .CO(w6347), .CI(w6346), .A(w4686), .B(w4682) );
	vdp_fa g4450 (.SUM(w4660), .CO(w6348), .CI(w6347), .A(w4684), .B(w4659) );
	vdp_fa g4451 (.SUM(w4664), .CO(w6349), .CI(w6348), .A(w4696), .B(w4663) );
	vdp_fa g4452 (.SUM(w4666), .CO(w6350), .CI(w6349), .A(w4697), .B(w4665) );
	vdp_fa g4453 (.SUM(w4680), .CI(w6350), .A(w4701), .B(w4679) );
	vdp_fa g4454 (.SUM(w4691), .CO(w6333), .CI(1'b0), .A(VPOS[0]), .B(w4692) );
	vdp_fa g4455 (.SUM(w4690), .CO(w6334), .CI(w6333), .A(VPOS[1]), .B(w1) );
	vdp_fa g4456 (.SUM(w4689), .CO(w6335), .CI(w6334), .A(VPOS[2]), .B(1'b0) );
	vdp_fa g4457 (.SUM(w4688), .CO(w6336), .CI(w6335), .A(VPOS[3]), .B(1'b0) );
	vdp_fa g4458 (.SUM(w4687), .CO(w6337), .CI(w6336), .A(VPOS[4]), .B(1'b0) );
	vdp_fa g4459 (.SUM(w4686), .CO(w6338), .CI(w6337), .A(VPOS[5]), .B(1'b0) );
	vdp_fa g4460 (.SUM(w4684), .CO(w6339), .CI(w6338), .A(VPOS[6]), .B(1'b0) );
	vdp_fa g4461 (.SUM(w4696), .CO(w6340), .CI(w6339), .A(VPOS[7]), .B(w4692) );
	vdp_fa g4462 (.SUM(w4697), .CO(w6341), .CI(w6340), .A(VPOS[8]), .B(w1) );
	vdp_fa g4463 (.SUM(w4701), .CI(w6341), .A(VPOS[9]), .B(1'b0) );
	vdp_slatch g4464 (.nC(w4584), .C(w4583), .Q(w4629), .D(S[0]) );
	vdp_dlatch_inv g4465 (.nQ(w4628), .D(w4597), .nC(nHCLK2), .C(HCLK2) );
	vdp_slatch g4466 (.nC(w4569), .C(w4568), .Q(w4597), .D(w4586) );
	vdp_slatch g4467 (.nC(w4584), .C(w4583), .Q(w4626), .D(S[1]) );
	vdp_slatch g4468 (.nC(w4569), .C(w4568), .Q(w6372), .D(w4588) );
	vdp_slatch g4469 (.nC(w4584), .C(w4583), .Q(w4624), .D(S[2]) );
	vdp_slatch g4470 (.nC(w4569), .C(w4568), .Q(w6373), .D(w4579) );
	vdp_slatch g4471 (.nC(w4584), .C(w4583), .Q(w4622), .D(S[3]) );
	vdp_slatch g4472 (.nC(w4569), .C(w4568), .Q(w6374), .D(w4575) );
	vdp_slatch g4473 (.nC(w4584), .C(w4583), .Q(w4619), .D(S[4]) );
	vdp_slatch g4474 (.nC(w4569), .C(w4568), .Q(w6375), .D(w4571) );
	vdp_slatch g4475 (.nC(w4584), .C(w4583), .Q(w4618), .D(S[5]) );
	vdp_slatch g4476 (.nC(w4569), .C(w4568), .Q(w6376), .D(w4567) );
	vdp_slatch g4477 (.nC(w4584), .C(w4583), .Q(w4615), .D(S[6]) );
	vdp_slatch g4478 (.nC(w4569), .C(w4568), .Q(w6377), .D(w6319) );
	vdp_slatch g4479 (.nC(w4584), .C(w4583), .Q(w6378), .D(S[7]) );
	vdp_slatch g4480 (.nC(w4569), .C(w4568), .Q(w6379), .D(w4599) );
	vdp_slatch g4481 (.nC(w4569), .C(w4568), .Q(w4600), .D(w4601) );
	vdp_slatch g4482 (.nC(w4569), .C(w4568), .Q(w6380), .D(w4603) );
	vdp_dlatch_inv g4483 (.nQ(w4625), .D(w6372), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4484 (.nQ(w4623), .D(w6373), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4485 (.nQ(w4621), .D(w6374), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4486 (.nQ(w4620), .D(w6375), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4487 (.nQ(w4617), .D(w6376), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4488 (.nQ(w4614), .D(w6377), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4489 (.nQ(w4613), .D(w6379), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4490 (.nQ(w4612), .D(w4600), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4491 (.nQ(w4602), .D(w6380), .nC(nHCLK2), .C(HCLK2) );
	vdp_sr_bit g4492 (.Q(w4554), .D(w4485), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4493 (.Z(w4409), .B2(w4550), .B1(w4556), .A1(M5), .A2(w4555) );
	vdp_sr_bit g4494 (.Q(w4485), .D(w4551), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4495 (.Q(w4551), .D(w4552), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4496 (.Q(w4552), .D(w4530), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4497 (.Q(w4591), .D(w4593), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4498 (.Q(w4582), .D(w4596), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4499 (.Q(w4578), .D(w4589), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4500 (.Q(w4574), .D(w4590), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4501 (.Q(w4570), .D(w4572), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4502 (.Q(w4566), .D(w4564), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4503 (.Q(w4598), .D(w4565), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4504 (.Q(w6381), .D(w4563), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4505 (.Q(w4512), .D(w4562), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4506 (.Q(w4519), .D(w4557), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4507 (.Q(w4553), .D(w4486), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4508 (.Q(w4486), .D(w4508), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4509 (.Q(w4738), .D(w119), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4510 (.Q(w4740), .D(VRAMA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4511 (.Q(w4508), .D(w8), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4512 (.Q(w4741), .D(w6326), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4513 (.Q(w6326), .D(w4738), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4514 (.Q(w6370), .D(w4724), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4515 (.Q(w6368), .D(w4727), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4516 (.Q(w6366), .D(w4743), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4517 (.Q(w6364), .D(w4704), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4518 (.Q(w6362), .D(w4528), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4519 (.Q(w6360), .D(w4533), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4520 (.Q(w6358), .D(w4534), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4521 (.Q(w6356), .D(w4558), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4522 (.Q(w6354), .D(w4559), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4523 (.Q(w6352), .D(w4560), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4524 (.Q(w4722), .D(w4561), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4525 (.Q(w4714), .D(w6351), .nC(w4713), .C(w4705) );
	vdp_dlatch_inv g4526 (.nQ(w6351), .D(w4722), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4527 (.Q(w4715), .D(w6353), .nC(w4713), .C(w4705) );
	vdp_dlatch_inv g4528 (.nQ(w6353), .D(w6352), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4529 (.Q(w4716), .D(w6355), .nC(w4713), .C(w4705) );
	vdp_dlatch_inv g4530 (.nQ(w6355), .D(w6354), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4531 (.Q(w4717), .D(w6357), .nC(w4713), .C(w4705) );
	vdp_dlatch_inv g4532 (.nQ(w6357), .D(w6356), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4533 (.Q(w4718), .D(w6359), .nC(w4713), .C(w4705) );
	vdp_dlatch_inv g4534 (.nQ(w6359), .D(w6358), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4535 (.Q(w6325), .D(w6361), .nC(w4713), .C(w4705) );
	vdp_dlatch_inv g4536 (.nQ(w6361), .D(w6360), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4537 (.Q(w4719), .D(w6363), .nC(w4713), .C(w4705) );
	vdp_dlatch_inv g4538 (.nQ(w6363), .D(w6362), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4539 (.Q(w4709), .D(w6365), .nC(w4713), .C(w4705) );
	vdp_dlatch_inv g4540 (.nQ(w6365), .D(w6364), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4541 (.Q(w4712), .D(w6367), .nC(w4713), .C(w4705) );
	vdp_dlatch_inv g4542 (.nQ(w6367), .D(w6366), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4543 (.Q(w4710), .D(w6369), .nC(w4713), .C(w4705) );
	vdp_dlatch_inv g4544 (.nQ(w6369), .D(w6368), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4545 (.Q(w4711), .D(w6371), .nC(w4713), .C(w4705) );
	vdp_dlatch_inv g4546 (.nQ(w6371), .D(w6370), .nC(nHCLK1), .C(HCLK1) );
	vdp_aon22 g4547 (.Z(w6186), .B2(w4538), .B1(w4488), .A1(w4487), .A2(w6166) );
	vdp_aon22 g4548 (.Z(w6187), .B2(w4538), .B1(w4491), .A1(w4487), .A2(w4543) );
	vdp_aon22 g4549 (.Z(w6188), .B2(w4538), .B1(w4493), .A1(w4487), .A2(w4542) );
	vdp_aon22 g4550 (.Z(w6189), .B2(w4538), .B1(w4495), .A1(w4487), .A2(w4541) );
	vdp_aon22 g4551 (.Z(w6190), .B2(w4538), .B1(w4499), .A1(w4487), .A2(w4540) );
	vdp_aon22 g4552 (.Z(w6192), .B2(w4538), .B1(w4496), .A1(w4487), .A2(w4539) );
	vdp_aon22 g4553 (.Z(w6191), .B2(w4538), .B1(w4492), .A1(w4487), .A2(w4537) );
	vdp_aon22 g4554 (.Z(w4755), .B2(w4501), .B1(w3), .A1(w4497), .A2(w4492) );
	vdp_aon22 g4555 (.Z(w4650), .B2(w4610), .B1(w4619), .A1(w4620), .A2(w4634) );
	vdp_2x_sr_bit g4556 (.Q(w4549), .D(w4492), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4557 (.Z(w6167), .B2(w4501), .B1(w4549), .A1(w4497), .A2(w4496) );
	vdp_2x_sr_bit g4558 (.Q(w4498), .D(w4496), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4559 (.Z(w4808), .B2(w4501), .B1(w4498), .A1(w4497), .A2(w4499) );
	vdp_2x_sr_bit g4560 (.Q(w4536), .D(w4499), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4561 (.Z(w4814), .B2(w4501), .B1(w4536), .A1(w4497), .A2(w4495) );
	vdp_2x_sr_bit g4562 (.Q(w4500), .D(w4495), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4563 (.Z(w4863), .B2(w4501), .B1(w4500), .A1(w4497), .A2(w4493) );
	vdp_2x_sr_bit g4564 (.Q(w4503), .D(w4493), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4565 (.Z(w4914), .B2(w4501), .B1(w4503), .A1(w4497), .A2(w4491) );
	vdp_aon22 g4566 (.Z(w4928), .B2(w4501), .B1(1'b1), .A1(w4497), .A2(w4488) );
	vdp_aon22 g4567 (.Z(w4586), .B2(w4511), .B1(w4587), .A1(w4514), .A2(w4585) );
	vdp_dlatch_inv g4568 (.nQ(w4585), .D(w4591), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4569 (.nZ(w4587), .A(S[0]) );
	vdp_aon22 g4570 (.Z(w4588), .B2(w4511), .B1(w4581), .A1(w4514), .A2(w4580) );
	vdp_dlatch_inv g4571 (.nQ(w4580), .D(w4582), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4572 (.nZ(w4581), .A(S[1]) );
	vdp_aon22 g4573 (.Z(w4579), .B2(w4511), .B1(w4577), .A1(w4514), .A2(w4576) );
	vdp_dlatch_inv g4574 (.nQ(w4576), .D(w4578), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4575 (.nZ(w4577), .A(S[2]) );
	vdp_aon22 g4576 (.Z(w4575), .B2(w4511), .B1(w4535), .A1(w4514), .A2(w4573) );
	vdp_dlatch_inv g4577 (.nQ(w4573), .D(w4574), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4578 (.nZ(w4535), .A(S[3]) );
	vdp_aon22 g4579 (.Z(w4571), .B2(w4511), .B1(w4531), .A1(w4514), .A2(w4532) );
	vdp_dlatch_inv g4580 (.nQ(w4532), .D(w4570), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4581 (.nZ(w4531), .A(S[4]) );
	vdp_aon22 g4582 (.Z(w4567), .B2(w4511), .B1(w4527), .A1(w4514), .A2(w4526) );
	vdp_dlatch_inv g4583 (.nQ(w4526), .D(w4566), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4584 (.nZ(w4527), .A(S[5]) );
	vdp_aon22 g4585 (.Z(w6319), .B2(w4511), .B1(w4522), .A1(w4514), .A2(w4521) );
	vdp_dlatch_inv g4586 (.nQ(w4521), .D(w4598), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4587 (.nZ(w4522), .A(S[6]) );
	vdp_aon22 g4588 (.Z(w4599), .B2(w4511), .B1(w4515), .A1(w4514), .A2(w4513) );
	vdp_dlatch_inv g4589 (.nQ(w4513), .D(w6381), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4590 (.nZ(w4515), .A(S[7]) );
	vdp_aon22 g4591 (.Z(w4601), .B2(w4511), .B1(w4750), .A1(w4514), .A2(1'b1) );
	vdp_dlatch_inv g4592 (.nQ(w4750), .D(w4512), .nC(nHCLK1), .C(HCLK1) );
	vdp_aon22 g4593 (.Z(w4603), .B2(w4511), .B1(1'b1), .A1(w4514), .A2(w4520) );
	vdp_dlatch_inv g4594 (.nQ(w4520), .D(w4519), .nC(nHCLK1), .C(HCLK1) );
	vdp_sr_bit g4595 (.Q(w4490), .D(w6314), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4596 (.Q(w4502), .D(w28), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4597 (.Q(w4523), .D(w4502), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4598 (.Q(w4507), .D(w5), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4599 (.Q(w4517), .D(w4507), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4600 (.Q(w4530), .D(w6313), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_not g4601 (.nZ(w4525), .A(w4524) );
	vdp_not g4602 (.nZ(w4518), .A(M5) );
	vdp_not g4603 (.nZ(w6314), .A(w4516) );
	vdp_not g4604 (.nZ(w4506), .A(w4517) );
	vdp_not g4605 (.nZ(w6313), .A(w4509) );
	vdp_not g4606 (.nZ(w4504), .A(w4489) );
	vdp_aon22 g4607 (.Z(w4609), .B2(w4605), .B1(w4422), .A1(w4604), .A2(w4421) );
	vdp_aon22 g4608 (.Z(w4608), .B2(w4605), .B1(w4421), .A1(w4604), .A2(w4420) );
	vdp_aon22 g4609 (.Z(w4607), .B2(w4605), .B1(w4420), .A1(w4604), .A2(1'b0) );
	vdp_slatch g4610 (.nQ(w6390), .D(w4737), .nC(w4721), .C(w4726) );
	vdp_aon22 g4611 (.Z(w4737), .B2(w4720), .B1(w4593), .A1(w4725), .A2(w4561) );
	vdp_notif0 g4612 (.A(w6390), .nZ(AD_DATA[0]), .nE(w4731) );
	vdp_slatch g4613 (.nQ(w6389), .D(w4736), .nC(w4721), .C(w4726) );
	vdp_aon22 g4614 (.Z(w4736), .B2(w4720), .B1(w4596), .A1(w4725), .A2(w4560) );
	vdp_notif0 g4615 (.A(w6389), .nZ(AD_DATA[1]), .nE(w4731) );
	vdp_slatch g4616 (.nQ(w6388), .D(w4735), .nC(w4721), .C(w4726) );
	vdp_aon22 g4617 (.Z(w4735), .B2(w4720), .B1(w4589), .A1(w4725), .A2(w4559) );
	vdp_notif0 g4618 (.A(w6388), .nZ(AD_DATA[2]), .nE(w4731) );
	vdp_slatch g4619 (.nQ(w6387), .D(w6323), .nC(w4721), .C(w4726) );
	vdp_aon22 g4620 (.Z(w6323), .B2(w4720), .B1(w4590), .A1(w4725), .A2(w4558) );
	vdp_notif0 g4621 (.A(w6387), .nZ(AD_DATA[3]), .nE(w4731) );
	vdp_slatch g4622 (.nQ(w6386), .D(w6322), .nC(w4721), .C(w4726) );
	vdp_aon22 g4623 (.Z(w6322), .B2(w4720), .B1(w4572), .A1(w4725), .A2(w4534) );
	vdp_notif0 g4624 (.A(w6386), .nZ(AD_DATA[4]), .nE(w4731) );
	vdp_slatch g4625 (.nQ(w6385), .D(w6321), .nC(w4721), .C(w4726) );
	vdp_aon22 g4626 (.Z(w6321), .B2(w4720), .B1(w4564), .A1(w4725), .A2(w4533) );
	vdp_notif0 g4627 (.A(w6385), .nZ(AD_DATA[5]), .nE(w4731) );
	vdp_slatch g4628 (.nQ(w6384), .D(w4734), .nC(w4721), .C(w4726) );
	vdp_aon22 g4629 (.Z(w4734), .B2(w4720), .B1(w4565), .A1(w4725), .A2(w4528) );
	vdp_notif0 g4630 (.A(w6384), .nZ(AD_DATA[6]), .nE(w4731) );
	vdp_slatch g4631 (.nQ(w6383), .D(w4742), .nC(w4721), .C(w4726) );
	vdp_aon22 g4632 (.Z(w4742), .B2(w4720), .B1(w4563), .A1(w4725), .A2(w4704) );
	vdp_notif0 g4633 (.A(w6383), .nZ(AD_DATA[7]), .nE(w4731) );
	vdp_slatch g4634 (.nQ(w4733), .D(w4732), .nC(w4721), .C(w4726) );
	vdp_aon22 g4635 (.Z(w4732), .B2(w4720), .B1(w4562), .A1(w4725), .A2(w4743) );
	vdp_notif0 g4636 (.A(w4733), .nZ(RD_DATA[0]), .nE(w4731) );
	vdp_slatch g4637 (.nQ(w4730), .D(w4729), .nC(w4721), .C(w4726) );
	vdp_aon22 g4638 (.Z(w4729), .B2(w4720), .B1(w4557), .A1(w4725), .A2(w4727) );
	vdp_notif0 g4639 (.A(w4730), .nZ(RD_DATA[1]), .nE(w4731) );
	vdp_slatch g4640 (.nQ(w4728), .D(w4723), .nC(w4721), .C(w4726) );
	vdp_aon22 g4641 (.Z(w4723), .B2(w4720), .B1(1'b0), .A1(w4725), .A2(w4724) );
	vdp_notif0 g4642 (.A(w4728), .nZ(RD_DATA[2]), .nE(w4731) );
	vdp_not g4643 (.nZ(w4731), .A(w4741) );
	vdp_sr_bit g4644 (.Q(w4415), .D(w6394), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4645 (.Q(w4416), .D(w4699), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4646 (.Q(w4695), .D(w4693), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_dlatch_inv g4647 (.nQ(w4694), .D(w4595), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4648 (.nQ(w4693), .D(w4633), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g4649 (.nQ(w4639), .D(w4635), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4650 (.nQ(w6320), .D(w4636), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4651 (.nQ(w4643), .D(w4637), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4652 (.nQ(w4641), .D(w4638), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4653 (.nQ(w4647), .D(w4642), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4654 (.nQ(w4645), .D(w4644), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4655 (.nQ(w4649), .D(w4648), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4656 (.nQ(w4658), .D(w4646), .nC(nHCLK2), .C(HCLK2) );
	vdp_aon22 g4657 (.Z(w4648), .B2(w4610), .B1(w4622), .A1(w4621), .A2(w4634) );
	vdp_aon22 g4658 (.Z(w4642), .B2(w4610), .B1(w4624), .A1(w4623), .A2(w4634) );
	vdp_aon22 g4659 (.Z(w4637), .B2(w4610), .B1(w4626), .A1(w4625), .A2(w4634) );
	vdp_aon22 g4660 (.Z(w4635), .B2(w4610), .B1(w4629), .A1(w4628), .A2(w4634) );
	vdp_not g4661 (.nZ(w4632), .A(w4595) );
	vdp_not g4662 (.nZ(w4418), .A(w6320) );
	vdp_not g4663 (.nZ(w4419), .A(w4641) );
	vdp_not g4664 (.nZ(w4428), .A(w4645) );
	vdp_not g4665 (.nZ(w4422), .A(w4658) );
	vdp_not g4666 (.nZ(w4654), .A(w4650) );
	vdp_not g4667 (.nZ(w4421), .A(w4652) );
	vdp_dlatch_inv g4668 (.nQ(w4653), .D(w4650), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4669 (.nQ(w4652), .D(w4651), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g4670 (.nZ(w4420), .A(w4661) );
	vdp_dlatch_inv g4671 (.nQ(w4682), .D(w4616), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4672 (.nQ(w4661), .D(w4657), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g4673 (.nZ(w4662), .A(w4683) );
	vdp_dlatch_inv g4674 (.nQ(w4659), .D(w4683), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4675 (.nQ(w4672), .D(w4660), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g4676 (.nZ(w4656), .A(w4667) );
	vdp_dlatch_inv g4677 (.nQ(w4663), .D(w4667), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4678 (.nQ(w4673), .D(w4664), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4679 (.nQ(w4665), .D(w4655), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4680 (.nQ(w4670), .D(w4666), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4681 (.nQ(w4679), .D(w4668), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4682 (.nQ(w4681), .D(w4680), .nC(nHCLK2), .C(HCLK2) );
	vdp_sr_bit g4683 (.Q(w4414), .D(w6382), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4684 (.Z(w4668), .B2(w4610), .B1(1'b0), .A1(w4602), .A2(w4634) );
	vdp_aon22 g4685 (.Z(w4655), .B2(w4610), .B1(1'b0), .A1(w4612), .A2(w4634) );
	vdp_aon22 g4686 (.Z(w6382), .B2(w4708), .B1(M5), .A1(w120), .A2(w4746) );
	vdp_not g4687 (.nZ(w4698), .A(w1) );
	vdp_not g4688 (.nZ(w4749), .A(w4711) );
	vdp_not g4689 (.nZ(w4699), .A(w4710) );
	vdp_not g4690 (.nZ(w4747), .A(w4712) );
	vdp_not g4691 (.nZ(w4708), .A(w4709) );
	vdp_not g4692 (.nZ(w4746), .A(M5) );
	vdp_not g4693 (.nZ(w4703), .A(w4706) );
	vdp_not g4694 (.nZ(w4700), .A(w4414) );
	vdp_not g4695 (.nZ(w6391), .A(w4415) );
	vdp_not g4696 (.nZ(w4748), .A(M5) );
	vdp_not g4697 (.nZ(w4671), .A(w1) );
	vdp_not g4698 (.nZ(w4675), .A(w4607) );
	vdp_bufif0 g4699 (.A(1'b0), .Z(VRAMA[0]), .nE(w4504) );
	vdp_bufif0 g4700 (.A(w4492), .Z(VRAMA[1]), .nE(w4504) );
	vdp_bufif0 g4701 (.A(w4496), .Z(VRAMA[2]), .nE(w4504) );
	vdp_bufif0 g4702 (.A(w4499), .Z(VRAMA[3]), .nE(w4504) );
	vdp_bufif0 g4703 (.A(w4495), .Z(VRAMA[4]), .nE(w4504) );
	vdp_bufif0 g4704 (.A(w4493), .Z(VRAMA[5]), .nE(w4504) );
	vdp_bufif0 g4705 (.A(1'b0), .Z(VRAMA[6]), .nE(w4504) );
	vdp_bufif0 g4706 (.A(1'b0), .Z(VRAMA[7]), .nE(w4504) );
	vdp_aon22 g4707 (.Z(w4667), .B2(w4610), .B1(w6378), .A1(w4613), .A2(w4634) );
	vdp_aon22 g4708 (.Z(w4683), .B2(w4610), .B1(w4615), .A1(w4614), .A2(w4634) );
	vdp_aon22 g4709 (.Z(w4616), .B2(w4610), .B1(w4618), .A1(w4617), .A2(w4634) );
	vdp_comp_str g4710 (.A(w4631), .nZ(w4569), .Z(w4568) );
	vdp_and g4711 (.Z(w4594), .B(w4554), .A(w4550) );
	vdp_comp_we g4712 (.A(w4594), .nZ(w4634), .Z(w4610) );
	vdp_comp_str g4713 (.A(w4627), .nZ(w4584), .Z(w4583) );
	vdp_not g4714 (.nZ(w4550), .A(M5) );
	vdp_comp_str g4715 (.A(w4702), .nZ(w4713), .Z(w4705) );
	vdp_comp_str g4716 (.A(w4739), .nZ(w4721), .Z(w4726) );
	vdp_comp_we g4717 (.A(M5), .nZ(w4511), .Z(w4514) );
	vdp_comp_we g4718 (.A(w4545), .nZ(w4538), .Z(w4487) );
	vdp_comp_we g4719 (.A(w4525), .nZ(w4494), .Z(w4529) );
	vdp_comp_we g4720 (.A(M5), .nZ(w4501), .Z(w4497) );
	vdp_comp_we g4721 (.A(w1), .nZ(w4605), .Z(w4604) );
	vdp_comp_we g4722 (.nZ(w4720), .A(w4740), .Z(w4725) );
	vdp_and g4723 (.Z(w4631), .B(w4693), .A(DCLK2) );
	vdp_and g4724 (.Z(w4627), .B(w4695), .A(DCLK2) );
	vdp_and g4725 (.Z(w4692), .B(M5), .A(w4698) );
	vdp_and g4726 (.Z(w6394), .B(w4747), .A(M5) );
	vdp_and g4727 (.Z(w6393), .B(w4700), .A(w4415) );
	vdp_and g4728 (.Z(w4739), .B(w4738), .A(HCLK1) );
	vdp_or g4729 (.Z(w4674), .B(w4671), .A(w4681) );
	vdp_or g4730 (.Z(w6395), .B(w4748), .A(w4670) );
	vdp_and g4731 (.Z(w4489), .B(w4518), .A(w4502) );
	vdp_and g4732 (.Z(w4546), .B(w4483), .A(w4548) );
	vdp_and g4733 (.Z(w6183), .B(w4548), .A(w4484) );
	vdp_and g4734 (.Z(w6184), .B(w4482), .A(w4484) );
	vdp_and g4735 (.Z(w6185), .B(w4483), .A(w4482) );
	vdp_and g4736 (.Z(w6159), .B(H40), .A(VRAMA[9]) );
	vdp_or g4737 (.Z(w4556), .B(w4485), .A(w4554) );
	vdp_or g4738 (.Z(w4555), .B(w4485), .A(w4551) );
	vdp_not g4739 (.nZ(w4482), .A(w4548) );
	vdp_oai21 g4740 (.Z(w4509), .B(w28), .A1(w29), .A2(w5) );
	vdp_oai21 g4741 (.Z(w4706), .B(w4409), .A1(w4630), .A2(w4707) );
	vdp_aoi22 g4742 (.Z(w4595), .B2(w4550), .B1(w4551), .A1(M5), .A2(w4592) );
	vdp_or3 g4743 (.Z(w4592), .B(w4551), .A(w4552), .C(w4553) );
	vdp_and3 g4744 (.Z(w4702), .B(DCLK1), .A(HCLK2), .C(w4694) );
	vdp_oai21 g4745 (.Z(w4524), .B(M5), .A1(w4502), .A2(w4523) );
	vdp_2a3oi g4746 (.Z(w4516), .B(w4507), .A1(w4506), .A2(w4), .C(SYSRES) );
	vdp_or8 g4747 (.Z(w4707), .B(w4719), .A(M5), .C(w6325), .D(w4718), .F(w4716), .E(w4717), .G(w4715), .H(w4714) );
	vdp_and9 g4748 (.Z(w4376), .B(w4676), .A(w4678), .C(w4677), .D(w4675), .F(w4673), .E(w4674), .G(w4672), .H(w4669), .I(w6395) );
	vdp_nor12 g4749 (.Z(w4630), .B(w4616), .A(1'b0), .C(w4656), .D(M5), .F(w4668), .E(w4655), .G(w4662), .H(w4654), .J(w4637), .I(w4642), .K(w4635), .L(w4648) );
	vdp_or4 g4750 (.Z(w4545), .B(w4484), .A(w4483), .C(w4544), .D(w4486) );
	vdp_nand g4751 (.Z(w4633), .B(w4632), .A(HCLK1) );
	vdp_nand g4752 (.Z(w4678), .B(w4609), .A(w6392) );
	vdp_nand g4753 (.Z(w4677), .B(w4608), .A(w6391) );
	vdp_nor g4754 (.Z(w6392), .B(w4414), .A(w4415) );
	vdp_nand3 g4755 (.Z(w4676), .B(w4608), .A(w6393), .C(w4609) );
	vdp_sr_bit g4756 (.Q(w4417), .D(w4749), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4757 (.Q(w4757), .D(w26), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4758 (.Q(w4437), .D(w6315), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4759 (.Q(w4756), .D(w6299), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4760 (.Q(w6299), .D(w6300), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4761 (.Q(w6300), .D(w4755), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4762 (.Z(w4760), .B2(w4756), .B1(w5108), .A1(DB[4]), .A2(w5109) );
	vdp_notif0 g4763 (.A(HPOS[1]), .nZ(VRAMA[1]), .nE(w4971) );
	vdp_aon22 g4764 (.Z(w6315), .B2(w4754), .B1(w4757), .A1(M5), .A2(w26) );
	vdp_not g4765 (.nZ(w4754), .A(M5) );
	vdp_lfsr_bit g4766 (.Q(w4761), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6567), .A1(w4760), .A2(w6568) );
	vdp_lfsr_bit g4767 (.Q(w4764), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6565), .A1(w4761), .A2(w6566) );
	vdp_lfsr_bit g4768 (.Q(w4766), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6563), .A1(w4764), .A2(w6564) );
	vdp_lfsr_bit g4769 (.Q(w4767), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6561), .A1(w4766), .A2(w6562) );
	vdp_lfsr_bit g4770 (.Q(w4771), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6559), .A1(w4767), .A2(w6560) );
	vdp_lfsr_bit g4771 (.Q(w4769), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6557), .A1(w4771), .A2(w6558) );
	vdp_lfsr_bit g4772 (.Q(w4773), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6555), .A1(w4769), .A2(w6556) );
	vdp_lfsr_bit g4773 (.Q(w4753), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6554), .A1(w4773), .A2(w6553) );
	vdp_lfsr_bit g4774 (.Q(w4777), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4951), .A1(w4753), .A2(w6552) );
	vdp_lfsr_bit g4775 (.Q(w4779), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5112), .A1(w4777), .A2(w5113) );
	vdp_lfsr_bit g4776 (.Q(w4783), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4997), .A1(w4779), .A2(w4998) );
	vdp_lfsr_bit g4777 (.Q(w4780), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4994), .A1(w4783), .A2(w4995) );
	vdp_lfsr_bit g4778 (.Q(w4782), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4992), .A1(w4780), .A2(w4993) );
	vdp_lfsr_bit g4779 (.Q(w4786), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6550), .A1(w4782), .A2(w6549) );
	vdp_lfsr_bit g4780 (.Q(w4787), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4989), .A1(w4786), .A2(w4990) );
	vdp_lfsr_bit g4781 (.Q(w4791), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6547), .A1(w4787), .A2(w6548) );
	vdp_lfsr_bit g4782 (.Q(w4790), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6551), .A1(w4791), .A2(w6318) );
	vdp_lfsr_bit g4783 (.Q(w4795), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4986), .A1(w4790), .A2(w4987) );
	vdp_lfsr_bit g4784 (.Q(w4797), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4985), .A1(w4795), .A2(w4984) );
	vdp_lfsr_bit g4785 (.Q(w4752), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4982), .A1(w4797), .A2(w4983) );
	vdp_bufif0 g4786 (.A(w4753), .Z(VRAMA[1]), .nE(w6317) );
	vdp_bufif0 g4787 (.A(1'b0), .Z(VRAMA[1]), .nE(w5005) );
	vdp_notif0 g4788 (.A(w4752), .nZ(DB[4]), .nE(w5114) );
	vdp_sr_bit g4789 (.Q(w4802), .D(w6302), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4790 (.Q(w6302), .D(w6301), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4791 (.Q(w6301), .D(w6167), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4792 (.Z(w4759), .B2(w4802), .B1(w5108), .A1(DB[5]), .A2(w5109) );
	vdp_notif0 g4793 (.A(w4810), .nZ(VRAMA[2]), .nE(w4971) );
	vdp_lfsr_bit g4794 (.Q(w4762), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6567), .A1(w4759), .A2(w6568) );
	vdp_lfsr_bit g4795 (.Q(w4763), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6565), .A1(w4762), .A2(w6566) );
	vdp_lfsr_bit g4796 (.Q(w4765), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6563), .A1(w4763), .A2(w6564) );
	vdp_lfsr_bit g4797 (.Q(w4768), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6561), .A1(w4765), .A2(w6562) );
	vdp_lfsr_bit g4798 (.Q(w4772), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6559), .A1(w4768), .A2(w6560) );
	vdp_lfsr_bit g4799 (.Q(w4770), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6557), .A1(w4772), .A2(w6558) );
	vdp_lfsr_bit g4800 (.Q(w4774), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6555), .A1(w4770), .A2(w6556) );
	vdp_lfsr_bit g4801 (.Q(w4775), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6554), .A1(w4774), .A2(w6553) );
	vdp_lfsr_bit g4802 (.Q(w4778), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4951), .A1(w4775), .A2(w6552) );
	vdp_lfsr_bit g4803 (.Q(w4776), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5112), .A1(w4778), .A2(w5113) );
	vdp_lfsr_bit g4804 (.Q(w4784), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4997), .A1(w4776), .A2(w4998) );
	vdp_lfsr_bit g4805 (.Q(w4781), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4994), .A1(w4784), .A2(w4995) );
	vdp_lfsr_bit g4806 (.Q(w4785), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4992), .A1(w4781), .A2(w4993) );
	vdp_lfsr_bit g4807 (.Q(w4789), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6550), .A1(w4785), .A2(w6549) );
	vdp_lfsr_bit g4808 (.Q(w4788), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4989), .A1(w4789), .A2(w4990) );
	vdp_lfsr_bit g4809 (.Q(w4792), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6547), .A1(w4788), .A2(w6548) );
	vdp_lfsr_bit g4810 (.Q(w4793), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6551), .A1(w4792), .A2(w6318) );
	vdp_lfsr_bit g4811 (.Q(w4794), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4986), .A1(w4793), .A2(w4987) );
	vdp_lfsr_bit g4812 (.Q(w4798), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4985), .A1(w4794), .A2(w4984) );
	vdp_lfsr_bit g4813 (.Q(w4800), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4982), .A1(w4798), .A2(w4983) );
	vdp_bufif0 g4814 (.A(w4775), .Z(VRAMA[2]), .nE(w6317) );
	vdp_bufif0 g4815 (.A(1'b1), .Z(VRAMA[2]), .nE(w5005) );
	vdp_notif0 g4816 (.A(w4800), .nZ(DB[5]), .nE(w5114) );
	vdp_aon22 g4817 (.Z(w4799), .B2(w4791), .B1(w4979), .A1(w4978), .A2(w4752) );
	vdp_dlatch_inv g4818 (.nQ(w4811), .D(w4804), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g4819 (.nQ(w4806), .D(w4758), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g4820 (.Z(w4805), .B(w4806), .A(DCLK2) );
	vdp_nand g4821 (.Z(w4804), .B(HCLK1), .A(w4437) );
	vdp_nand g4822 (.Z(w4758), .B(HCLK1), .A(w26) );
	vdp_sr_bit g4823 (.Q(w4803), .D(w6304), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4824 (.Q(w6304), .D(w6303), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4825 (.Q(w6303), .D(w4808), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4826 (.Z(w4819), .B2(w4803), .B1(w5108), .A1(DB[6]), .A2(w5109) );
	vdp_notif0 g4827 (.A(w4817), .nZ(VRAMA[3]), .nE(w4971) );
	vdp_lfsr_bit g4828 (.Q(w4821), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6567), .A1(w4819), .A2(w6568) );
	vdp_lfsr_bit g4829 (.Q(w4822), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6565), .A1(w4821), .A2(w6566) );
	vdp_lfsr_bit g4830 (.Q(w4825), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6563), .A1(w4822), .A2(w6564) );
	vdp_lfsr_bit g4831 (.Q(w4826), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6561), .A1(w4825), .A2(w6562) );
	vdp_lfsr_bit g4832 (.Q(w4831), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6559), .A1(w4826), .A2(w6560) );
	vdp_lfsr_bit g4833 (.Q(w4830), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6557), .A1(w4831), .A2(w6558) );
	vdp_lfsr_bit g4834 (.Q(w4833), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6555), .A1(w4830), .A2(w6556) );
	vdp_lfsr_bit g4835 (.Q(w4835), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6554), .A1(w4833), .A2(w6553) );
	vdp_lfsr_bit g4836 (.Q(w4837), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4951), .A1(w4835), .A2(w6552) );
	vdp_lfsr_bit g4837 (.Q(w4839), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5112), .A1(w4837), .A2(w5113) );
	vdp_lfsr_bit g4838 (.Q(w4841), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4997), .A1(w4839), .A2(w4998) );
	vdp_lfsr_bit g4839 (.Q(w4843), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4994), .A1(w4841), .A2(w4995) );
	vdp_lfsr_bit g4840 (.Q(w4845), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4992), .A1(w4843), .A2(w4993) );
	vdp_lfsr_bit g4841 (.Q(w4848), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6550), .A1(w4845), .A2(w6549) );
	vdp_lfsr_bit g4842 (.Q(w4849), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4989), .A1(w4848), .A2(w4990) );
	vdp_lfsr_bit g4843 (.Q(w4850), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6547), .A1(w4849), .A2(w6548) );
	vdp_lfsr_bit g4844 (.Q(w4855), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6551), .A1(w4850), .A2(w6318) );
	vdp_lfsr_bit g4845 (.Q(w4854), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4986), .A1(w4855), .A2(w4987) );
	vdp_lfsr_bit g4846 (.Q(w4857), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4985), .A1(w4854), .A2(w4984) );
	vdp_lfsr_bit g4847 (.Q(w4801), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4982), .A1(w4857), .A2(w4983) );
	vdp_bufif0 g4848 (.A(w4835), .Z(VRAMA[3]), .nE(w6317) );
	vdp_bufif0 g4849 (.A(w4799), .Z(VRAMA[3]), .nE(w5005) );
	vdp_notif0 g4850 (.A(w4801), .nZ(DB[6]), .nE(w5114) );
	vdp_aon22 g4851 (.Z(w4858), .B2(w4792), .B1(w4979), .A1(w4978), .A2(w4800) );
	vdp_sr_bit g4852 (.Q(w4813), .D(w4811), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g4853 (.Q(w4807), .D(w4806), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_and g4854 (.Z(w4809), .B(w4811), .A(DCLK2) );
	vdp_and g4855 (.Z(w4815), .B(DCLK2), .A(w4813) );
	vdp_and g4856 (.Z(w4812), .B(w4807), .A(DCLK2) );
	vdp_sr_bit g4857 (.Q(w4870), .D(w6305), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4858 (.Q(w6305), .D(w6306), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4859 (.Q(w6306), .D(w4814), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4860 (.Z(w4818), .B2(w4870), .B1(w5108), .A1(DB[7]), .A2(w5109) );
	vdp_notif0 g4861 (.A(w4868), .nZ(VRAMA[4]), .nE(w4971) );
	vdp_lfsr_bit g4862 (.Q(w4820), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6567), .A1(w4818), .A2(w6568) );
	vdp_lfsr_bit g4863 (.Q(w4823), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6565), .A1(w4820), .A2(w6566) );
	vdp_lfsr_bit g4864 (.Q(w4824), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6563), .A1(w4823), .A2(w6564) );
	vdp_lfsr_bit g4865 (.Q(w4827), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6561), .A1(w4824), .A2(w6562) );
	vdp_lfsr_bit g4866 (.Q(w4828), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6559), .A1(w4827), .A2(w6560) );
	vdp_lfsr_bit g4867 (.Q(w4829), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6557), .A1(w4828), .A2(w6558) );
	vdp_lfsr_bit g4868 (.Q(w4832), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6555), .A1(w4829), .A2(w6556) );
	vdp_lfsr_bit g4869 (.Q(w4834), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6554), .A1(w4832), .A2(w6553) );
	vdp_lfsr_bit g4870 (.Q(w4836), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4951), .A1(w4834), .A2(w6552) );
	vdp_lfsr_bit g4871 (.Q(w4838), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5112), .A1(w4836), .A2(w5113) );
	vdp_lfsr_bit g4872 (.Q(w4840), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4997), .A1(w4838), .A2(w4998) );
	vdp_lfsr_bit g4873 (.Q(w4842), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4994), .A1(w4840), .A2(w4995) );
	vdp_lfsr_bit g4874 (.Q(w4844), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4992), .A1(w4842), .A2(w4993) );
	vdp_lfsr_bit g4875 (.Q(w4847), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6550), .A1(w4844), .A2(w6549) );
	vdp_lfsr_bit g4876 (.Q(w4846), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4989), .A1(w4847), .A2(w4990) );
	vdp_lfsr_bit g4877 (.Q(w4851), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6547), .A1(w4846), .A2(w6548) );
	vdp_lfsr_bit g4878 (.Q(w4852), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6551), .A1(w4851), .A2(w6318) );
	vdp_lfsr_bit g4879 (.Q(w4853), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4986), .A1(w4852), .A2(w4987) );
	vdp_lfsr_bit g4880 (.Q(w4856), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4985), .A1(w4853), .A2(w4984) );
	vdp_lfsr_bit g4881 (.Q(w4872), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4982), .A1(w4856), .A2(w4983) );
	vdp_bufif0 g4882 (.A(w4834), .Z(VRAMA[4]), .nE(w6317) );
	vdp_bufif0 g4883 (.A(w4858), .Z(VRAMA[4]), .nE(w5005) );
	vdp_notif0 g4884 (.A(w4872), .nZ(DB[7]), .nE(w5114) );
	vdp_aon22 g4885 (.Z(w4873), .B2(w4850), .B1(w4979), .A1(w4978), .A2(w4801) );
	vdp_aon22 g4886 (.Z(w4867), .B2(w4860), .B1(w120), .A1(w4816), .A2(w4866) );
	vdp_not g4887 (.nZ(w4816), .A(w120) );
	vdp_comp_str g4888 (.nZ(w4861), .A(w4812), .Z(w4862) );
	vdp_comp_str g4889 (.nZ(w4865), .A(w4815), .Z(w4864) );
	vdp_sr_bit g4890 (.Q(w4869), .D(w6308), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4891 (.Q(w6308), .D(w6307), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4892 (.Q(w6307), .D(w4863), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4893 (.Z(w4913), .B2(w4869), .B1(w5108), .A1(DB[8]), .A2(w5109) );
	vdp_notif0 g4894 (.A(w4867), .nZ(VRAMA[5]), .nE(w4971) );
	vdp_lfsr_bit g4895 (.Q(w4911), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6567), .A1(w4913), .A2(w6568) );
	vdp_lfsr_bit g4896 (.Q(w4908), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6565), .A1(w4911), .A2(w6566) );
	vdp_lfsr_bit g4897 (.Q(w4907), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6563), .A1(w4908), .A2(w6564) );
	vdp_lfsr_bit g4898 (.Q(w4904), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6561), .A1(w4907), .A2(w6562) );
	vdp_lfsr_bit g4899 (.Q(w4903), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6559), .A1(w4904), .A2(w6560) );
	vdp_lfsr_bit g4900 (.Q(w4900), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6557), .A1(w4903), .A2(w6558) );
	vdp_lfsr_bit g4901 (.Q(w4899), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6555), .A1(w4900), .A2(w6556) );
	vdp_lfsr_bit g4902 (.Q(w4877), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6554), .A1(w4899), .A2(w6553) );
	vdp_lfsr_bit g4903 (.Q(w4896), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4951), .A1(w4877), .A2(w6552) );
	vdp_lfsr_bit g4904 (.Q(w4871), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5112), .A1(w4896), .A2(w5113) );
	vdp_lfsr_bit g4905 (.Q(w4893), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4997), .A1(w4871), .A2(w4998) );
	vdp_lfsr_bit g4906 (.Q(w4892), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4994), .A1(w4893), .A2(w4995) );
	vdp_lfsr_bit g4907 (.Q(w4889), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4992), .A1(w4892), .A2(w4993) );
	vdp_lfsr_bit g4908 (.Q(w4887), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6550), .A1(w4889), .A2(w6549) );
	vdp_lfsr_bit g4909 (.Q(w4886), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4989), .A1(w4887), .A2(w4990) );
	vdp_lfsr_bit g4910 (.Q(w4875), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6547), .A1(w4886), .A2(w6548) );
	vdp_lfsr_bit g4911 (.Q(w4882), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6551), .A1(w4875), .A2(w6318) );
	vdp_lfsr_bit g4912 (.Q(w4880), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4986), .A1(w4882), .A2(w4987) );
	vdp_lfsr_bit g4913 (.Q(w4878), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4985), .A1(w4880), .A2(w4984) );
	vdp_lfsr_bit g4914 (.Q(w4895), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4982), .A1(w4878), .A2(w4983) );
	vdp_bufif0 g4915 (.A(w4877), .Z(VRAMA[5]), .nE(w6317) );
	vdp_bufif0 g4916 (.A(w4873), .Z(VRAMA[5]), .nE(w5005) );
	vdp_notif0 g4917 (.A(w4895), .nZ(DB[8]), .nE(w5114) );
	vdp_aon22 g4918 (.Z(w4874), .B2(w4851), .B1(w4979), .A1(w4978), .A2(w4872) );
	vdp_slatch g4919 (.D(S[0]), .nC(w4865), .C(w4864), .Q(w4918) );
	vdp_slatch g4920 (.D(S[0]), .nC(w4861), .C(w4862), .Q(w4859) );
	vdp_aoi22 g4921 (.Z(w4866), .B2(w4917), .B1(w4918), .A1(w4916), .A2(w4859) );
	vdp_sr_bit g4922 (.Q(w4925), .D(w6310), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4923 (.Q(w6310), .D(w6309), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4924 (.Q(w6309), .D(w4914), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4925 (.Z(w4912), .B2(w4925), .B1(w5108), .A1(DB[9]), .A2(w5109) );
	vdp_notif0 g4926 (.A(w4915), .nZ(VRAMA[6]), .nE(w4971) );
	vdp_lfsr_bit g4927 (.Q(w4910), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6567), .A1(w4912), .A2(w6568) );
	vdp_lfsr_bit g4928 (.Q(w4909), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6565), .A1(w4910), .A2(w6566) );
	vdp_lfsr_bit g4929 (.Q(w4906), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6563), .A1(w4909), .A2(w6564) );
	vdp_lfsr_bit g4930 (.Q(w4905), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6561), .A1(w4906), .A2(w6562) );
	vdp_lfsr_bit g4931 (.Q(w4902), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6559), .A1(w4905), .A2(w6560) );
	vdp_lfsr_bit g4932 (.Q(w4901), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6557), .A1(w4902), .A2(w6558) );
	vdp_lfsr_bit g4933 (.Q(w4898), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6555), .A1(w4901), .A2(w6556) );
	vdp_lfsr_bit g4934 (.Q(w4876), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6554), .A1(w4898), .A2(w6553) );
	vdp_lfsr_bit g4935 (.Q(w4897), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4951), .A1(w4876), .A2(w6552) );
	vdp_lfsr_bit g4936 (.Q(w4923), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5112), .A1(w4897), .A2(w5113) );
	vdp_lfsr_bit g4937 (.Q(w4894), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4997), .A1(w4923), .A2(w4998) );
	vdp_lfsr_bit g4938 (.Q(w4891), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4994), .A1(w4894), .A2(w4995) );
	vdp_lfsr_bit g4939 (.Q(w4890), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4992), .A1(w4891), .A2(w4993) );
	vdp_lfsr_bit g4940 (.Q(w4888), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6550), .A1(w4890), .A2(w6549) );
	vdp_lfsr_bit g4941 (.Q(w4885), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4989), .A1(w4888), .A2(w4990) );
	vdp_lfsr_bit g4942 (.Q(w4884), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6547), .A1(w4885), .A2(w6548) );
	vdp_lfsr_bit g4943 (.Q(w4883), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6551), .A1(w4884), .A2(w6318) );
	vdp_lfsr_bit g4944 (.Q(w4881), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4986), .A1(w4883), .A2(w4987) );
	vdp_lfsr_bit g4945 (.Q(w4879), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4985), .A1(w4881), .A2(w4984) );
	vdp_lfsr_bit g4946 (.Q(w4920), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4982), .A1(w4879), .A2(w4983) );
	vdp_bufif0 g4947 (.A(w4876), .Z(VRAMA[6]), .nE(w6317) );
	vdp_bufif0 g4948 (.A(w4874), .Z(VRAMA[6]), .nE(w5005) );
	vdp_notif0 g4949 (.A(w4920), .nZ(DB[9]), .nE(w5114) );
	vdp_aon22 g4950 (.Z(w4922), .B2(w4875), .B1(w4979), .A1(w4978), .A2(w4895) );
	vdp_aoi22 g4951 (.Z(w4915), .B2(w4917), .B1(w4927), .A1(w4916), .A2(w4919) );
	vdp_slatch g4952 (.D(S[1]), .nC(w4865), .C(w4864), .Q(w4927) );
	vdp_slatch g4953 (.D(S[1]), .nC(w4861), .C(w4862), .Q(w4919) );
	vdp_sr_bit g4954 (.Q(w4924), .D(w6312), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4955 (.Q(w6312), .D(w6311), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4956 (.Q(w6311), .D(w4928), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4957 (.Z(w4970), .B2(w4924), .B1(w5108), .A1(DB[10]), .A2(w5109) );
	vdp_notif0 g4958 (.A(w4973), .nZ(VRAMA[7]), .nE(w4974) );
	vdp_lfsr_bit g4959 (.Q(w4969), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6567), .A1(w4970), .A2(w6568) );
	vdp_lfsr_bit g4960 (.Q(w4964), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6565), .A1(w4969), .A2(w6566) );
	vdp_lfsr_bit g4961 (.Q(w4965), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6563), .A1(w4964), .A2(w6564) );
	vdp_lfsr_bit g4962 (.Q(w4959), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6561), .A1(w4965), .A2(w6562) );
	vdp_lfsr_bit g4963 (.Q(w4960), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6559), .A1(w4959), .A2(w6560) );
	vdp_lfsr_bit g4964 (.Q(w4957), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6557), .A1(w4960), .A2(w6558) );
	vdp_lfsr_bit g4965 (.Q(w4955), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6555), .A1(w4957), .A2(w6556) );
	vdp_lfsr_bit g4966 (.Q(w4921), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6554), .A1(w4955), .A2(w6553) );
	vdp_lfsr_bit g4967 (.Q(w4952), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4951), .A1(w4921), .A2(w6552) );
	vdp_lfsr_bit g4968 (.Q(w4947), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5112), .A1(w4952), .A2(w5113) );
	vdp_lfsr_bit g4969 (.Q(w4949), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4997), .A1(w4947), .A2(w4998) );
	vdp_lfsr_bit g4970 (.Q(w4946), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4994), .A1(w4949), .A2(w4995) );
	vdp_lfsr_bit g4971 (.Q(w4945), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4992), .A1(w4946), .A2(w4993) );
	vdp_lfsr_bit g4972 (.Q(w4942), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6550), .A1(w4945), .A2(w6549) );
	vdp_lfsr_bit g4973 (.Q(w4940), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4989), .A1(w4942), .A2(w4990) );
	vdp_lfsr_bit g4974 (.Q(w4938), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6547), .A1(w4940), .A2(w6548) );
	vdp_lfsr_bit g4975 (.Q(w4936), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6551), .A1(w4938), .A2(w6318) );
	vdp_lfsr_bit g4976 (.Q(w4934), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4986), .A1(w4936), .A2(w4987) );
	vdp_lfsr_bit g4977 (.Q(w4932), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4985), .A1(w4934), .A2(w4984) );
	vdp_lfsr_bit g4978 (.Q(w4930), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4982), .A1(w4932), .A2(w4983) );
	vdp_bufif0 g4979 (.A(w4921), .Z(VRAMA[7]), .nE(w6317) );
	vdp_bufif0 g4980 (.A(w4922), .Z(VRAMA[7]), .nE(w5005) );
	vdp_notif0 g4981 (.A(w4930), .nZ(DB[10]), .nE(w5114) );
	vdp_aon22 g4982 (.Z(w4929), .B2(w4884), .B1(w4979), .A1(w4978), .A2(w4920) );
	vdp_aoi22 g4983 (.Z(w4973), .B2(w4917), .B1(w4975), .A1(w4916), .A2(w4926) );
	vdp_slatch g4984 (.D(S[2]), .nC(w4865), .C(w4864), .Q(w4975) );
	vdp_slatch g4985 (.D(S[2]), .nC(w4861), .C(w4862), .Q(w4926) );
	vdp_sr_bit g4986 (.Q(w5000), .D(w27), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4987 (.Q(w4999), .D(w21), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4988 (.Z(w4967), .B2(w4412), .B1(w5108), .A1(DB[11]), .A2(w5109) );
	vdp_notif0 g4989 (.A(w4972), .nZ(VRAMA[8]), .nE(w4974) );
	vdp_lfsr_bit g4990 (.Q(w4968), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6567), .A1(w4967), .A2(w6568) );
	vdp_lfsr_bit g4991 (.Q(w4963), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6565), .A1(w4968), .A2(w6566) );
	vdp_lfsr_bit g4992 (.Q(w4966), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6563), .A1(w4963), .A2(w6564) );
	vdp_lfsr_bit g4993 (.Q(w4962), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6561), .A1(w4966), .A2(w6562) );
	vdp_lfsr_bit g4994 (.Q(w4961), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6559), .A1(w4962), .A2(w6560) );
	vdp_lfsr_bit g4995 (.Q(w4958), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6557), .A1(w4961), .A2(w6558) );
	vdp_lfsr_bit g4996 (.Q(w4956), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6555), .A1(w4958), .A2(w6556) );
	vdp_lfsr_bit g4997 (.Q(w4954), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6554), .A1(w4956), .A2(w6553) );
	vdp_lfsr_bit g4998 (.Q(w4953), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4951), .A1(w4954), .A2(w6552) );
	vdp_lfsr_bit g4999 (.Q(w4950), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5112), .A1(w4953), .A2(w5113) );
	vdp_lfsr_bit g5000 (.Q(w4948), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4997), .A1(w4950), .A2(w4998) );
	vdp_lfsr_bit g5001 (.Q(w4944), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4994), .A1(w4948), .A2(w4995) );
	vdp_lfsr_bit g5002 (.Q(w4943), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4992), .A1(w4944), .A2(w4993) );
	vdp_lfsr_bit g5003 (.Q(w4941), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6550), .A1(w4943), .A2(w6549) );
	vdp_lfsr_bit g5004 (.Q(w4939), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4989), .A1(w4941), .A2(w4990) );
	vdp_lfsr_bit g5005 (.Q(w4937), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6547), .A1(w4939), .A2(w6548) );
	vdp_lfsr_bit g5006 (.Q(w4935), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6551), .A1(w4937), .A2(w6318) );
	vdp_lfsr_bit g5007 (.Q(w4933), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4986), .A1(w4935), .A2(w4987) );
	vdp_lfsr_bit g5008 (.Q(w4931), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4985), .A1(w4933), .A2(w4984) );
	vdp_lfsr_bit g5009 (.Q(w4996), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4982), .A1(w4931), .A2(w4983) );
	vdp_bufif0 g5010 (.A(1'b0), .Z(VRAMA[0]), .nE(w6317) );
	vdp_bufif0 g5011 (.A(w4929), .Z(VRAMA[8]), .nE(w5005) );
	vdp_notif0 g5012 (.A(w4996), .nZ(DB[11]), .nE(w5114) );
	vdp_aon22 g5013 (.Z(w5006), .B2(w4980), .B1(w4979), .A1(w4978), .A2(w4930) );
	vdp_aoi22 g5014 (.Z(w4972), .B2(w4917), .B1(w4976), .A1(w4916), .A2(w4977) );
	vdp_slatch g5015 (.D(S[3]), .nC(w4865), .C(w4864), .Q(w4976) );
	vdp_slatch g5016 (.D(S[3]), .nC(w4861), .C(w4862), .Q(w4977) );
	vdp_bufif0 g5017 (.A(1'b0), .Z(VRAMA[0]), .nE(w5005) );
	vdp_bufif0 g5018 (.A(w5008), .Z(VRAMA[8]), .nE(w5012) );
	vdp_aon22 g5019 (.Z(w5035), .B2(w4422), .B1(w5108), .A1(DB[3]), .A2(w5109) );
	vdp_lfsr_bit g5020 (.Q(w5033), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6567), .A1(w5035), .A2(w6568) );
	vdp_lfsr_bit g5021 (.Q(w5031), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6565), .A1(w5033), .A2(w6566) );
	vdp_lfsr_bit g5022 (.Q(w5029), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6563), .A1(w5031), .A2(w6564) );
	vdp_lfsr_bit g5023 (.Q(w5027), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6561), .A1(w5029), .A2(w6562) );
	vdp_lfsr_bit g5024 (.Q(w5024), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6559), .A1(w5027), .A2(w6560) );
	vdp_lfsr_bit g5025 (.Q(w5023), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6557), .A1(w5024), .A2(w6558) );
	vdp_lfsr_bit g5026 (.Q(w5021), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6555), .A1(w5023), .A2(w6556) );
	vdp_lfsr_bit g5027 (.Q(w5019), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6554), .A1(w5021), .A2(w6553) );
	vdp_lfsr_bit g5028 (.Q(w5004), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4951), .A1(w5019), .A2(w6552) );
	vdp_lfsr_bit g5029 (.Q(w5002), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5112), .A1(w5004), .A2(w5113) );
	vdp_notif0 g5030 (.A(w5002), .nZ(DB[3]), .nE(w5114) );
	vdp_not g5031 (.nZ(w4991), .A(M5) );
	vdp_not g5032 (.nZ(w5001), .A(H40) );
	vdp_notif0 g5033 (.A(1'b1), .nZ(VRAMA[0]), .nE(w4971) );
	vdp_aoi22 g5034 (.Z(w4860), .B2(w5039), .B1(w5004), .A1(w4916), .A2(w5002) );
	vdp_not g5035 (.nZ(w5037), .A(M5) );
	vdp_or g5036 (.Z(w5038), .B(w5000), .A(w4999) );
	vdp_sr_bit g5037 (.Q(w5009), .D(w8), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5038 (.Q(w5015), .D(w28), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_comp_we g5039 (.nZ(w4982), .A(w5007), .Z(w4983) );
	vdp_comp_we g5040 (.nZ(w4985), .A(w5007), .Z(w4984) );
	vdp_comp_we g5041 (.nZ(w4986), .A(w5007), .Z(w4987) );
	vdp_comp_we g5042 (.nZ(w6551), .A(w5007), .Z(w6318) );
	vdp_comp_we g5043 (.nZ(w6547), .A(w5007), .Z(w6548) );
	vdp_comp_we g5044 (.nZ(w4979), .A(H40), .Z(w4978) );
	vdp_comp_we g5045 (.nZ(w4989), .A(w5007), .Z(w4990) );
	vdp_comp_we g5046 (.nZ(w6550), .A(w5007), .Z(w6549) );
	vdp_comp_we g5047 (.nZ(w4992), .A(w5007), .Z(w4993) );
	vdp_comp_we g5048 (.nZ(w4994), .A(w5007), .Z(w4995) );
	vdp_comp_we g5049 (.nZ(w4997), .A(w5007), .Z(w4998) );
	vdp_comp_we g5050 (.nZ(w4917), .A(w4999), .Z(w4916) );
	vdp_not g5051 (.nZ(w4974), .A(w5003) );
	vdp_not g5052 (.nZ(w4971), .A(w5003) );
	vdp_not g5053 (.nZ(w5005), .A(w5011) );
	vdp_not g5054 (.nZ(w6317), .A(w4988) );
	vdp_and g5055 (.Z(w4988), .B(w5009), .A(w4991) );
	vdp_oai21 g5056 (.Z(w5014), .B(w4991), .A1(w5015), .A2(w5009) );
	vdp_aon333 g5057 (.Z(w4375), .B1(M5), .A1(1'b1), .C1(M5), .A2(w4991), .A3(w4954), .B2(w4937), .B3(w5001), .C2(H40), .C3(w4996) );
	vdp_aon22 g5058 (.Z(w5034), .B2(w4428), .B1(w5108), .A1(DB[2]), .A2(w5109) );
	vdp_lfsr_bit g5059 (.Q(w5032), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6567), .A1(w5034), .A2(w6568) );
	vdp_lfsr_bit g5060 (.Q(w5030), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6565), .A1(w5032), .A2(w6566) );
	vdp_lfsr_bit g5061 (.Q(w5028), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6563), .A1(w5030), .A2(w6564) );
	vdp_lfsr_bit g5062 (.Q(w5026), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6561), .A1(w5028), .A2(w6562) );
	vdp_lfsr_bit g5063 (.Q(w5025), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6559), .A1(w5026), .A2(w6560) );
	vdp_lfsr_bit g5064 (.Q(w5022), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6557), .A1(w5025), .A2(w6558) );
	vdp_lfsr_bit g5065 (.Q(w5020), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6555), .A1(w5022), .A2(w6556) );
	vdp_lfsr_bit g5066 (.Q(w5018), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6554), .A1(w5020), .A2(w6553) );
	vdp_lfsr_bit g5067 (.Q(w5017), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4951), .A1(w5018), .A2(w6552) );
	vdp_lfsr_bit g5068 (.Q(w5016), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5112), .A1(w5017), .A2(w5113) );
	vdp_notif0 g5069 (.A(w5016), .nZ(DB[2]), .nE(w5114) );
	vdp_aoi22 g5070 (.Z(w4868), .B2(w5039), .B1(w5017), .A1(w4916), .A2(w5016) );
	vdp_aoi22 g5071 (.Z(w5051), .B2(w5039), .B1(w5052), .A1(w4916), .A2(w4377) );
	vdp_notif0 g5072 (.A(w5051), .nZ(VRAMA[9]), .nE(w4974) );
	vdp_slatch g5074 (.D(S[4]), .nC(w4862), .C(w4861), .Q(w4377) );
	vdp_and g5075 (.Z(w5003), .B(w5037), .A(w5038) );
	vdp_slatch g5076 (.D(REG_BUS[0]), .nC(w5111), .C(w5110), .Q(w4980) );
	vdp_slatch g5077 (.D(REG_BUS[7]), .nC(w5111), .C(w5110), .Q(w5010) );
	vdp_bufif0 g5078 (.A(w5006), .Z(VRAMA[9]), .nE(w5041) );
	vdp_bufif0 g5079 (.A(w5010), .Z(VRAMA[16]), .nE(w5041) );
	vdp_and g5080 (.Z(w5011), .B(w5009), .A(M5) );
	vdp_not g5081 (.nZ(w5041), .A(w5011) );
	vdp_not g5082 (.nZ(w5012), .A(w5013) );
	vdp_not g5083 (.nZ(w5013), .A(w5014) );
	vdp_xor g5084 (.Z(w5040), .B(w5010), .A(VRAMA[16]) );
	vdp_xor g5085 (.Z(w5044), .B(w5046), .A(w5045) );
	vdp_and3 g5086 (.Z(w6165), .B(w5050), .A(w5047), .C(M5) );
	vdp_nor g5087 (.Z(w5046), .B(H40), .A(w4980) );
	vdp_nor g5088 (.Z(w5045), .B(H40), .A(VRAMA[9]) );
	vdp_aon22 g5089 (.Z(w5070), .B2(w4419), .B1(w5108), .A1(DB[1]), .A2(w5109) );
	vdp_lfsr_bit g5090 (.Q(w5069), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6567), .A1(w5070), .A2(w6568) );
	vdp_lfsr_bit g5091 (.Q(w5068), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6565), .A1(w5069), .A2(w6566) );
	vdp_lfsr_bit g5092 (.Q(w5067), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6563), .A1(w5068), .A2(w6564) );
	vdp_lfsr_bit g5093 (.Q(w5066), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6561), .A1(w5067), .A2(w6562) );
	vdp_lfsr_bit g5094 (.Q(w5065), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6559), .A1(w5066), .A2(w6560) );
	vdp_lfsr_bit g5095 (.Q(w5064), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6557), .A1(w5065), .A2(w6558) );
	vdp_lfsr_bit g5096 (.Q(w5063), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6555), .A1(w5064), .A2(w6556) );
	vdp_lfsr_bit g5097 (.Q(w5062), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6554), .A1(w5063), .A2(w6553) );
	vdp_lfsr_bit g5098 (.Q(w5049), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4951), .A1(w5062), .A2(w6552) );
	vdp_lfsr_bit g5099 (.Q(w5060), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5112), .A1(w5049), .A2(w5113) );
	vdp_notif0 g5100 (.A(w5060), .nZ(DB[1]), .nE(w5114) );
	vdp_slatch g5101 (.D(REG_BUS[1]), .nC(w5111), .C(w5110), .Q(w5008) );
	vdp_slatch g5102 (.D(REG_BUS[6]), .nC(w5111), .C(w5110), .Q(w5059) );
	vdp_xor g5103 (.Z(w5043), .B(w5059), .A(VRAMA[15]) );
	vdp_xor g5104 (.Z(w5042), .B(w5008), .A(VRAMA[10]) );
	vdp_aon22 g5105 (.Z(w5079), .B2(w4418), .B1(w5108), .A1(DB[0]), .A2(w5109) );
	vdp_lfsr_bit g5106 (.Q(w5080), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6567), .A1(w5079), .A2(w6568) );
	vdp_lfsr_bit g5107 (.Q(w5081), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6565), .A1(w5080), .A2(w6566) );
	vdp_lfsr_bit g5108 (.Q(w5082), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6563), .A1(w5081), .A2(w6564) );
	vdp_lfsr_bit g5109 (.Q(w5084), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6561), .A1(w5082), .A2(w6562) );
	vdp_lfsr_bit g5110 (.Q(w5083), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6559), .A1(w5084), .A2(w6560) );
	vdp_lfsr_bit g5111 (.Q(w5086), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6557), .A1(w5083), .A2(w6558) );
	vdp_lfsr_bit g5112 (.Q(w5085), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6555), .A1(w5086), .A2(w6556) );
	vdp_lfsr_bit g5113 (.Q(w5087), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6554), .A1(w5085), .A2(w6553) );
	vdp_lfsr_bit g5114 (.Q(w5061), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4951), .A1(w5087), .A2(w6552) );
	vdp_lfsr_bit g5115 (.Q(w6316), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5112), .A1(w5061), .A2(w5113) );
	vdp_notif0 g5116 (.A(w6316), .nZ(DB[0]), .nE(w5114) );
	vdp_slatch g5117 (.D(REG_BUS[2]), .nC(w5111), .C(w5110), .Q(w5058) );
	vdp_slatch g5118 (.D(REG_BUS[5]), .nC(w5111), .C(w5110), .Q(w5102) );
	vdp_xor g5119 (.Z(w5055), .B(w5102), .A(VRAMA[14]) );
	vdp_xor g5120 (.Z(w5054), .B(w5058), .A(VRAMA[11]) );
	vdp_slatch g5121 (.D(S[5]), .nC(w4864), .C(w4865), .Q(w5073) );
	vdp_slatch g5122 (.D(S[5]), .nC(w4862), .C(w4861), .Q(w5053) );
	vdp_slatch g5123 (.D(S[6]), .nC(w4864), .C(w4865), .Q(w5074) );
	vdp_slatch g5124 (.D(S[6]), .nC(w4862), .C(w4861), .Q(w5072) );
	vdp_slatch g5125 (.D(S[7]), .nC(w4864), .C(w4865), .Q(w5107) );
	vdp_slatch g5126 (.D(S[7]), .nC(w4862), .C(w4861), .Q(w5039) );
	vdp_slatch g5127 (.D(REG_BUS[2]), .nC(w5077), .C(w5078), .Q(w5075) );
	vdp_slatch g5128 (.D(REG_BUS[5]), .nC(w5077), .C(w5078), .Q(w5071) );
	vdp_bufif0 g5129 (.A(w5058), .Z(VRAMA[9]), .nE(w5012) );
	vdp_bufif0 g5130 (.A(w5008), .Z(VRAMA[10]), .nE(w5041) );
	vdp_bufif0 g5131 (.A(w5096), .Z(VRAMA[10]), .nE(w5012) );
	vdp_bufif0 g5132 (.A(w5059), .Z(VRAMA[13]), .nE(w5012) );
	vdp_bufif0 g5133 (.A(w5102), .Z(VRAMA[14]), .nE(w5041) );
	vdp_bufif0 g5134 (.A(w5058), .Z(VRAMA[11]), .nE(w5041) );
	vdp_bufif0 g5135 (.A(w5095), .Z(VRAMA[13]), .nE(w5041) );
	vdp_bufif0 g5136 (.A(w5096), .Z(VRAMA[12]), .nE(w5041) );
	vdp_bufif0 g5137 (.A(w5095), .Z(VRAMA[11]), .nE(w5012) );
	vdp_bufif0 g5138 (.A(w5102), .Z(VRAMA[12]), .nE(w5012) );
	vdp_bufif0 g5139 (.A(w5059), .Z(VRAMA[15]), .nE(w5041) );
	vdp_slatch g5140 (.D(REG_BUS[3]), .nC(w5111), .C(w5110), .Q(w5096) );
	vdp_slatch g5141 (.D(REG_BUS[4]), .nC(w5111), .C(w5110), .Q(w5095) );
	vdp_xor g5142 (.Z(w5057), .B(w5095), .A(VRAMA[13]) );
	vdp_xor g5143 (.Z(w5056), .B(w5096), .A(VRAMA[12]) );
	vdp_dlatch_inv g5144 (.nQ(w5094), .D(w5099), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5145 (.nQ(w5093), .D(w5100), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5146 (.nQ(w5092), .D(w6422), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5147 (.nQ(w5091), .D(w6424), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5148 (.nQ(w5090), .D(w5101), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5149 (.nQ(w5089), .D(w5098), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5150 (.nQ(w5088), .D(w6423), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5151 (.nQ(w6160), .D(w5097), .nC(nDCLK1), .C(DCLK1) );
	vdp_comp_we g5152 (.nZ(w5112), .A(w5007), .Z(w5113) );
	vdp_comp_we g5153 (.nZ(w4951), .A(w5007), .Z(w6552) );
	vdp_comp_we g5154 (.nZ(w6554), .A(w5007), .Z(w6553) );
	vdp_comp_we g5155 (.nZ(w6555), .A(w5007), .Z(w6556) );
	vdp_comp_we g5156 (.nZ(w6557), .A(w5007), .Z(w6558) );
	vdp_comp_we g5157 (.nZ(w6559), .A(w5007), .Z(w6560) );
	vdp_comp_we g5158 (.nZ(w6561), .A(w5007), .Z(w6562) );
	vdp_comp_we g5159 (.nZ(w6563), .A(w5007), .Z(w6564) );
	vdp_comp_we g5160 (.nZ(w6565), .A(w5007), .Z(w6566) );
	vdp_comp_we g5161 (.nZ(w6567), .A(w5007), .Z(w6568) );
	vdp_comp_we g5162 (.nZ(w5108), .A(w110), .Z(w5109) );
	vdp_notif0 g5163 (.A(w5048), .nZ(VRAMA[10]), .nE(w4974) );
	vdp_notif0 g5164 (.A(w5076), .nZ(VRAMA[13]), .nE(w4974) );
	vdp_notif0 g5165 (.A(w5106), .nZ(VRAMA[11]), .nE(w4974) );
	vdp_notif0 g5166 (.A(w5105), .nZ(VRAMA[12]), .nE(w4974) );
	vdp_not g5167 (.nZ(w5050), .A(VRAMA[2]) );
	vdp_not g5168 (.nZ(w5076), .A(w5075) );
	vdp_not g5169 (.nZ(w5104), .A(w106) );
	vdp_aoi22 g5170 (.Z(w4817), .B2(w5039), .B1(w5049), .A1(w4916), .A2(w5060) );
	vdp_aoi22 g5171 (.Z(w5048), .B2(w5039), .B1(w5073), .A1(w4916), .A2(w5053) );
	vdp_aoi22 g5172 (.Z(w4810), .B2(w5039), .B1(w5061), .A1(w4916), .A2(w6316) );
	vdp_aoi22 g5173 (.Z(w5106), .B2(w5039), .B1(w5074), .A1(w4916), .A2(w5072) );
	vdp_aoi22 g5174 (.Z(w5105), .B2(w5039), .B1(w5107), .A1(w4916), .A2(w5039) );
	vdp_and g5175 (.Z(w5103), .B(w5104), .A(w4410) );
	vdp_nor8 g5176 (.Z(w5047), .B(w5056), .A(w5057), .C(w5055), .D(w5054), .F(w5044), .E(w5040), .G(w5042), .H(w5043) );
	vdp_not g5177 (.nZ(w5114), .A(w109) );
	vdp_comp_str g5178 (.nZ(w5111), .A(w159), .Z(w5110) );
	vdp_comp_str g5179 (.nZ(w5078), .A(w160), .Z(w5077) );
	vdp_or3 g5180 (.Z(w5007), .B(w110), .A(w109), .C(w5103) );
	vdp_not g5181 (.nZ(S[7]), .A(w5094) );
	vdp_not g5182 (.nZ(S[6]), .A(w5093) );
	vdp_not g5183 (.nZ(S[5]), .A(w5092) );
	vdp_not g5184 (.nZ(S[4]), .A(w5091) );
	vdp_not g5185 (.nZ(S[3]), .A(w5090) );
	vdp_not g5186 (.nZ(S[2]), .A(w5089) );
	vdp_not g5187 (.nZ(S[1]), .A(w5088) );
	vdp_not g5188 (.nZ(S[0]), .A(w6160) );
	vdp_aon21_sr g5189 (.Q(w5182), .A1(w5181), .A2(w6230), .B(w6231), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5190 (.Q(w6231), .A1(w5176), .A2(w6230), .B(w6569), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5191 (.Q(w6569), .A1(w5177), .A2(w6230), .B(w6570), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5192 (.Q(w6570), .A1(w5126), .A2(w6230), .B(w6571), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5193 (.Q(w6571), .A1(w5175), .A2(w6230), .B(w6572), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5194 (.Q(w6572), .A1(w5174), .A2(w6230), .B(w6573), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5195 (.Q(w6573), .A1(w5173), .A2(w6230), .B(w6574), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5196 (.Q(w6574), .A1(w5172), .A2(w6230), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5197 (.Q(w6575), .A1(w5162), .A2(w6232), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5198 (.Q(w6576), .A1(w5156), .A2(w6232), .B(w6575), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5199 (.Q(w6577), .A1(w5158), .A2(w6232), .B(w6576), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5200 (.Q(w6578), .A1(w5155), .A2(w6232), .B(w6577), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5201 (.Q(w6579), .A1(w5125), .A2(w6232), .B(w6578), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5202 (.Q(w6580), .A1(w5153), .A2(w6232), .B(w6579), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5203 (.Q(w6581), .A1(w5154), .A2(w6232), .B(w6580), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5204 (.Q(w5146), .A1(w5152), .A2(w6232), .B(w6581), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5205 (.Q(w5288), .A1(w5143), .A2(w6229), .B(w6582), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5206 (.Q(w6582), .A1(w5141), .A2(w6229), .B(w6583), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5207 (.Q(w6583), .A1(w5144), .A2(w6229), .B(w6584), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5208 (.Q(w6584), .A1(w5139), .A2(w6229), .B(w6585), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5209 (.Q(w6585), .A1(w5117), .A2(w6229), .B(w6586), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5210 (.Q(w6586), .A1(w5138), .A2(w6229), .B(w6587), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5211 (.Q(w6587), .A1(w5140), .A2(w6229), .B(w6588), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5212 (.Q(w6588), .A1(w5135), .A2(w6229), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5213 (.Q(w6590), .A1(w5187), .A2(w6228), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5214 (.Q(w6591), .A1(w5186), .A2(w6228), .B(w6590), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5215 (.Q(w6592), .A1(w5511), .A2(w6228), .B(w6591), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5216 (.Q(w6593), .A1(w5194), .A2(w6228), .B(w6592), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5217 (.Q(w6594), .A1(w5192), .A2(w6228), .B(w6593), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5218 (.Q(w6595), .A1(w5198), .A2(w6228), .B(w6594), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5219 (.Q(w6596), .A1(w5191), .A2(w6228), .B(w6595), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5220 (.Q(w5115), .A1(w5124), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .A2(w6228), .B(w6596) );
	vdp_not g5221 (.nZ(w6229), .A(w5167) );
	vdp_not g5222 (.nZ(w6228), .A(w5167) );
	vdp_not g5223 (.nZ(w6232), .A(w5167) );
	vdp_not g5224 (.nZ(w6230), .A(w5167) );
	vdp_or4 g5225 (.Z(w5180), .B(w5169), .A(w6161), .D(w5170), .C(w5168) );
	vdp_or4 g5226 (.Z(w5150), .B(w5166), .A(w5159), .D(w5164), .C(w5165) );
	vdp_or4 g5227 (.Z(w5183), .B(w5123), .A(w5124), .D(w5507), .C(w5122) );
	vdp_or4 g5228 (.Z(w5149), .B(w5121), .A(w5504), .D(w5191), .C(w5120) );
	vdp_or4 g5229 (.Z(w5145), .B(w5119), .A(w5503), .D(w5198), .C(w5118) );
	vdp_or4 g5230 (.Z(w5188), .B(w5128), .A(w5129), .D(w6162), .C(w5127) );
	vdp_or4 g5231 (.Z(w5134), .B(w5132), .A(w5133), .D(w5116), .C(w5131) );
	vdp_slatch g5232 (.Q(w5170), .D(w5235), .nC(w5160), .C(w5161) );
	vdp_comp_str g5233 (.nZ(w5160), .A(w5207), .Z(w5161) );
	vdp_slatch g5234 (.Q(w5168), .D(w5233), .nC(w5160), .C(w5161) );
	vdp_slatch g5235 (.Q(w5169), .D(w5232), .nC(w5160), .C(w5161) );
	vdp_slatch g5236 (.Q(w6161), .D(w5231), .nC(w5160), .C(w5161) );
	vdp_slatch g5237 (.Q(w5164), .D(w5230), .nC(w5160), .C(w5161) );
	vdp_slatch g5238 (.Q(w5165), .D(w5229), .nC(w5160), .C(w5161) );
	vdp_slatch g5239 (.Q(w5166), .D(w5227), .nC(w5160), .C(w5161) );
	vdp_slatch g5240 (.Q(w5159), .D(w5223), .nC(w5160), .C(w5161) );
	vdp_slatch g5241 (.Q(w5116), .D(w6225), .nC(w5130), .C(w5190) );
	vdp_slatch g5242 (.Q(w5131), .D(w6226), .nC(w5130), .C(w5190) );
	vdp_slatch g5243 (.Q(w5132), .D(w6227), .nC(w5130), .C(w5190) );
	vdp_slatch g5244 (.Q(w5133), .D(w5213), .nC(w5130), .C(w5190) );
	vdp_slatch g5245 (.Q(w6162), .D(w5211), .nC(w5130), .C(w5190) );
	vdp_slatch g5246 (.Q(w5127), .D(w5210), .nC(w5130), .C(w5190) );
	vdp_slatch g5247 (.Q(w5128), .D(w5209), .nC(w5130), .C(w5190) );
	vdp_slatch g5248 (.Q(w5129), .D(w5206), .nC(w5130), .C(w5190) );
	vdp_aon22 g5249 (.Z(w5243), .B2(w5136), .B1(w5196), .A1(w5188), .A2(w5148) );
	vdp_comp_we g5250 (.nZ(w5136), .A(w5195), .Z(w5148) );
	vdp_notif0 g5251 (.A(w5189), .nZ(DB[11]), .nE(w5205) );
	vdp_notif0 g5252 (.A(w5193), .nZ(DB[3]), .nE(w5205) );
	vdp_notif0 g5253 (.A(w5137), .nZ(DB[10]), .nE(w5205) );
	vdp_notif0 g5254 (.A(w5142), .nZ(DB[2]), .nE(w5205) );
	vdp_notif0 g5255 (.A(w5157), .nZ(DB[1]), .nE(w5205) );
	vdp_notif0 g5256 (.A(w5199), .nZ(DB[9]), .nE(w5205) );
	vdp_notif0 g5257 (.A(w5178), .nZ(DB[8]), .nE(w5205) );
	vdp_notif0 g5258 (.A(w5179), .nZ(DB[0]), .nE(w5205) );
	vdp_not g5259 (.nZ(w5184), .A(w5183) );
	vdp_aon22 g5260 (.Z(w5216), .B2(w5136), .B1(w5147), .A1(w5134), .A2(w5148) );
	vdp_aon22 g5261 (.Z(w5221), .B2(w5136), .B1(w5151), .A1(w5150), .A2(w5148) );
	vdp_aon22 g5262 (.Z(w5238), .B2(w5136), .B1(w5184), .A1(w5180), .A2(w5148) );
	vdp_comp_str g5263 (.nZ(w5130), .A(w5207), .Z(w5190) );
	vdp_not g5264 (.nZ(w5196), .A(w5197) );
	vdp_not g5265 (.nZ(w5147), .A(w5145) );
	vdp_not g5266 (.nZ(w5151), .A(w5149) );
	vdp_and3 g5267 (.Z(w6210), .B(w5219), .A(w5150), .C(w5149) );
	vdp_and3 g5268 (.Z(w5225), .B(w5239), .A(w5180), .C(w5183) );
	vdp_and3 g5269 (.Z(w5241), .B(w5217), .A(w5134), .C(w5145) );
	vdp_and3 g5270 (.Z(w5570), .B(w5188), .A(w5200), .C(w5197) );
	vdp_aon2222 g5271 (.Z(w5193), .B2(w5194), .B1(w5203), .A1(w5204), .A2(w5186), .D2(w5124), .D1(w5201), .C1(w5202), .C2(w5198) );
	vdp_aon2222 g5272 (.Z(w5189), .B2(w5511), .B1(w5203), .A1(w5204), .A2(w5187), .D2(w5191), .D1(w5201), .C1(w5202), .C2(w5192) );
	vdp_aon2222 g5273 (.Z(w5137), .B2(w5138), .B1(w5203), .A1(w5204), .A2(w5135), .D2(w5141), .D1(w5201), .C1(w5202), .C2(w5139) );
	vdp_aon2222 g5274 (.Z(w5142), .B2(w5117), .B1(w5203), .A1(w5204), .A2(w5140), .D2(w5143), .D1(w5201), .C1(w5202), .C2(w5144) );
	vdp_aon2222 g5275 (.Z(w5157), .B2(w5155), .B1(w5203), .A1(w5204), .A2(w5156), .D2(w5152), .D1(w5201), .C1(w5202), .C2(w5153) );
	vdp_aon2222 g5276 (.Z(w5199), .B2(w5158), .B1(w5203), .A1(w5204), .A2(w5162), .D2(w5154), .D1(w5201), .C1(w5202), .C2(w5125) );
	vdp_aon2222 g5277 (.Z(w5178), .B2(w5174), .B1(w5203), .A1(w5204), .A2(w5172), .D2(w5176), .D1(w5201), .C1(w5202), .C2(w5126) );
	vdp_aon2222 g5278 (.Z(w5179), .B2(w5175), .B1(w5203), .A1(w5204), .A2(w5173), .D2(w5181), .D1(w5201), .C1(w5202), .C2(w5177) );
	vdp_slatch g5279 (.Q(w5235), .D(w5255), .nC(w5254), .C(w5234) );
	vdp_comp_str g5280 (.nZ(w5254), .A(w5253), .Z(w5234) );
	vdp_slatch g5281 (.Q(w5233), .D(w5259), .nC(w5254), .C(w5234) );
	vdp_slatch g5282 (.Q(w5232), .D(w5260), .nC(w5254), .C(w5234) );
	vdp_slatch g5283 (.Q(w5231), .D(w5263), .nC(w5254), .C(w5234) );
	vdp_slatch g5284 (.Q(w5230), .D(w5268), .nC(w5269), .C(w5228) );
	vdp_comp_str g5285 (.nZ(w5269), .A(w5264), .Z(w5228) );
	vdp_slatch g5286 (.Q(w5229), .D(w5271), .nC(w5269), .C(w5228) );
	vdp_slatch g5287 (.Q(w5227), .D(w5272), .nC(w5269), .C(w5228) );
	vdp_slatch g5288 (.Q(w5223), .D(w5274), .nC(w5269), .C(w5228) );
	vdp_sr_bit g5289 (.Q(w5276), .D(w5146), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5290 (.nQ(w5222), .D(w5278), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5291 (.nQ(w5280), .D(w5220), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5292 (.nQ(w5218), .D(w5287), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5293 (.nQ(w5293), .D(w6203), .nC(nDCLK2), .C(DCLK2) );
	vdp_slatch g5294 (.Q(w5213), .D(w5255), .nC(w5295), .C(w5215) );
	vdp_slatch g5295 (.Q(w6225), .D(w5259), .nC(w5295), .C(w5215) );
	vdp_slatch g5296 (.Q(w6226), .D(w5260), .nC(w5295), .C(w5215) );
	vdp_slatch g5297 (.Q(w6227), .D(w5263), .nC(w5295), .C(w5215) );
	vdp_comp_str g5298 (.nZ(w5295), .A(w5294), .Z(w5215) );
	vdp_slatch g5299 (.Q(w5211), .D(w5268), .nC(w5306), .C(w5208) );
	vdp_slatch g5300 (.Q(w5210), .D(w5271), .nC(w5306), .C(w5208) );
	vdp_slatch g5301 (.Q(w5209), .D(w5272), .nC(w5306), .C(w5208) );
	vdp_slatch g5302 (.Q(w5206), .D(w5274), .nC(w5306), .C(w5208) );
	vdp_comp_str g5303 (.nZ(w5306), .A(w5311), .Z(w5208) );
	vdp_dlatch_inv g5304 (.nQ(w5304), .D(w5303), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5305 (.nQ(w5307), .D(w6202), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5306 (.nQ(w5242), .D(w5310), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5307 (.Z(w5309), .B(w5242), .A(w5246) );
	vdp_xor g5308 (.Z(w6221), .B(w5218), .A(w5246) );
	vdp_xor g5309 (.Z(w5277), .B(w5222), .A(w5246) );
	vdp_xor g5310 (.Z(w6170), .B(w6169), .A(w5246) );
	vdp_sr_bit g5311 (.Q(w6224), .D(w5182), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5312 (.nQ(w6169), .D(w5244), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5313 (.nQ(w6171), .D(w5237), .nC(nDCLK2), .C(DCLK2) );
	vdp_and g5314 (.Z(w5239), .B(w6170), .A(w5247) );
	vdp_and g5315 (.Z(w5240), .B(w6171), .A(DCLK1) );
	vdp_and g5316 (.Z(w5224), .B(w5280), .A(DCLK1) );
	vdp_and g5317 (.Z(w5219), .B(w5277), .A(w5247) );
	vdp_and g5318 (.Z(w5201), .B(w5282), .A(w5281) );
	vdp_and g5319 (.Z(w5202), .B(w74), .A(w5282) );
	vdp_and g5320 (.Z(w5203), .B(w75), .A(w5281) );
	vdp_and g5321 (.Z(w5204), .B(w74), .A(w75) );
	vdp_and g5322 (.Z(w5217), .B(w6221), .A(w5247) );
	vdp_and g5323 (.Z(w5236), .B(w5293), .A(DCLK1) );
	vdp_and g5324 (.Z(w5226), .B(w5307), .A(DCLK1) );
	vdp_and g5325 (.Z(w5200), .B(w5309), .A(w5247) );
	vdp_sr_bit g5326 (.Q(w5285), .D(w5288), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5327 (.Q(w5296), .D(w5266), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_not g5328 (.nZ(w5207), .A(w5214) );
	vdp_not g5329 (.nZ(w5212), .A(w114) );
	vdp_not g5330 (.nZ(w5281), .A(w74) );
	vdp_not g5331 (.nZ(w5282), .A(w75) );
	vdp_aoi21 g5332 (.Z(w5237), .B(w5250), .A1(w5238), .A2(w5239) );
	vdp_aoi21 g5333 (.Z(w5220), .B(w5250), .A1(w5221), .A2(w5219) );
	vdp_aoi21 g5334 (.Z(w6203), .B(w5292), .A1(w5216), .A2(w5217) );
	vdp_oai21 g5335 (.Z(w5214), .B(DCLK2), .A1(w5297), .A2(w5296) );
	vdp_aoi21 g5336 (.Z(w6202), .B(w5292), .A1(w5200), .A2(w5243) );
	vdp_not g5337 (.nZ(w5205), .A(w115) );
	vdp_nand g5338 (.Z(w5266), .B(w5304), .A(w5212) );
	vdp_sr_bit g5339 (.Q(w5257), .D(w5313), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5340 (.Q(w5262), .D(w6172), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5341 (.Q(w5273), .D(w6223), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5342 (.Q(w5258), .D(w5275), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5343 (.Q(w5279), .D(w2612), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5344 (.Q(w5283), .D(w5284), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5345 (.Q(w6214), .D(w5300), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5346 (.Q(w5300), .D(w5312), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5347 (.Q(w5314), .D(w5115), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g5348 (.Z(w5312), .B2(w5115), .B1(w5318), .A1(w5317), .A2(w5314) );
	vdp_aon22 g5349 (.Z(w5284), .B2(w5288), .B1(w5318), .A1(w5317), .A2(w5285) );
	vdp_aon22 g5350 (.Z(w5275), .B2(w5146), .B1(w5318), .A1(w5317), .A2(w5276) );
	vdp_aon22 g5351 (.Z(w5313), .B2(w5182), .B1(w5318), .A1(w5317), .A2(w6224) );
	vdp_not g5352 (.nZ(w5256), .A(w5310) );
	vdp_not g5353 (.nZ(w5248), .A(w75) );
	vdp_not g5354 (.nZ(w5253), .A(w5330) );
	vdp_not g5355 (.nZ(w5261), .A(M5) );
	vdp_not g5356 (.nZ(w5264), .A(w5265) );
	vdp_not g5357 (.nZ(w5251), .A(w5323) );
	vdp_not g5358 (.nZ(w5245), .A(w5321) );
	vdp_not g5359 (.nZ(w5294), .A(w5291) );
	vdp_not g5360 (.nZ(w5311), .A(w5299) );
	vdp_not g5361 (.nZ(w5305), .A(w5300) );
	vdp_comp_we g5362 (.nZ(w5318), .A(M5), .Z(w5317) );
	vdp_and g5363 (.Z(w2729), .B(w5258), .A(w5257) );
	vdp_or g5364 (.Z(w6172), .B(w5257), .A(w5261) );
	vdp_or g5365 (.Z(w5267), .B(w5270), .A(w5266) );
	vdp_and g5366 (.Z(w6223), .B(w5258), .A(M5) );
	vdp_and g5367 (.Z(w2612), .B(w5283), .A(M5) );
	vdp_or g5368 (.Z(w5308), .B(w5266), .A(w5298) );
	vdp_not g5369 (.nZ(w5329), .A(SPR_PRIO) );
	vdp_bufif0 g5370 (.A(w6214), .Z(COL[0]), .nE(w5329) );
	vdp_oai21 g5371 (.Z(w5291), .B(DCLK2), .A1(w5267), .A2(w5290) );
	vdp_bufif0 g5372 (.A(w5279), .Z(COL[6]), .nE(w5329) );
	vdp_bufif0 g5373 (.A(w5273), .Z(COL[5]), .nE(w5329) );
	vdp_bufif0 g5374 (.A(w5262), .Z(COL[4]), .nE(w5329) );
	vdp_oai21 g5375 (.Z(w5265), .B(DCLK2), .A1(w5267), .A2(w5252) );
	vdp_oai21 g5376 (.Z(w5330), .B(DCLK2), .A1(w5324), .A2(w5252) );
	vdp_and3 g5377 (.Z(w5252), .B(w5328), .A(w5251), .C(w5327) );
	vdp_and3 g5378 (.Z(w5270), .B(w5328), .A(w5251), .C(w5315) );
	vdp_and3 g5379 (.Z(w5290), .B(w5327), .A(w5316), .C(w5251) );
	vdp_and3 g5380 (.Z(w5298), .B(w5315), .A(w5316), .C(w5251) );
	vdp_or4 g5381 (.Z(w2611), .B(w5320), .A(w5302), .D(w5300), .C(w5301) );
	vdp_and4 g5382 (.Z(w2669), .B(w5301), .A(w5320), .D(w5305), .C(w5302) );
	vdp_and4 g5383 (.Z(w2668), .B(w5301), .A(w5320), .D(w5300), .C(w5302) );
	vdp_oai21 g5384 (.Z(w5299), .B(DCLK2), .A1(w5290), .A2(w5308) );
	vdp_nand3 g5385 (.Z(w5244), .B(w5245), .A(w5256), .C(w5326) );
	vdp_nand3 g5386 (.Z(w5249), .B(w5325), .A(w105), .C(w5248) );
	vdp_nand3 g5387 (.Z(w5289), .B(w74), .A(w105), .C(w5248) );
	vdp_nand g5388 (.Z(w5292), .B(w5289), .A(w5319) );
	vdp_nand g5389 (.Z(w5286), .B(w5322), .A(w5321) );
	vdp_nand g5390 (.Z(w5287), .B(w5256), .A(w5286) );
	vdp_nand g5391 (.Z(w5278), .B(w5245), .A(w5256) );
	vdp_nand g5392 (.Z(w5250), .B(w5249), .A(w5319) );
	vdp_sr_bit g5393 (.Q(w6175), .D(w6174), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5394 (.Q(w6176), .D(w6175), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5395 (.Q(w5394), .D(w6176), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5396 (.Q(w5401), .D(w5394), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5397 (.Q(w5303), .D(w6177), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5398 (.Q(w6222), .D(w5402), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5399 (.Q(w5404), .D(w6233), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5400 (.Q(w5385), .D(w6173), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_dlatch_inv g5401 (.nQ(w5352), .D(w5344), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5402 (.nQ(w5357), .D(w5343), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5403 (.nQ(w5363), .D(w5342), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5404 (.nQ(w5368), .D(w5341), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5405 (.nQ(w5369), .D(w5340), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5406 (.nQ(w5372), .D(w5339), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5407 (.nQ(w5373), .D(w5338), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5408 (.nQ(w5376), .D(w5336), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5409 (.nQ(w5398), .D(w5399), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5410 (.nQ(w5396), .D(w5381), .nC(nDCLK1), .C(DCLK1) );
	vdp_cnt_bit_load g5411 (.Q(w5399), .D(w5400), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1), .R(1'b0), .CI(w6235), .L(w5333), .nL(w5378) );
	vdp_cnt_bit_load g5412 (.Q(w5381), .D(w5380), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1), .R(1'b0), .CI(w5334), .L(w5333), .nL(w5378), .CO(w6235) );
	vdp_aon22 g5413 (.Z(w5268), .B2(w5335), .B1(DB[11]), .A1(w5376), .A2(w5353) );
	vdp_aon22 g5414 (.Z(w5336), .B2(w5337), .B1(w5365), .A1(w5364), .A2(w5356) );
	vdp_aon22 g5415 (.Z(w5271), .B2(w5335), .B1(DB[12]), .A1(w5373), .A2(w5353) );
	vdp_aon22 g5416 (.Z(w5338), .B2(w5337), .B1(w5361), .A1(w5362), .A2(w5356) );
	vdp_aon22 g5417 (.Z(w5272), .B2(w5335), .B1(DB[13]), .A1(w5372), .A2(w5353) );
	vdp_aon22 g5418 (.Z(w5339), .B2(w5337), .B1(w5354), .A1(w5355), .A2(w5356) );
	vdp_aon22 g5419 (.Z(w5274), .B2(w5335), .B1(DB[14]), .A1(w5369), .A2(w5353) );
	vdp_aon22 g5420 (.Z(w5340), .B2(w5337), .B1(w5345), .A1(w5346), .A2(w5356) );
	vdp_aon22 g5421 (.Z(w5255), .B2(w5335), .B1(DB[3]), .A1(w5368), .A2(w5353) );
	vdp_aon22 g5422 (.Z(w5341), .B2(w5337), .B1(w5364), .A1(w5365), .A2(w5356) );
	vdp_aon22 g5423 (.Z(w5259), .B2(w5335), .B1(DB[4]), .A1(w5363), .A2(w5353) );
	vdp_aon22 g5424 (.Z(w5342), .B2(w5337), .B1(w5362), .A1(w5361), .A2(w5356) );
	vdp_aon22 g5425 (.Z(w5260), .B2(w5335), .B1(DB[5]), .A1(w5357), .A2(w5353) );
	vdp_aon22 g5426 (.Z(w5343), .B2(w5337), .B1(w5355), .A1(w5354), .A2(w5356) );
	vdp_aon22 g5427 (.Z(w5263), .B2(w5335), .B1(DB[6]), .A1(w5352), .A2(w5353) );
	vdp_aon22 g5428 (.Z(w5344), .B2(w5337), .B1(w5346), .A1(w5345), .A2(w5356) );
	vdp_slatch g5429 (.Q(w6173), .D(w5388), .nC(w5332), .C(w5389) );
	vdp_dlatch_inv g5430 (.nQ(w5386), .D(w5385), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5431 (.nQ(w5402), .D(w25), .nC(nHCLK1), .C(HCLK1) );
	vdp_xnor g5432 (.Z(w5316), .B(1'b0), .A(w5396) );
	vdp_xor g5433 (.Z(w5377), .B(w5385), .A(w5387) );
	vdp_aon22 g5434 (.Z(w6233), .B2(w5394), .B1(M5), .A1(w5401), .A2(w6234) );
	vdp_not g5435 (.nZ(w5403), .A(w5402) );
	vdp_not g5436 (.nZ(w6234), .A(M5) );
	vdp_not g5437 (.nZ(w5332), .A(w5389) );
	vdp_not g5438 (.nZ(w6174), .A(w5392) );
	vdp_not g5439 (.nZ(w5315), .A(w5386) );
	vdp_not g5440 (.nZ(w5323), .A(w5398) );
	vdp_not g5441 (.nZ(w5334), .A(w5389) );
	vdp_comp_we g5442 (.nZ(w5353), .A(w114), .Z(w5335) );
	vdp_comp_we g5443 (.nZ(w5356), .A(w5377), .Z(w5337) );
	vdp_comp_we g5444 (.nZ(w5378), .A(w5389), .Z(w5333) );
	vdp_and g5445 (.Z(w6177), .B(w6222), .A(w5403) );
	vdp_aoi21 g5446 (.Z(w5392), .B(w24), .A1(M5), .A2(w21) );
	vdp_sr_bit g5447 (.Q(w5387), .D(w5448), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_aon22 g5448 (.Z(w5456), .B2(w5450), .B1(w5449), .A1(w5446), .A2(w5395) );
	vdp_aon22 g5449 (.Z(w5455), .B2(w5450), .B1(w5453), .A1(w5451), .A2(w5395) );
	vdp_aon22 g5450 (.Z(w5452), .B2(w5450), .B1(w5451), .A1(w5453), .A2(w5395) );
	vdp_aon22 g5451 (.Z(w5457), .B2(w5450), .B1(w5446), .A1(w5449), .A2(w5395) );
	vdp_not g5452 (.nZ(w5413), .A(w5449) );
	vdp_not g5453 (.nZ(w5414), .A(w5453) );
	vdp_not g5454 (.nZ(w5419), .A(w5451) );
	vdp_not g5455 (.nZ(w5418), .A(w5446) );
	vdp_not g5456 (.nZ(w5348), .A(w5455) );
	vdp_not g5457 (.nZ(w5349), .A(w5456) );
	vdp_not g5458 (.nZ(w5350), .A(w5457) );
	vdp_not g5459 (.nZ(w5351), .A(w5452) );
	vdp_not g5460 (.nZ(w5393), .A(M5) );
	vdp_comp_we g5461 (.nZ(w5450), .A(w5387), .Z(w5395) );
	vdp_not g5462 (.nZ(w5389), .A(w5447) );
	vdp_not g5463 (.nZ(w5445), .A(w5444) );
	vdp_dlatch_inv g5464 (.nQ(w5444), .D(w5443), .nC(nHCLK1), .C(HCLK1) );
	vdp_aon2222 g5465 (.Z(w5347), .B2(w5349), .B1(w5407), .A1(w5406), .A2(w5348), .D2(w5351), .D1(w5424), .C1(w5423), .C2(w5350) );
	vdp_aon2222 g5466 (.Z(w5397), .B2(w5419), .B1(w5411), .A1(w5418), .A2(w5406), .D2(w5413), .D1(w5415), .C1(w5414), .C2(w5458) );
	vdp_aon2222 g5467 (.Z(w5367), .B2(w5349), .B1(w5412), .A1(w5411), .A2(w5348), .D2(w5351), .D1(w5416), .C1(w5459), .C2(w5350) );
	vdp_aon2222 g5468 (.Z(w5358), .B2(w5419), .B1(w5412), .A1(w5418), .A2(w5407), .D2(w5413), .D1(w5426), .C1(w5414), .C2(w5420) );
	vdp_aon2222 g5469 (.Z(w5375), .B2(w5349), .B1(w5420), .A1(w5458), .A2(w5348), .D2(w5351), .D1(w5422), .C1(w5421), .C2(w5350) );
	vdp_aon2222 g5470 (.Z(w5366), .B2(w5419), .B1(w5459), .A1(w5418), .A2(w5423), .D2(w5413), .D1(w5425), .C1(w5414), .C2(w5421) );
	vdp_aon2222 g5471 (.Z(w6201), .B2(w5349), .B1(w5426), .A1(w5415), .A2(w5348), .D2(w5351), .D1(w5427), .C1(w5425), .C2(w5350) );
	vdp_aon2222 g5472 (.Z(w5370), .B2(w5419), .B1(w5416), .A1(w5418), .A2(w5424), .D2(w5413), .D1(w5427), .C1(w5414), .C2(w5422) );
	vdp_aon2222 g5473 (.Z(w5359), .B2(w5349), .B1(w5429), .A1(w5428), .A2(w5348), .D2(w5351), .D1(w5441), .C1(w5430), .C2(w5350) );
	vdp_aon2222 g5474 (.Z(w5374), .B2(w5419), .B1(w5431), .A1(w5418), .A2(w5428), .D2(w5413), .D1(w5432), .C1(w5414), .C2(w5433) );
	vdp_aon2222 g5475 (.Z(w5371), .B2(w5349), .B1(w5435), .A1(w5431), .A2(w5348), .D2(w5351), .D1(w5434), .C1(w5436), .C2(w5350) );
	vdp_aon2222 g5476 (.Z(w5383), .B2(w5419), .B1(w5435), .A1(w5418), .A2(w5429), .D2(w5413), .D1(w5437), .C1(w5414), .C2(w5438) );
	vdp_aon2222 g5477 (.Z(w5382), .B2(w5349), .B1(w5438), .A1(w5433), .A2(w5348), .D2(w5351), .D1(w5439), .C1(w5440), .C2(w5350) );
	vdp_aon2222 g5478 (.Z(w5384), .B2(w5419), .B1(w5436), .A1(w5418), .A2(w5430), .D2(w5413), .D1(w5442), .C1(w5414), .C2(w5440) );
	vdp_aon2222 g5479 (.Z(w5391), .B2(w5349), .B1(w5437), .A1(w5432), .A2(w5348), .D2(w5351), .D1(w5454), .C1(w5442), .C2(w5350) );
	vdp_aon2222 g5480 (.Z(w5390), .B2(w5419), .B1(w5434), .A1(w5418), .A2(w5441), .D2(w5413), .D1(w5454), .C1(w5414), .C2(w5439) );
	vdp_aoi22 g5481 (.Z(w5345), .B2(w5405), .B1(w5347), .A1(w5360), .A2(w5397) );
	vdp_aoi22 g5482 (.Z(w5354), .B2(w5405), .B1(w5359), .A1(w5360), .A2(w5358) );
	vdp_aoi22 g5483 (.Z(w5361), .B2(w5405), .B1(w5367), .A1(w5360), .A2(w5366) );
	vdp_aoi22 g5484 (.Z(w5365), .B2(w5405), .B1(w5371), .A1(w5360), .A2(w5370) );
	vdp_aoi22 g5485 (.Z(w5346), .B2(w5405), .B1(w5375), .A1(w5360), .A2(w5374) );
	vdp_aoi22 g5486 (.Z(w5355), .B2(w5405), .B1(w5382), .A1(w5360), .A2(w5383) );
	vdp_aoi22 g5487 (.Z(w5362), .B2(w5405), .B1(w6201), .A1(w5360), .A2(w5384) );
	vdp_aoi22 g5488 (.Z(w5364), .B2(w5405), .B1(w5391), .A1(w5360), .A2(w5390) );
	vdp_nand g5489 (.Z(w5447), .B(w5445), .A(HCLK2) );
	vdp_nor g5490 (.Z(w5405), .B(w5393), .A(w5303) );
	vdp_nor g5491 (.Z(w5360), .B(M5), .A(w5303) );
	vdp_sr_bit g5492 (.Q(w5449), .D(w5453), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5493 (.Q(w5453), .D(w5451), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5494 (.Q(w5451), .D(w5446), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5495 (.Q(w5446), .D(w5447), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_dlatch_inv g5496 (.nQ(w5297), .D(w5449), .nC(nDCLK1), .C(DCLK1) );
	vdp_comp_str g5497 (.nZ(w5410), .A(w5460), .Z(w5462) );
	vdp_comp_str g5498 (.nZ(w5409), .A(w5460), .Z(w5465) );
	vdp_comp_str g5499 (.nZ(w5417), .A(w5460), .Z(w5466) );
	vdp_comp_str g5500 (.nZ(w5408), .A(w5460), .Z(w5461) );
	vdp_slatch g5501 (.D(w5475), .Q(w5406), .nC(w5408), .C(w5461) );
	vdp_slatch g5502 (.D(w6259), .Q(w5407), .nC(w5417), .C(w5466) );
	vdp_slatch g5503 (.D(w6258), .Q(w5423), .nC(w5409), .C(w5465) );
	vdp_slatch g5504 (.D(w6257), .Q(w5424), .nC(w5410), .C(w5462) );
	vdp_slatch g5505 (.D(w5474), .Q(w5411), .nC(w5408), .C(w5461) );
	vdp_slatch g5506 (.D(w6256), .Q(w5412), .nC(w5417), .C(w5466) );
	vdp_slatch g5507 (.D(w6255), .Q(w5459), .nC(w5409), .C(w5465) );
	vdp_slatch g5508 (.D(w6254), .Q(w5416), .nC(w5410), .C(w5462) );
	vdp_slatch g5509 (.D(w5473), .Q(w5458), .nC(w5408), .C(w5461) );
	vdp_slatch g5510 (.D(w6253), .Q(w5420), .nC(w5417), .C(w5466) );
	vdp_slatch g5511 (.D(w6252), .Q(w5421), .nC(w5409), .C(w5465) );
	vdp_slatch g5512 (.D(w6251), .Q(w5422), .nC(w5410), .C(w5462) );
	vdp_slatch g5513 (.D(w5472), .Q(w5415), .nC(w5408), .C(w5461) );
	vdp_slatch g5514 (.D(w6250), .Q(w5426), .nC(w5417), .C(w5466) );
	vdp_slatch g5515 (.D(w6249), .Q(w5425), .nC(w5409), .C(w5465) );
	vdp_slatch g5516 (.D(w6248), .Q(w5427), .nC(w5410), .C(w5462) );
	vdp_slatch g5517 (.D(w5471), .Q(w5428), .nC(w5408), .C(w5461) );
	vdp_slatch g5518 (.D(w6247), .Q(w5429), .nC(w5417), .C(w5466) );
	vdp_slatch g5519 (.D(w6246), .Q(w5430), .nC(w5409), .C(w5465) );
	vdp_slatch g5520 (.D(w6245), .Q(w5441), .nC(w5410), .C(w5462) );
	vdp_slatch g5521 (.D(w5470), .Q(w5431), .nC(w5408), .C(w5461) );
	vdp_slatch g5522 (.D(w6244), .Q(w5435), .nC(w5417), .C(w5466) );
	vdp_slatch g5523 (.D(w6243), .Q(w5436), .nC(w5409), .C(w5465) );
	vdp_slatch g5524 (.D(w6242), .Q(w5434), .nC(w5410), .C(w5462) );
	vdp_slatch g5525 (.D(w5469), .Q(w5433), .nC(w5408), .C(w5461) );
	vdp_slatch g5526 (.D(w6241), .Q(w5438), .nC(w5417), .C(w5466) );
	vdp_slatch g5527 (.D(w6240), .Q(w5440), .nC(w5409), .C(w5465) );
	vdp_slatch g5528 (.D(w6239), .Q(w5439), .nC(w5410), .C(w5462) );
	vdp_slatch g5529 (.D(w5468), .Q(w5432), .nC(w5408), .C(w5461) );
	vdp_slatch g5530 (.D(w6238), .Q(w5437), .nC(w5417), .C(w5466) );
	vdp_slatch g5531 (.D(w6237), .Q(w5442), .nC(w5409), .C(w5465) );
	vdp_slatch g5532 (.D(w6236), .nC(w5410), .C(w5462), .Q(w5454) );
	vdp_sr_bit g5533 (.Q(w5476), .D(w5477), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g5534 (.Q(w6178), .D(w5476), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g5535 (.Q(w5489), .D(w6178), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_comp_str g5536 (.nZ(w5479), .A(w5490), .Z(w5467) );
	vdp_comp_str g5537 (.nZ(w5482), .A(w5490), .Z(w5464) );
	vdp_comp_str g5538 (.nZ(w5484), .A(w5490), .Z(w5463) );
	vdp_dlatch_inv g5539 (.nQ(w5477), .D(w5485), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g5540 (.Z(w5460), .B(DCLK2), .A(w5489) );
	vdp_and g5541 (.Z(w5490), .B(DCLK2), .A(w5476) );
	vdp_and g5542 (.Z(w5491), .B(DCLK2), .A(w5477) );
	vdp_slatch g5543 (.Q(w6238), .D(w6262), .nC(w5479), .C(w5467) );
	vdp_slatch g5544 (.Q(w6237), .D(w6261), .nC(w5482), .C(w5464) );
	vdp_slatch g5545 (.Q(w6236), .D(w6260), .nC(w5484), .C(w5463) );
	vdp_slatch g5546 (.Q(w6241), .D(w6265), .nC(w5479), .C(w5467) );
	vdp_slatch g5547 (.Q(w6240), .D(w6264), .nC(w5482), .C(w5464) );
	vdp_slatch g5548 (.Q(w6239), .D(w6263), .nC(w5484), .C(w5463) );
	vdp_slatch g5549 (.Q(w6244), .D(w6268), .nC(w5479), .C(w5467) );
	vdp_slatch g5550 (.Q(w6243), .D(w6267), .nC(w5482), .C(w5464) );
	vdp_slatch g5551 (.Q(w6242), .D(w6266), .nC(w5484), .C(w5463) );
	vdp_slatch g5552 (.Q(w6247), .D(w6271), .nC(w5479), .C(w5467) );
	vdp_slatch g5553 (.Q(w6246), .D(w6270), .nC(w5482), .C(w5464) );
	vdp_slatch g5554 (.Q(w6245), .D(w6269), .nC(w5484), .C(w5463) );
	vdp_slatch g5555 (.Q(w6250), .D(w6274), .nC(w5479), .C(w5467) );
	vdp_slatch g5556 (.Q(w6249), .D(w6273), .nC(w5482), .C(w5464) );
	vdp_slatch g5557 (.Q(w6248), .D(w6272), .nC(w5484), .C(w5463) );
	vdp_slatch g5558 (.Q(w6253), .D(w6277), .nC(w5479), .C(w5467) );
	vdp_slatch g5559 (.Q(w6252), .D(w6276), .nC(w5482), .C(w5464) );
	vdp_slatch g5560 (.Q(w6251), .D(w6275), .nC(w5484), .C(w5463) );
	vdp_slatch g5561 (.Q(w6256), .D(w6280), .nC(w5479), .C(w5467) );
	vdp_slatch g5562 (.Q(w6255), .D(w6279), .nC(w5482), .C(w5464) );
	vdp_slatch g5563 (.Q(w6254), .D(w6278), .nC(w5484), .C(w5463) );
	vdp_slatch g5564 (.Q(w6259), .D(w6283), .nC(w5479), .C(w5467) );
	vdp_slatch g5565 (.Q(w6258), .D(w6282), .nC(w5482), .C(w5464) );
	vdp_slatch g5566 (.Q(w6257), .D(w6281), .nC(w5484), .C(w5463) );
	vdp_sr_bit g5567 (.Q(w5488), .D(w5487), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_dlatch_inv g5568 (.nQ(w5487), .D(w5486), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g5569 (.Z(w5497), .B(w5487), .A(DCLK2) );
	vdp_nand g5570 (.Z(w5486), .B(w5394), .A(HCLK1) );
	vdp_nand g5571 (.Z(w5485), .B(w5404), .A(HCLK1) );
	vdp_and g5572 (.Z(w5496), .B(w5488), .A(DCLK2) );
	vdp_comp_str g5573 (.nZ(w5483), .A(w5497), .Z(w5495) );
	vdp_comp_str g5574 (.nZ(w5481), .A(w5496), .Z(w5494) );
	vdp_comp_str g5575 (.nZ(w5480), .A(w5491), .Z(w5493) );
	vdp_comp_str g5576 (.nZ(w5478), .A(w5490), .Z(w5492) );
	vdp_slatch g5577 (.D(S[7]), .Q(w5475), .nC(w5478), .C(w5492) );
	vdp_slatch g5578 (.D(S[7]), .Q(w6283), .nC(w5480), .C(w5493) );
	vdp_slatch g5579 (.D(S[7]), .Q(w6282), .nC(w5481), .C(w5494) );
	vdp_slatch g5580 (.D(S[7]), .Q(w6281), .nC(w5483), .C(w5495) );
	vdp_slatch g5581 (.D(S[5]), .Q(w5474), .nC(w5478), .C(w5492) );
	vdp_slatch g5582 (.D(S[5]), .Q(w6280), .nC(w5480), .C(w5493) );
	vdp_slatch g5583 (.D(S[5]), .Q(w6279), .nC(w5481), .C(w5494) );
	vdp_slatch g5584 (.D(S[5]), .Q(w6278), .nC(w5483), .C(w5495) );
	vdp_slatch g5585 (.D(S[3]), .Q(w5473), .nC(w5478), .C(w5492) );
	vdp_slatch g5586 (.D(S[3]), .Q(w6277), .nC(w5480), .C(w5493) );
	vdp_slatch g5587 (.D(S[3]), .Q(w6276), .nC(w5481), .C(w5494) );
	vdp_slatch g5588 (.D(S[3]), .Q(w6275), .nC(w5483), .C(w5495) );
	vdp_slatch g5589 (.D(S[1]), .Q(w5472), .nC(w5478), .C(w5492) );
	vdp_slatch g5590 (.D(S[1]), .Q(w6274), .nC(w5480), .C(w5493) );
	vdp_slatch g5591 (.D(S[1]), .Q(w6273), .nC(w5481), .C(w5494) );
	vdp_slatch g5592 (.D(S[1]), .Q(w6272), .nC(w5483), .C(w5495) );
	vdp_slatch g5593 (.D(S[6]), .Q(w5471), .nC(w5478), .C(w5492) );
	vdp_slatch g5594 (.D(S[6]), .Q(w6271), .nC(w5480), .C(w5493) );
	vdp_slatch g5595 (.D(S[6]), .Q(w6270), .nC(w5481), .C(w5494) );
	vdp_slatch g5596 (.D(S[6]), .Q(w6269), .nC(w5483), .C(w5495) );
	vdp_slatch g5597 (.D(S[4]), .Q(w5470), .nC(w5478), .C(w5492) );
	vdp_slatch g5598 (.D(S[4]), .Q(w6268), .nC(w5480), .C(w5493) );
	vdp_slatch g5599 (.D(S[4]), .Q(w6267), .nC(w5481), .C(w5494) );
	vdp_slatch g5600 (.D(S[4]), .Q(w6266), .nC(w5483), .C(w5495) );
	vdp_slatch g5601 (.D(S[2]), .Q(w5469), .nC(w5478), .C(w5492) );
	vdp_slatch g5602 (.D(S[2]), .Q(w6265), .nC(w5480), .C(w5493) );
	vdp_slatch g5603 (.D(S[2]), .Q(w6264), .nC(w5481), .C(w5494) );
	vdp_slatch g5604 (.D(S[2]), .Q(w6263), .nC(w5483), .C(w5495) );
	vdp_slatch g5605 (.D(S[0]), .Q(w5468), .nC(w5478), .C(w5492) );
	vdp_slatch g5606 (.D(S[0]), .Q(w6262), .nC(w5480), .C(w5493) );
	vdp_slatch g5607 (.D(S[0]), .Q(w6261), .nC(w5481), .C(w5494) );
	vdp_slatch g5608 (.D(S[0]), .nC(w5483), .C(w5495), .Q(w6260) );
	vdp_aon21_sr g5609 (.Q(w5551), .A1(w5123), .A2(w6443), .B(w6597), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5610 (.Q(w6597), .A1(w5120), .A2(w6443), .B(w6598), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5611 (.Q(w6598), .A1(w5118), .A2(w6443), .B(w6599), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5612 (.Q(w6599), .A1(w5536), .A2(w6443), .B(w6600), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5613 (.Q(w6600), .A1(w5546), .A2(w6443), .B(w6601), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5614 (.Q(w6601), .A1(w5513), .A2(w6443), .B(w6602), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5615 (.Q(w6602), .A1(w5515), .A2(w6443), .B(w6603), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5616 (.Q(w6603), .A1(w5505), .A2(w6443), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5617 (.Q(w6604), .A1(w5510), .A2(w6444), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5618 (.Q(w6605), .A1(w5516), .A2(w6444), .B(w6604), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5619 (.Q(w6606), .A1(w5514), .A2(w6444), .B(w6605), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5620 (.Q(w6607), .A1(w5553), .A2(w6444), .B(w6606), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5621 (.Q(w6608), .A1(w5537), .A2(w6444), .B(w6607), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5622 (.Q(w6609), .A1(w5119), .A2(w6444), .B(w6608), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5623 (.Q(w6610), .A1(w5121), .A2(w6444), .B(w6609), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5624 (.Q(w5556), .A1(w5122), .A2(w6444), .B(w6610), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5625 (.Q(w5561), .A1(w5507), .A2(w6445), .B(w6611), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5626 (.Q(w6611), .A1(w5504), .A2(w6445), .B(w6612), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5627 (.Q(w6612), .A1(w5503), .A2(w6445), .B(w6613), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5628 (.Q(w6613), .A1(w5509), .A2(w6445), .B(w6614), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5629 (.Q(w6614), .A1(w5512), .A2(w6445), .B(w6615), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5630 (.Q(w6615), .A1(w5517), .A2(w6445), .B(w6616), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5631 (.Q(w6616), .A1(w5529), .A2(w6445), .B(w6617), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5632 (.Q(w6617), .A1(w5532), .A2(w6445), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_or4 g5633 (.Z(w5542), .B(w5546), .A(w5194), .C(w5553), .D(w5512) );
	vdp_or4 g5634 (.Z(w5197), .B(w5536), .A(w5192), .C(w5537), .D(w5509) );
	vdp_aon22 g5635 (.Z(w5525), .B2(w4361), .B1(w5530), .A1(w5566), .A2(DB[0]) );
	vdp_aon22 g5636 (.Z(w5524), .B2(w4362), .B1(w5530), .A1(w5566), .A2(DB[1]) );
	vdp_aon22 g5637 (.Z(w5523), .B2(w4370), .B1(w5530), .A1(w5566), .A2(DB[2]) );
	vdp_aon22 g5638 (.Z(w5522), .B2(w4361), .B1(w5530), .A1(w5566), .A2(DB[8]) );
	vdp_aon22 g5639 (.Z(w5521), .B2(w4362), .B1(w5530), .A1(w5566), .A2(DB[9]) );
	vdp_aon22 g5640 (.Z(w5520), .B2(w4370), .B1(w5530), .A1(w5566), .A2(DB[10]) );
	vdp_or4 g5641 (.Z(w5552), .B(w5501), .A(w5502), .C(w5534), .D(w5535) );
	vdp_or4 g5642 (.Z(w5543), .B(w5540), .A(w5541), .C(w5539), .D(w5538) );
	vdp_or4 g5643 (.Z(w5560), .B(w5515), .A(w5186), .C(w5516), .D(w5529) );
	vdp_or4 g5644 (.Z(w5557), .B(w5514), .A(w5517), .C(w5513), .D(w5511) );
	vdp_or4 g5645 (.Z(w5567), .B(w5506), .A(w5508), .C(w5519), .D(w5518) );
	vdp_or4 g5646 (.Z(w5558), .B(w5527), .A(w5528), .C(w5533), .D(w5526) );
	vdp_or4 g5647 (.Z(w5569), .B(w5505), .A(w5187), .C(w5510), .D(w5532) );
	vdp_comp_we g5648 (.nZ(w5530), .A(w114), .Z(w5566) );
	vdp_not g5649 (.nZ(w6443), .A(w5167) );
	vdp_not g5650 (.nZ(w6444), .A(w5167) );
	vdp_not g5651 (.nZ(w6445), .A(w5167) );
	vdp_slatch g5652 (.Q(w5538), .D(w5583), .nC(w5549), .C(w5582) );
	vdp_comp_str g5653 (.nZ(w5549), .A(w5207), .Z(w5582) );
	vdp_slatch g5654 (.Q(w5539), .D(w5585), .nC(w5549), .C(w5582) );
	vdp_slatch g5655 (.Q(w5540), .D(w5586), .nC(w5549), .C(w5582) );
	vdp_slatch g5656 (.Q(w5541), .D(w5587), .nC(w5549), .C(w5582) );
	vdp_slatch g5657 (.Q(w5502), .D(w5588), .nC(w5549), .C(w5582) );
	vdp_slatch g5658 (.Q(w5501), .D(w5590), .nC(w5549), .C(w5582) );
	vdp_slatch g5659 (.Q(w5534), .D(w5591), .nC(w5549), .C(w5582) );
	vdp_slatch g5660 (.Q(w5535), .D(w5592), .nC(w5549), .C(w5582) );
	vdp_slatch g5661 (.Q(w5526), .D(w5601), .nC(w5564), .C(w5600) );
	vdp_comp_str g5662 (.nZ(w5564), .A(w5207), .Z(w5600) );
	vdp_slatch g5663 (.Q(w5533), .D(w5603), .nC(w5564), .C(w5600) );
	vdp_slatch g5664 (.Q(w5527), .D(w5604), .nC(w5564), .C(w5600) );
	vdp_slatch g5665 (.Q(w5528), .D(w5605), .nC(w5564), .C(w5600) );
	vdp_slatch g5666 (.Q(w5508), .D(w5606), .nC(w5564), .C(w5600) );
	vdp_slatch g5667 (.Q(w5506), .D(w5608), .nC(w5564), .C(w5600) );
	vdp_slatch g5668 (.Q(w5519), .D(w5609), .nC(w5564), .C(w5600) );
	vdp_slatch g5669 (.Q(w5518), .D(w5610), .nC(w5564), .C(w5600) );
	vdp_comp_we g5670 (.nZ(w5545), .A(1'b0), .Z(w5195) );
	vdp_aon22 g5671 (.Z(w5612), .B2(w5545), .B1(w5568), .A1(w5567), .A2(w5195) );
	vdp_not g5672 (.nZ(w5167), .A(w4372) );
	vdp_not g5673 (.nZ(w5568), .A(w5569) );
	vdp_not g5674 (.nZ(w5559), .A(w5560) );
	vdp_not g5675 (.nZ(w5555), .A(w5557) );
	vdp_not g5676 (.nZ(w5544), .A(w5542) );
	vdp_and3 g5677 (.Z(w5572), .B(w5571), .A(w5543), .C(w5542) );
	vdp_aon22 g5678 (.Z(w5580), .B2(w5545), .B1(w5544), .A1(w5543), .A2(w5195) );
	vdp_notif0 g5679 (.A(w5547), .nZ(DB[4]), .nE(w5548) );
	vdp_aon2222 g5680 (.Z(w5547), .B2(w5546), .B1(w5578), .A1(w5579), .A2(w5515), .D2(w5123), .D1(w5576), .C1(w5577), .C2(w5118) );
	vdp_notif0 g5681 (.A(w5550), .nZ(DB[12]), .nE(w5548) );
	vdp_aon2222 g5682 (.Z(w5550), .B2(w5513), .B1(w5578), .A1(w5579), .A2(w5505), .D2(w5120), .D1(w5576), .C1(w5577), .C2(w5536) );
	vdp_notif0 g5683 (.A(w6213), .nZ(DB[13]), .nE(w5548) );
	vdp_aon2222 g5684 (.Z(w6213), .B2(w5514), .B1(w5578), .A1(w5579), .A2(w5510), .D2(w5121), .D1(w5576), .C1(w5577), .C2(w5537) );
	vdp_notif0 g5685 (.A(w5554), .nZ(DB[5]), .nE(w5548) );
	vdp_aon2222 g5686 (.Z(w5554), .B2(w5553), .B1(w5578), .A1(w5579), .A2(w5516), .D2(w5122), .D1(w5576), .C1(w5577), .C2(w5119) );
	vdp_notif0 g5687 (.A(w5563), .nZ(DB[14]), .nE(w5548) );
	vdp_aon2222 g5688 (.Z(w5563), .B2(w5517), .B1(w5578), .A1(w5579), .A2(w5532), .D2(w5504), .D1(w5576), .C1(w5577), .C2(w5509) );
	vdp_notif0 g5689 (.A(w5562), .nZ(DB[6]), .nE(w5548) );
	vdp_aon2222 g5690 (.Z(w5562), .B2(w5512), .B1(w5578), .A1(w5579), .A2(w5529), .D2(w5507), .D1(w5576), .C1(w5577), .C2(w5503) );
	vdp_aon22 g5691 (.Z(w5593), .B2(w5545), .B1(w5555), .A1(w5552), .A2(w5195) );
	vdp_aon22 g5692 (.Z(w5596), .B2(w5545), .B1(w5559), .A1(w5558), .A2(w5195) );
	vdp_and3 g5693 (.Z(w5574), .B(w5595), .A(w5552), .C(w5557) );
	vdp_and3 g5694 (.Z(w5575), .B(w5597), .A(w5558), .C(w5560) );
	vdp_and3 g5695 (.Z(w5573), .B(w5611), .A(w5567), .C(w5569) );
	vdp_not g5696 (.nZ(w5548), .A(w115) );
	vdp_slatch g5697 (.Q(w5606), .D(w5268), .nC(w5640), .C(w5607) );
	vdp_slatch g5698 (.Q(w5608), .D(w5271), .nC(w5640), .C(w5607) );
	vdp_slatch g5699 (.Q(w5609), .D(w5272), .nC(w5640), .C(w5607) );
	vdp_slatch g5700 (.Q(w5610), .D(w5274), .nC(w5640), .C(w5607) );
	vdp_comp_str g5701 (.nZ(w5640), .A(w5641), .Z(w5607) );
	vdp_slatch g5702 (.Q(w5601), .D(w5255), .nC(w5635), .C(w5602) );
	vdp_slatch g5703 (.Q(w5603), .D(w5259), .nC(w5635), .C(w5602) );
	vdp_slatch g5704 (.Q(w5604), .D(w5260), .nC(w5635), .C(w5602) );
	vdp_slatch g5705 (.Q(w5605), .D(w5263), .nC(w5635), .C(w5602) );
	vdp_comp_str g5706 (.nZ(w5635), .A(w5639), .Z(w5602) );
	vdp_slatch g5707 (.Q(w5588), .D(w5268), .nC(w5622), .C(w5589) );
	vdp_slatch g5708 (.Q(w5590), .D(w5271), .nC(w5622), .C(w5589) );
	vdp_slatch g5709 (.Q(w5591), .D(w5272), .nC(w5622), .C(w5589) );
	vdp_slatch g5710 (.Q(w5592), .D(w5274), .nC(w5622), .C(w5589) );
	vdp_comp_str g5711 (.nZ(w5622), .A(w6440), .Z(w5589) );
	vdp_slatch g5712 (.Q(w5583), .D(w5255), .nC(w5621), .C(w5584) );
	vdp_slatch g5713 (.Q(w5585), .D(w5259), .nC(w5621), .C(w5584) );
	vdp_slatch g5714 (.Q(w5586), .D(w5260), .nC(w5621), .C(w5584) );
	vdp_slatch g5715 (.Q(w5587), .D(w5263), .nC(w5621), .C(w5584) );
	vdp_comp_str g5716 (.nZ(w5621), .A(w5619), .Z(w5584) );
	vdp_dlatch_inv g5717 (.nQ(w6212), .D(w5614), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5718 (.Z(w5616), .B(w5246), .A(w6212) );
	vdp_sr_bit g5719 (.Q(COLLISION), .D(w6209), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g5720 (.Q(w5613), .D(w5551), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5721 (.nQ(w5618), .D(w5581), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5722 (.nQ(w6204), .D(w5594), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5723 (.nQ(w6206), .D(w5628), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5724 (.Z(w6205), .B(w6206), .A(w5246) );
	vdp_sr_bit g5725 (.Q(w6215), .D(w5556), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5726 (.nQ(w5598), .D(w6438), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5727 (.Z(w6207), .B(w5598), .A(w5246) );
	vdp_sr_bit g5728 (.Q(w5632), .D(w5561), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5729 (.nQ(w5629), .D(w6211), .nC(nDCLK2), .C(DCLK2) );
	vdp_not g5730 (.nZ(w5645), .A(w5246) );
	vdp_not g5731 (.nZ(w5599), .A(w75) );
	vdp_not g5732 (.nZ(w5633), .A(w74) );
	vdp_dlatch_inv g5733 (.nQ(w5643), .D(w6208), .nC(nDCLK2), .C(DCLK2) );
	vdp_and g5734 (.Z(w5611), .B(w5645), .A(w5247) );
	vdp_aoi21 g5735 (.Z(w6208), .B(w5630), .A1(w5612), .A2(w5611) );
	vdp_and g5736 (.Z(w5498), .B(w5643), .A(DCLK1) );
	vdp_and g5737 (.Z(w5499), .B(w5629), .A(DCLK1) );
	vdp_and g5738 (.Z(w5597), .B(w6207), .A(w5247) );
	vdp_aoi21 g5739 (.Z(w6211), .B(w5630), .A1(w5596), .A2(w5597) );
	vdp_and g5740 (.Z(w5595), .B(w6205), .A(w5247) );
	vdp_aoi21 g5741 (.Z(w5594), .B(w5617), .A1(w5593), .A2(w5595) );
	vdp_and g5742 (.Z(w5571), .B(w5247), .A(w5616) );
	vdp_aoi21 g5743 (.Z(w5581), .B(w5617), .A1(w5580), .A2(w5571) );
	vdp_and g5744 (.Z(w5531), .B(DCLK1), .A(w5618) );
	vdp_and g5745 (.Z(w5500), .B(w6204), .A(DCLK1) );
	vdp_and g5746 (.Z(w5576), .B(w5599), .A(w5633) );
	vdp_and g5747 (.Z(w5578), .B(w75), .A(w5633) );
	vdp_and g5748 (.Z(w5577), .B(w5599), .A(w74) );
	vdp_and g5749 (.Z(w5579), .B(w75), .A(w74) );
	vdp_or8 g5750 (.Z(w6209), .B(w5572), .A(w5241), .C(w5573), .D(w6210), .F(w5575), .E(w5570), .G(w5225), .H(w5574) );
	vdp_sr_bit g5751 (.Q(w5302), .D(w5650), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5752 (.Q(w5615), .D(w5302), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5753 (.Q(w5301), .D(w5627), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5754 (.Q(w5646), .D(w5301), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5755 (.Q(w5320), .D(w6193), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5756 (.Q(w5634), .D(w5320), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_comp_we g5757 (.nZ(w5648), .A(M5), .Z(w5647) );
	vdp_not g5758 (.nZ(w5641), .A(w5642) );
	vdp_or g5759 (.Z(w5324), .B(w5644), .A(w5266) );
	vdp_and3 g5760 (.Z(w5644), .B(w5316), .A(w5323), .C(w5315) );
	vdp_and3 g5761 (.Z(w5637), .B(w5316), .A(w5323), .C(w5327) );
	vdp_and3 g5762 (.Z(w6438), .B(w5321), .A(w5310), .C(w5322) );
	vdp_and3 g5763 (.Z(w5624), .B(w5328), .A(w5323), .C(w5315) );
	vdp_and3 g5764 (.Z(w5626), .B(w5328), .A(w5323), .C(w5327) );
	vdp_aoi21 g5765 (.Z(w5614), .B(w5256), .A1(w5245), .A2(w5326) );
	vdp_aon22 g5766 (.Z(w5650), .B2(w5551), .B1(w5648), .A1(w5647), .A2(w5613) );
	vdp_aon22 g5767 (.Z(w5627), .B2(w5556), .B1(w5648), .A1(w5647), .A2(w6215) );
	vdp_aon22 g5768 (.Z(w6193), .B2(w5561), .B1(w5648), .A1(w5647), .A2(w5632) );
	vdp_bufif0 g5769 (.A(w5646), .Z(COL[2]), .nE(w5649) );
	vdp_oai21 g5770 (.Z(w5625), .B(DCLK2), .A1(w5638), .A2(w5626) );
	vdp_and g5771 (.Z(w5628), .B(w5321), .A(w5310) );
	vdp_or g5772 (.Z(w5638), .B(w5624), .A(w5266) );
	vdp_bufif0 g5773 (.A(w5634), .Z(COL[3]), .nE(w5649) );
	vdp_oai21 g5774 (.Z(w5636), .B(DCLK2), .A1(w5638), .A2(w5637) );
	vdp_oai21 g5775 (.Z(w5642), .B(DCLK2), .A1(w5637), .A2(w5324) );
	vdp_not g5776 (.nZ(w5327), .A(w5315) );
	vdp_not g5777 (.nZ(w5639), .A(w5636) );
	vdp_not g5778 (.nZ(w5325), .A(w74) );
	vdp_not g5779 (.nZ(w5328), .A(w5316) );
	vdp_not g5780 (.nZ(w6440), .A(w5625) );
	vdp_not g5781 (.nZ(w5326), .A(w5322) );
	vdp_not g5782 (.nZ(w5619), .A(w5620) );
	vdp_bufif0 g5783 (.A(w5615), .Z(COL[1]), .nE(w5649) );
	vdp_oai21 g5784 (.Z(w5620), .B(DCLK2), .A1(w5308), .A2(w5626) );
	vdp_not g5785 (.nZ(w5649), .A(SPR_PRIO) );
	vdp_nand3 g5786 (.Z(w5623), .B(w105), .A(w75), .C(w5325) );
	vdp_nand g5787 (.Z(w5617), .B(w5319), .A(w5623) );
	vdp_nand3 g5788 (.Z(w5631), .B(w105), .A(w75), .C(w74) );
	vdp_nand g5789 (.Z(w5630), .B(w5319), .A(w5631) );
	vdp_sr_bit g5790 (.Q(w5673), .D(w5714), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5791 (.Q(w5674), .D(w5712), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5792 (.Q(w5671), .D(w5719), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5793 (.Q(w5672), .D(w5711), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5794 (.Z(w4367), .B2(w5673), .B1(w5708), .A1(w5707), .A2(w73), .C1(w5662), .C2(w5674) );
	vdp_aon222 g5795 (.Z(w4366), .B2(w5671), .B1(w5708), .A1(w5707), .A2(w72), .C1(w5662), .C2(w5672) );
	vdp_sr_bit g5796 (.Q(w5669), .D(w5718), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5797 (.Q(w5670), .D(w5710), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5798 (.Z(w4365), .B2(w5669), .B1(w5708), .A1(w5707), .A2(w71), .C1(w5662), .C2(w5670) );
	vdp_sr_bit g5799 (.Q(w5667), .D(w5717), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5800 (.Q(w5668), .D(w5709), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5801 (.Z(w4364), .B2(w5667), .B1(w5708), .A1(w5707), .A2(w70), .C1(w5662), .C2(w5668) );
	vdp_sr_bit g5802 (.Q(w5663), .D(w5716), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5803 (.Q(w5666), .D(w5720), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5804 (.Z(w4363), .B2(w5663), .B1(w5708), .A1(w5707), .A2(w69), .C1(w5662), .C2(w5666) );
	vdp_sr_bit g5805 (.Q(w5664), .D(w5715), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5806 (.Q(w5665), .D(w5706), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5807 (.Z(w4368), .B2(w5664), .B1(w5708), .A1(w5707), .A2(w68), .C1(w5662), .C2(w5665) );
	vdp_sr_bit g5808 (.Q(w5310), .D(w6417), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_slatch g5809 (.Q(w6417), .D(w5400), .nC(w5698), .C(w5659) );
	vdp_sr_bit g5810 (.Q(w5321), .D(w6415), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_slatch g5811 (.Q(w6415), .D(w5380), .nC(w5698), .C(w5659) );
	vdp_sr_bit g5812 (.Q(w5322), .D(w6416), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_slatch g5813 (.Q(w6416), .D(w5388), .nC(w5698), .C(w5659) );
	vdp_sr_bit g5814 (.Q(w5675), .D(w25), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5815 (.Q(w5658), .D(w5675), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5816 (.Q(w5657), .D(w5703), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5817 (.Q(w5691), .D(w5701), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5818 (.Q(w5690), .D(w5700), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5819 (.Q(w5654), .D(w4372), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5820 (.Q(w5653), .D(w5686), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5821 (.Q(w5681), .D(w6218), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5822 (.Q(w6218), .D(w5722), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_xor g5823 (.Z(w5683), .B(w5681), .A(w5682) );
	vdp_dlatch_inv g5824 (.nQ(w5652), .D(w5686), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5825 (.nQ(w5684), .D(w5683), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5826 (.nQ(w5655), .D(w5656), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5827 (.nQ(w5689), .D(w5688), .nC(nHCLK1), .C(HCLK1) );
	vdp_comp_str g5828 (.nZ(w5698), .A(w5695), .Z(w5659) );
	vdp_oai21 g5829 (.Z(w6217), .B(w5685), .A1(w5722), .A2(w5681) );
	vdp_and g5830 (.Z(w4361), .B(w5679), .A(w5651) );
	vdp_not g5831 (.nZ(w5246), .A(w5684) );
	vdp_not g5832 (.nZ(w5686), .A(w6217) );
	vdp_and g5833 (.Z(w4362), .B(w5678), .A(w5651) );
	vdp_and g5834 (.Z(w4370), .B(w5677), .A(w5651) );
	vdp_or g5835 (.Z(w5687), .B(w5653), .A(w5686) );
	vdp_not g5836 (.nZ(w5705), .A(w114) );
	vdp_not g5837 (.nZ(w4372), .A(w5688) );
	vdp_not g5838 (.nZ(w5721), .A(M5) );
	vdp_not g5839 (.nZ(w5708), .A(w6408) );
	vdp_not g5840 (.nZ(w5660), .A(w5659) );
	vdp_not g5841 (.nZ(w5707), .A(w5705) );
	vdp_not g5842 (.nZ(w5662), .A(w5661) );
	vdp_or4 g5843 (.Z(w4369), .B(w4372), .A(w114), .C(w5654), .D(w5687) );
	vdp_or4 g5844 (.Z(w5688), .B(w5691), .A(w5651), .C(w5657), .D(w5690) );
	vdp_nand g5845 (.Z(w5656), .B(w5689), .A(HCLK2) );
	vdp_nand g5846 (.Z(w5319), .B(w5705), .A(w5655) );
	vdp_nor g5847 (.Z(w5247), .B(w5652), .A(w114) );
	vdp_nand g5848 (.Z(w5661), .B(w5705), .A(w5660) );
	vdp_nand g5849 (.Z(w6408), .B(w5705), .A(w5651) );
	vdp_aoi22 g5850 (.Z(w5651), .B2(w5721), .B1(w25), .A1(M5), .A2(w5658) );
	vdp_cnt_bit_load g5851 (.Q(w5750), .D(w5699), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w38), .CI(w5807), .L(w5697), .nL(w5743) );
	vdp_cnt_bit_load g5852 (.Q(w5696), .D(w5747), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w38), .CI(w5692), .L(w5697), .nL(w5743), .CO(w5807) );
	vdp_sr_bit g5853 (.Q(w5685), .D(w6200), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5854 (.SUM(w5703), .CO(w6396), .CI(1'b1), .A(HPOS[0]), .B(M5) );
	vdp_fa g5855 (.SUM(w5701), .CO(w6397), .CI(w6396), .A(HPOS[1]), .B(1'b0) );
	vdp_fa g5856 (.SUM(w5700), .CO(w6398), .CI(w6397), .A(HPOS[2]), .B(1'b1) );
	vdp_fa g5857 (.SUM(w5706), .CO(w6399), .CI(w6398), .A(HPOS[3]), .B(M5) );
	vdp_fa g5858 (.SUM(w5720), .CO(w6400), .CI(w6399), .A(HPOS[4]), .B(w5758) );
	vdp_fa g5859 (.SUM(w5709), .CO(w6401), .CI(w6400), .A(HPOS[5]), .B(1'b1) );
	vdp_fa g5860 (.SUM(w5710), .CO(w6402), .CI(w6401), .A(HPOS[6]), .B(1'b1) );
	vdp_fa g5861 (.SUM(w5711), .CO(w6403), .CI(w6402), .A(HPOS[7]), .B(1'b1) );
	vdp_fa g5862 (.SUM(w5712), .CI(w6403), .A(HPOS[8]), .B(1'b1) );
	vdp_not g5863 (.nZ(w5758), .A(M5) );
	vdp_aoi33 g5864 (.Z(w6200), .B2(w6414), .B1(w5714), .A1(H40), .A2(w5714), .A3(w5713), .B3(w6414) );
	vdp_not g5865 (.nZ(w6414), .A(H40) );
	vdp_or g5866 (.Z(w5713), .B(w5718), .A(w5719) );
	vdp_and g5867 (.Z(w5694), .B(w5692), .A(w5693) );
	vdp_sr_bit g5868 (.Q(w5692), .D(w6216), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5869 (.Q(w6216), .D(w5443), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5870 (.nQ(w5740), .D(w5297), .nC(nDCLK2), .C(DCLK2) );
	vdp_slatch g5871 (.Q(w5739), .D(w5726), .nC(w5680), .C(w5730) );
	vdp_slatch g5872 (.Q(w5679), .D(w5739), .nC(w5676), .C(w5732) );
	vdp_slatch g5873 (.Q(w5733), .D(w5724), .nC(w5680), .C(w5730) );
	vdp_slatch g5874 (.Q(w5677), .D(w5733), .nC(w5676), .C(w5732) );
	vdp_slatch g5875 (.Q(w5734), .D(w5725), .nC(w5680), .C(w5730) );
	vdp_slatch g5876 (.Q(w5678), .D(w5734), .nC(w5676), .C(w5732) );
	vdp_slatch g5877 (.Q(w6219), .D(w5448), .nC(w5680), .C(w5730) );
	vdp_sr_bit g5878 (.Q(w5682), .D(w6219), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_and g5879 (.Z(w5723), .B(DCLK2), .A(w5297) );
	vdp_comp_str g5880 (.nZ(w5676), .A(w5723), .Z(w5732) );
	vdp_comp_str g5881 (.nZ(w5680), .A(w5695), .Z(w5730) );
	vdp_not g5882 (.nZ(w5722), .A(w5740) );
	vdp_comp_we g5883 (.nZ(w5743), .A(w5694), .Z(w5697) );
	vdp_and3 g5884 (.Z(w5695), .B(HCLK1), .A(w5693), .C(w5692) );
	vdp_nand g5885 (.Z(w5747), .B(w5728), .A(M5) );
	vdp_nand g5886 (.Z(w5699), .B(w5727), .A(M5) );
	vdp_nor g5887 (.Z(w5693), .B(w5750), .A(w5696) );
	vdp_fa g5888 (.SUM(w5714), .CI(w5768), .A(w5767), .B(w5778) );
	vdp_aon22 g5889 (.Z(w5767), .B2(w5770), .B1(w5766), .A1(w5801), .A2(w5736) );
	vdp_sr_bit g5890 (.Q(w5766), .D(w5714), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5891 (.Q(w5801), .D(w5802), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5892 (.SUM(w5802), .CI(w5764), .A(w5765), .B(w5797) );
	vdp_aon22 g5893 (.Z(w5765), .B2(w5775), .B1(w5800), .A1(1'b0), .A2(w5729) );
	vdp_fa g5894 (.SUM(w5719), .CO(w5768), .CI(w5763), .A(w5762), .B(w5778) );
	vdp_aon22 g5895 (.Z(w5762), .B2(w5770), .B1(w5761), .A1(w5798), .A2(w5736) );
	vdp_sr_bit g5896 (.Q(w5761), .D(w5719), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5897 (.Q(w5798), .D(w5804), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5898 (.SUM(w5804), .CO(w5764), .CI(w5760), .A(w5759), .B(w5797) );
	vdp_aon22 g5899 (.Z(w5759), .B2(w5775), .B1(w5795), .A1(w5796), .A2(w5729) );
	vdp_fa g5900 (.SUM(w5718), .CO(w5763), .CI(w5757), .A(w5756), .B(w5778) );
	vdp_aon22 g5901 (.Z(w5756), .B2(w5770), .B1(w5755), .A1(w5794), .A2(w5736) );
	vdp_fa g5902 (.SUM(w5805), .CO(w5760), .CI(w5754), .A(w5753), .B(w5781) );
	vdp_aon22 g5903 (.Z(w5753), .B2(w5775), .B1(w5792), .A1(w5793), .A2(w5729) );
	vdp_sr_bit g5904 (.Q(w5755), .D(w5718), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5905 (.Q(w5794), .D(w5805), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5906 (.SUM(w5717), .CO(w5757), .CI(w5769), .A(w5752), .B(w5778) );
	vdp_aon22 g5907 (.Z(w5752), .B2(w5770), .B1(w5751), .A1(w5791), .A2(w5736) );
	vdp_sr_bit g5908 (.Q(w5751), .D(w5717), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5909 (.Q(w5791), .D(w5790), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5910 (.SUM(w5790), .CO(w5754), .CI(w5748), .A(w5749), .B(w5781) );
	vdp_aon22 g5911 (.Z(w5749), .B2(w5775), .B1(w6411), .A1(w5789), .A2(w5729) );
	vdp_fa g5912 (.SUM(w5716), .CO(w5769), .CI(w5745), .A(w5746), .B(w5778) );
	vdp_aon22 g5913 (.Z(w5746), .B2(w5770), .B1(w5744), .A1(w5788), .A2(w5736) );
	vdp_sr_bit g5914 (.Q(w5744), .D(w5716), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5915 (.Q(w5788), .D(w6404), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5916 (.SUM(w6404), .CO(w5748), .CI(w5742), .A(w5741), .B(w5787) );
	vdp_aon22 g5917 (.Z(w5741), .B2(w5775), .B1(w5806), .A1(w5786), .A2(w5729) );
	vdp_fa g5918 (.SUM(w5715), .CO(w5745), .CI(w5738), .A(w5737), .B(w5778) );
	vdp_aon22 g5919 (.Z(w5737), .B2(w5770), .B1(w5735), .A1(w5785), .A2(w5736) );
	vdp_sr_bit g5920 (.Q(w5735), .D(w5715), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5921 (.Q(w5785), .D(w5784), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5922 (.SUM(w5784), .CO(w5742), .CI(w5448), .A(w5731), .B(w5780) );
	vdp_aon22 g5923 (.Z(w5731), .B2(w5775), .B1(w5782), .A1(w5783), .A2(w5729) );
	vdp_aon22 g5924 (.Z(w5400), .B2(w5775), .B1(w5779), .A1(w5803), .A2(w5729) );
	vdp_aon22 g5925 (.Z(w5380), .B2(w5775), .B1(w5774), .A1(w5777), .A2(w5729) );
	vdp_aon22 g5926 (.Z(w5388), .B2(w5775), .B1(w5773), .A1(w5776), .A2(w5729) );
	vdp_and g5927 (.Z(w5738), .B(w5772), .A(w6410) );
	vdp_comp_we g5928 (.nZ(w5729), .A(M5), .Z(w5775) );
	vdp_comp_we g5929 (.nZ(w5770), .A(w6409), .Z(w5736) );
	vdp_sr_bit g5930 (.Q(w6409), .D(w5695), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5931 (.Q(w5771), .D(w5740), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5932 (.Q(w5817), .D(w5820), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5933 (.Q(w5820), .D(w5821), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5934 (.Q(w5821), .D(w5825), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5935 (.Q(w5825), .D(w5826), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5936 (.Q(w5826), .D(w5827), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5937 (.nQ(w5827), .D(w5830), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5938 (.nZ(w5779), .A(w5817) );
	vdp_sr_bit g5939 (.Q(w5831), .D(w5832), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5940 (.Q(w5832), .D(w5836), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5941 (.Q(w5836), .D(w5837), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5942 (.Q(w5837), .D(w5839), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5943 (.Q(w5839), .D(w5842), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5944 (.nQ(w5842), .D(w5841), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5945 (.nZ(w5782), .A(w5831) );
	vdp_sr_bit g5946 (.Q(w5843), .D(w6220), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5947 (.Q(w6220), .D(w5846), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5948 (.Q(w5846), .D(w5848), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5949 (.Q(w5848), .D(w5849), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5950 (.Q(w5849), .D(w5850), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5951 (.nQ(w5850), .D(w5854), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5952 (.nZ(w5806), .A(w5843) );
	vdp_sr_bit g5953 (.Q(w5855), .D(w5858), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5954 (.Q(w5858), .D(w5862), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5955 (.Q(w5862), .D(w5861), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5956 (.Q(w5861), .D(w5863), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5957 (.Q(w5863), .D(w5866), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5958 (.nQ(w5866), .D(w5867), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5959 (.nZ(w6411), .A(w5855) );
	vdp_sr_bit g5960 (.Q(w5870), .D(w5873), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5961 (.Q(w5873), .D(w5874), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5962 (.Q(w5874), .D(w5875), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5963 (.Q(w5875), .D(w5899), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5964 (.Q(w5899), .D(w5900), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5965 (.nQ(w5900), .D(w5880), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5966 (.nZ(w5792), .A(w5870) );
	vdp_sr_bit g5967 (.Q(w5901), .D(w5895), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5968 (.Q(w5895), .D(w5894), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5969 (.Q(w5894), .D(w5892), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5970 (.Q(w5892), .D(w5891), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5971 (.Q(w5891), .D(w5889), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5972 (.nQ(w5889), .D(w5879), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5973 (.nZ(w5795), .A(w5901) );
	vdp_sr_bit g5974 (.Q(w6412), .D(w5885), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5975 (.Q(w5885), .D(w5886), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5976 (.Q(w5886), .D(w5882), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5977 (.Q(w5882), .D(w5881), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5978 (.Q(w5881), .D(w5877), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5979 (.nQ(w5877), .D(w5878), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5980 (.nZ(w5800), .A(w6412) );
	vdp_and g5981 (.Z(w5778), .B(w5772), .A(w5682) );
	vdp_and g5982 (.Z(w5813), .B(w5448), .A(w5728) );
	vdp_and g5983 (.Z(w5814), .B(w5448), .A(w5727) );
	vdp_or g5984 (.Z(w5780), .B(w5813), .A(w5781) );
	vdp_and g5985 (.B(w5816), .A(M5), .Z(w5448) );
	vdp_or g5986 (.Z(w5787), .B(w5814), .A(w5781) );
	vdp_and g5987 (.Z(w5781), .B(w22), .A(w6421) );
	vdp_or g5988 (.Z(w5797), .B(w5781), .A(M5) );
	vdp_not g5989 (.nZ(w6421), .A(M5) );
	vdp_not g5990 (.nZ(w6410), .A(w5682) );
	vdp_nor g5991 (.Z(w5772), .B(w6409), .A(w5771) );
	vdp_sr_bit g5992 (.Q(w5829), .D(w5833), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5993 (.Q(w5833), .D(w5834), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5994 (.Q(w5834), .D(w5835), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5995 (.Q(w5835), .D(w5838), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5996 (.Q(w5838), .D(w6413), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5997 (.nQ(w6413), .D(w5907), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5998 (.nZ(w5725), .A(w5829) );
	vdp_sr_bit g5999 (.Q(w5818), .D(w5819), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6000 (.Q(w5819), .D(w5822), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6001 (.Q(w5822), .D(w5823), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6002 (.Q(w5823), .D(w5824), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6003 (.Q(w5824), .D(w5828), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6004 (.nQ(w5828), .D(w5906), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6005 (.nZ(w5726), .A(w5818) );
	vdp_sr_bit g6006 (.Q(w5808), .D(w5809), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6007 (.Q(w5809), .D(w5810), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6008 (.Q(w5810), .D(w5812), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6009 (.Q(w5812), .D(w5811), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6010 (.Q(w5811), .D(w5815), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6011 (.nQ(w5815), .D(w5905), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6012 (.nZ(w5816), .A(w5808) );
	vdp_sr_bit g6013 (.Q(w5840), .D(w5844), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6014 (.Q(w5844), .D(w5845), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6015 (.Q(w5845), .D(w5847), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6016 (.Q(w5847), .D(w5851), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6017 (.Q(w5851), .D(w5852), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6018 (.nQ(w5852), .D(w5912), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6019 (.nZ(w5724), .A(w5840) );
	vdp_sr_bit g6020 (.Q(w5853), .D(w5856), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6021 (.Q(w5856), .D(w5857), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6022 (.Q(w5857), .D(w5859), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6023 (.Q(w5859), .D(w5860), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6024 (.Q(w5860), .D(w5864), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6025 (.nQ(w5864), .D(w5908), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6026 (.nZ(w5728), .A(w5853) );
	vdp_sr_bit g6027 (.Q(w5865), .D(w5868), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6028 (.Q(w5868), .D(w5869), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6029 (.Q(w5869), .D(w5871), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6030 (.Q(w5871), .D(w5872), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6031 (.Q(w5872), .D(w5876), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6032 (.nQ(w5876), .D(w5909), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6033 (.nZ(w5727), .A(w5865) );
	vdp_sr_bit g6034 (.Q(w5897), .D(w5898), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6035 (.Q(w5898), .D(w5902), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6036 (.Q(w5902), .D(w5903), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6037 (.Q(w5903), .D(w5896), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6038 (.Q(w5896), .D(w5893), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6039 (.nQ(w5893), .D(w5910), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6040 (.nZ(w5773), .A(w5897) );
	vdp_sr_bit g6041 (.Q(w5888), .D(w5890), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6042 (.Q(w5890), .D(w5887), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6043 (.Q(w5887), .D(w5884), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6044 (.Q(w5884), .D(w5883), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6045 (.Q(w5883), .D(w5904), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6046 (.nQ(w5904), .D(w5911), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6047 (.nZ(w5774), .A(w5888) );
	vdp_slatch g6048 (.D(w5937), .nC(w5974), .C(w5915), .nQ(w5776) );
	vdp_slatch g6049 (.D(S[1]), .nC(w5975), .C(w5919), .Q(w5936) );
	vdp_slatch g6050 (.D(S[1]), .nC(w5976), .C(w5918), .Q(w5935) );
	vdp_aoi22 g6051 (.Z(w5934), .B2(w5980), .B1(w5936), .A1(w5935), .A2(w5916) );
	vdp_slatch g6052 (.D(S[0]), .nC(w5975), .C(w5919), .Q(w5939) );
	vdp_slatch g6053 (.D(S[0]), .nC(w5976), .C(w5918), .Q(w5938) );
	vdp_aoi22 g6054 (.Z(w5937), .B2(w5980), .B1(w5939), .A1(w5938), .A2(w5916) );
	vdp_slatch g6055 (.D(w5934), .nC(w5974), .C(w5915), .nQ(w5777) );
	vdp_slatch g6056 (.D(S[2]), .nC(w5975), .C(w5919), .Q(w5933) );
	vdp_slatch g6057 (.D(S[2]), .nC(w5976), .C(w5918), .Q(w5932) );
	vdp_aoi22 g6058 (.Z(w6016), .B2(w5980), .B1(w5933), .A1(w5932), .A2(w5916) );
	vdp_slatch g6059 (.D(w6016), .nC(w5974), .C(w5915), .nQ(w5803) );
	vdp_slatch g6060 (.D(S[3]), .nC(w5975), .C(w5919), .Q(w5931) );
	vdp_slatch g6061 (.D(S[3]), .nC(w5976), .C(w5918), .Q(w5930) );
	vdp_aoi22 g6062 (.Z(w5929), .B2(w5980), .B1(w5931), .A1(w5930), .A2(w5916) );
	vdp_slatch g6063 (.D(w5929), .nC(w5974), .C(w5915), .nQ(w5783) );
	vdp_slatch g6064 (.D(S[4]), .nC(w5975), .C(w5919), .Q(w5928) );
	vdp_slatch g6065 (.D(S[4]), .nC(w5976), .C(w5918), .Q(w5927) );
	vdp_aoi22 g6066 (.Z(w5926), .B2(w5980), .B1(w5928), .A1(w5927), .A2(w5916) );
	vdp_slatch g6067 (.D(w5926), .nC(w5974), .C(w5915), .nQ(w5786) );
	vdp_slatch g6068 (.D(S[5]), .nC(w5975), .C(w5919), .Q(w5925) );
	vdp_slatch g6069 (.D(S[5]), .nC(w5976), .C(w5918), .Q(w5924) );
	vdp_aoi22 g6070 (.Z(w5923), .B2(w5980), .B1(w5925), .A1(w5924), .A2(w5916) );
	vdp_slatch g6071 (.D(w5923), .nC(w5974), .C(w5915), .nQ(w5789) );
	vdp_slatch g6072 (.D(S[6]), .nC(w5975), .C(w5919), .Q(w5922) );
	vdp_slatch g6073 (.D(S[6]), .nC(w5976), .C(w5918), .Q(w5920) );
	vdp_aoi22 g6074 (.Z(w5921), .B2(w5980), .B1(w5922), .A1(w5920), .A2(w5916) );
	vdp_slatch g6075 (.D(w5921), .nC(w5974), .C(w5915), .nQ(w5793) );
	vdp_slatch g6076 (.D(S[7]), .nC(w5975), .C(w5919), .Q(w5917) );
	vdp_slatch g6077 (.D(S[7]), .nC(w5976), .C(w5918), .Q(w5913) );
	vdp_aoi22 g6078 (.Z(w5914), .B2(w5980), .B1(w5917), .A1(w5913), .A2(w5916) );
	vdp_slatch g6079 (.D(w5914), .nC(w5974), .C(w5915), .nQ(w5796) );
	vdp_comp_str g6080 (.nZ(w5974), .A(w5443), .Z(w5915) );
	vdp_comp_str g6081 (.nZ(w5975), .A(w4805), .Z(w5919) );
	vdp_comp_str g6082 (.nZ(w5976), .A(w4809), .Z(w5918) );
	vdp_comp_we g6083 (.nZ(w5980), .A(w5973), .Z(w5916) );
	vdp_sr_bit g6084 (.Q(w5971), .D(w5967), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6085 (.Z(w5967), .B(w5972), .A(w5940) );
	vdp_fa g6086 (.SUM(w5972), .CI(w5942), .A(w5971), .B(1'b0) );
	vdp_sr_bit g6087 (.Q(w6006), .D(w5962), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6088 (.Z(w5962), .B(w5968), .A(w5940) );
	vdp_fa g6089 (.SUM(w5968), .CO(w5942), .CI(w5943), .A(w6006), .B(1'b0) );
	vdp_sr_bit g6090 (.Q(w5963), .D(w5986), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6091 (.Z(w5986), .B(w5964), .A(w5940) );
	vdp_fa g6092 (.SUM(w5964), .CO(w5943), .CI(w5945), .A(w5963), .B(w5944) );
	vdp_sr_bit g6093 (.Q(w5959), .D(w5958), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6094 (.Z(w5958), .B(w5960), .A(w5940) );
	vdp_fa g6095 (.SUM(w5960), .CO(w5945), .CI(w5947), .A(w5959), .B(w5946) );
	vdp_sr_bit g6096 (.Q(w5950), .D(w6418), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6097 (.Q(w6418), .D(w21), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6098 (.nQ(w5948), .D(w5950), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g6099 (.nQ(w5940), .D(w5949), .nC(nHCLK1), .C(HCLK1) );
	vdp_and g6100 (.Z(w5944), .B(w5947), .A(w5955) );
	vdp_and g6101 (.Z(w5946), .B(w5947), .A(w5954) );
	vdp_and g6102 (.Z(w4448), .B(w6418), .A(w6030) );
	vdp_or g6103 (.Z(w5949), .B(w5952), .A(w6017) );
	vdp_not g6104 (.nZ(w5951), .A(M5) );
	vdp_not g6105 (.nZ(w5947), .A(w5948) );
	vdp_fa g6106 (.SUM(w5991), .CO(w5994), .CI(w5992), .A(w6044), .B(w5965) );
	vdp_aoi22 g6107 (.Z(w6055), .B2(w5977), .B1(w5993), .A1(w5991), .A2(w6040) );
	vdp_notif0 g6108 (.A(w6055), .nZ(VRAMA[9]), .nE(w6033) );
	vdp_fa g6109 (.SUM(w5982), .CO(w5992), .CI(w5988), .A(w6043), .B(w5969) );
	vdp_aoi22 g6110 (.Z(w5990), .B2(w5977), .B1(w5991), .A1(w5982), .A2(w6040) );
	vdp_notif0 g6111 (.A(w5990), .nZ(VRAMA[8]), .nE(w6033) );
	vdp_fa g6112 (.SUM(w5978), .CO(w5988), .CI(w5981), .A(w6042), .B(w5961) );
	vdp_aoi22 g6113 (.Z(w5989), .B2(w5977), .B1(w5982), .A1(w5978), .A2(w6040) );
	vdp_notif0 g6114 (.A(w5989), .nZ(VRAMA[7]), .nE(w6033) );
	vdp_fa g6115 (.SUM(w5984), .CO(w5981), .CI(1'b0), .A(w6041), .B(w5957) );
	vdp_aoi22 g6116 (.Z(w5979), .B2(w5977), .B1(w5978), .A1(w5984), .A2(w6040) );
	vdp_notif0 g6117 (.A(w5979), .nZ(VRAMA[6]), .nE(w6033) );
	vdp_not g6118 (.nZ(w6033), .A(w6047) );
	vdp_ha g6119 (.SUM(w5993), .B(w6045), .A(w5994), .CO(w5995) );
	vdp_aoi22 g6120 (.Z(w5997), .B2(w5977), .B1(w5996), .A1(w5993), .A2(w6040) );
	vdp_notif0 g6121 (.A(w5997), .nZ(VRAMA[10]), .nE(w6050) );
	vdp_ha g6122 (.SUM(w5996), .B(w6046), .A(w5995), .CO(w5998) );
	vdp_aoi22 g6123 (.Z(w5999), .B2(w5977), .B1(w6007), .A1(w5996), .A2(w6040) );
	vdp_notif0 g6124 (.A(w5999), .nZ(VRAMA[11]), .nE(w6050) );
	vdp_ha g6125 (.SUM(w6007), .B(w6049), .A(w5998), .CO(w6000) );
	vdp_aoi22 g6126 (.Z(w6002), .B2(w5977), .B1(w6001), .A1(w6007), .A2(w6040) );
	vdp_notif0 g6127 (.A(w6002), .nZ(VRAMA[12]), .nE(w6050) );
	vdp_ha g6128 (.SUM(w6001), .B(w6048), .A(w6000), .CO(w6004) );
	vdp_aoi22 g6129 (.Z(w6005), .B2(w5977), .B1(w6003), .A1(w6001), .A2(w6040) );
	vdp_notif0 g6130 (.A(w6005), .nZ(VRAMA[13]), .nE(w6050) );
	vdp_ha g6131 (.SUM(w6003), .B(w6052), .A(w6004), .CO(w6010) );
	vdp_aoi22 g6132 (.Z(w6008), .B2(w5977), .B1(w6009), .A1(w6003), .A2(w6040) );
	vdp_notif0 g6133 (.A(w6008), .nZ(VRAMA[14]), .nE(w6050) );
	vdp_ha g6134 (.SUM(w6009), .B(w6051), .A(w6010), .CO(w6011) );
	vdp_aoi22 g6135 (.Z(w6014), .B2(w5977), .B1(w6015), .A1(w6009), .A2(w6040) );
	vdp_notif0 g6136 (.A(w6014), .nZ(VRAMA[15]), .nE(w6050) );
	vdp_ha g6137 (.SUM(w6015), .B(w6054), .A(w6011) );
	vdp_aoi22 g6138 (.Z(w6013), .B2(w5977), .B1(w5071), .A1(w6015), .A2(w6040) );
	vdp_notif0 g6139 (.A(w6013), .nZ(VRAMA[16]), .nE(w6050) );
	vdp_not g6140 (.nZ(w6050), .A(w6047) );
	vdp_sr_bit g6141 (.Q(w6047), .D(w6199), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6142 (.nQ(w4371), .D(w6012), .nC(nHCLK2), .C(HCLK2) );
	vdp_and g6143 (.Z(w6199), .B(M5), .A(w21) );
	vdp_or9 g6144 (.Z(w6012), .B(w5911), .A(w5910), .C(w5830), .D(w5841), .F(w5867), .E(w5854), .G(w5880), .H(w5879), .I(w5878) );
	vdp_sr_bit g6145 (.Q(w4442), .D(w6298), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_sr_bit g6146 (.D(w6419), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_fa g6147 (.SUM(w5957), .CO(w6405), .CI(1'b0), .A(w6028), .B(w5958) );
	vdp_fa g6148 (.SUM(w5961), .CO(w6406), .CI(w6405), .A(w6029), .B(w5986) );
	vdp_fa g6149 (.SUM(w5969), .CO(w6407), .CI(w6406), .A(1'b0), .B(w5962) );
	vdp_fa g6150 (.SUM(w5965), .CI(w6407), .A(1'b0), .B(w5967) );
	vdp_notif0 g6151 (.A(1'b1), .nZ(VRAMA[0]), .nE(w6033) );
	vdp_notif0 g6152 (.A(1'b1), .nZ(VRAMA[1]), .nE(w6033) );
	vdp_not g6153 (.nZ(w5966), .A(w6034) );
	vdp_notif0 g6154 (.A(w5966), .nZ(VRAMA[2]), .nE(w6033) );
	vdp_not g6155 (.nZ(w5970), .A(w6036) );
	vdp_notif0 g6156 (.A(w5970), .nZ(VRAMA[3]), .nE(w6033) );
	vdp_not g6157 (.nZ(w5983), .A(w6035) );
	vdp_notif0 g6158 (.A(w5983), .nZ(VRAMA[4]), .nE(w6033) );
	vdp_notif0 g6159 (.A(w5985), .nZ(VRAMA[5]), .nE(w6033) );
	vdp_aoi22 g6160 (.Z(w5985), .B2(w5977), .B1(w5984), .A1(w6026), .A2(w6040) );
	vdp_comp_we g6161 (.nZ(w5977), .A(w1), .Z(w6040) );
	vdp_aon22 g6162 (.Z(w6028), .B2(w5953), .B1(w6026), .A1(w6024), .A2(w6027) );
	vdp_aon22 g6163 (.Z(w6029), .B2(w5953), .B1(w6024), .A1(w6023), .A2(w6027) );
	vdp_comp_we g6164 (.nZ(w5953), .A(w1), .Z(w6027) );
	vdp_or g6165 (.Z(w6419), .B(w6017), .A(w4448) );
	vdp_nor g6166 (.Z(w6298), .B(w5952), .A(w5951) );
	vdp_comp_str g6167 (.nZ(w6081), .A(w6037), .Z(w6053) );
	vdp_slatch g6168 (.D(w6084), .nC(w6081), .C(w6053), .Q(w5910) );
	vdp_aon22 g6169 (.Z(w6085), .B2(w6056), .B1(w5938), .A1(DB[0]), .A2(w6038) );
	vdp_slatch g6170 (.D(w6086), .nC(w6081), .C(w6053), .Q(w5911) );
	vdp_aon22 g6171 (.Z(w6087), .B2(w6056), .B1(w5935), .A1(DB[1]), .A2(w6038) );
	vdp_slatch g6172 (.D(w6088), .nC(w6081), .C(w6053), .Q(w5830) );
	vdp_aon22 g6173 (.Z(w6089), .B2(w6056), .B1(w5932), .A1(DB[2]), .A2(w6038) );
	vdp_slatch g6174 (.D(w6090), .nC(w6081), .C(w6053), .Q(w5841) );
	vdp_aon22 g6175 (.Z(w6091), .B2(w6056), .B1(w5930), .A1(DB[3]), .A2(w6038) );
	vdp_slatch g6176 (.D(w6092), .nC(w6081), .C(w6053), .Q(w5854) );
	vdp_aon22 g6177 (.Z(w6093), .B2(w6056), .B1(w5927), .A1(DB[4]), .A2(w6038) );
	vdp_slatch g6178 (.D(w6094), .nC(w6081), .C(w6053), .Q(w5867) );
	vdp_aon22 g6179 (.Z(w6095), .B2(w6056), .B1(w5924), .A1(w6069), .A2(w6038) );
	vdp_slatch g6180 (.D(w6096), .nC(w6081), .C(w6053), .Q(w5880) );
	vdp_aon22 g6181 (.Z(w6097), .B2(w6056), .B1(w5920), .A1(w6074), .A2(w6038) );
	vdp_slatch g6182 (.D(w6099), .nC(w6081), .C(w6053), .Q(w5879) );
	vdp_aon22 g6183 (.Z(w6100), .B2(w6056), .B1(w5913), .A1(DB[7]), .A2(w6038) );
	vdp_slatch g6184 (.D(w6098), .nC(w6081), .C(w6053), .Q(w5878) );
	vdp_aon22 g6185 (.Z(w6101), .B2(w6056), .B1(w4918), .A1(DB[8]), .A2(w6038) );
	vdp_slatch g6186 (.D(w6071), .nC(w6067), .C(w6039), .Q(w6043) );
	vdp_aon22 g6187 (.Z(w6108), .B2(w6056), .B1(w5933), .A1(DB[2]), .A2(w6038) );
	vdp_slatch g6188 (.D(w6070), .nC(w6067), .C(w6039), .Q(w6044) );
	vdp_aon22 g6189 (.Z(w6103), .B2(w6056), .B1(w5931), .A1(DB[3]), .A2(w6038) );
	vdp_slatch g6190 (.D(w6078), .nC(w6067), .C(w6039), .Q(w6045) );
	vdp_aon22 g6191 (.Z(w6104), .B2(w6056), .B1(w5928), .A1(DB[4]), .A2(w6038) );
	vdp_slatch g6192 (.D(w6077), .nC(w6067), .C(w6039), .Q(w6046) );
	vdp_aon22 g6193 (.Z(w6107), .B2(w6056), .B1(w5925), .A1(w6069), .A2(w6038) );
	vdp_slatch g6194 (.D(w6075), .nC(w6067), .C(w6039), .Q(w6049) );
	vdp_aon22 g6195 (.Z(w6109), .B2(w6056), .B1(w5922), .A1(w6074), .A2(w6038) );
	vdp_slatch g6196 (.D(w6076), .nC(w6067), .C(w6039), .Q(w6048) );
	vdp_aon22 g6197 (.Z(w6110), .B2(w6056), .B1(w5917), .A1(DB[7]), .A2(w6038) );
	vdp_slatch g6198 (.D(w6073), .nC(w6067), .C(w6039), .Q(w6052) );
	vdp_aon22 g6199 (.Z(w6111), .B2(w6056), .B1(w4859), .A1(DB[8]), .A2(w6038) );
	vdp_slatch g6200 (.D(w6065), .nC(w6067), .C(w6039), .Q(w6051) );
	vdp_aon22 g6201 (.Z(w6064), .B2(w6056), .B1(w4919), .A1(DB[9]), .A2(w6038) );
	vdp_slatch g6202 (.D(w6082), .nC(w6067), .C(w6039), .Q(w6054) );
	vdp_aon22 g6203 (.Z(w6083), .B2(w6056), .B1(w4926), .A1(DB[10]), .A2(w6038) );
	vdp_slatch g6204 (.D(w6068), .nC(w6067), .C(w6039), .Q(w6041) );
	vdp_aon22 g6205 (.Z(w6105), .B2(w6056), .B1(w5939), .A1(DB[0]), .A2(w6038) );
	vdp_slatch g6206 (.D(w6112), .nC(w6067), .C(w6039), .Q(w6042) );
	vdp_aon22 g6207 (.Z(w6106), .B2(w6056), .B1(w5936), .A1(DB[1]), .A2(w6038) );
	vdp_comp_str g6208 (.nZ(w6067), .A(w6037), .Z(w6039) );
	vdp_not g6209 (.nZ(w6037), .A(w6194) );
	vdp_oai21 g6210 (.Z(w6194), .B(HCLK1), .A1(w5952), .A2(w112) );
	vdp_sr_bit g6211 (.Q(w6195), .D(w6197), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6212 (.Q(w5443), .D(w6196), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6213 (.Q(w5973), .D(w6198), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6214 (.Q(w6102), .D(w5404), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g6215 (.Q(w6020), .D(w6025), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w6017), .CI(w21), .L(w6022), .nL(w6059), .CO(w6060) );
	vdp_cnt_bit_load g6216 (.Q(w6058), .D(w6021), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w6017), .CI(w6060), .L(w6022), .nL(w6059) );
	vdp_comp_we g6217 (.nZ(w6059), .A(w5952), .Z(w6022) );
	vdp_not g6218 (.nZ(w6025), .A(w6061) );
	vdp_not g6219 (.nZ(w6021), .A(w6057) );
	vdp_not g6220 (.nZ(w6018), .A(w107) );
	vdp_nand g6221 (.Z(w6113), .B(w107), .A(w4442) );
	vdp_nand g6222 (.Z(w6019), .B(w6018), .A(w4442) );
	vdp_not g6223 (.nZ(w6056), .A(w6019) );
	vdp_nor g6224 (.Z(w6030), .B(w6058), .A(w6020) );
	vdp_and g6225 (.Z(w5952), .B(w6030), .A(w21) );
	vdp_rs_ff g6226 (.Q(w6197), .R(w6031), .S(w6017) );
	vdp_and3 g6227 (.Z(w6196), .B(w5404), .A(w4449), .C(w6195) );
	vdp_cnt_bit g6228 (.Q(w6198), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w38), .CI(w6102) );
	vdp_not g6229 (.nZ(w6038), .A(w6113) );
	vdp_not g6230 (.nZ(w6063), .A(w4406) );
	vdp_not g6231 (.nZ(w6066), .A(w4407) );
	vdp_comp_str g6232 (.nZ(w6062), .A(w6037), .Z(w6115) );
	vdp_not g6233 (.nZ(w6123), .A(w112) );
	vdp_aon22 g6234 (.Z(w6125), .B2(w6056), .B1(w4977), .A1(DB[0]), .A2(w6038) );
	vdp_slatch g6235 (.D(w6114), .nC(w6062), .C(w6115), .Q(w5905) );
	vdp_bufif0 g6236 (.A(w6122), .Z(DB[0]), .nE(w6123) );
	vdp_aon222 g6237 (.Z(w6122), .B2(w4408), .B1(w5910), .A1(w5905), .A2(w6063), .C1(w6041), .C2(w6066) );
	vdp_aon22 g6238 (.Z(w6128), .B2(w6056), .B1(w5053), .A1(DB[1]), .A2(w6038) );
	vdp_slatch g6239 (.D(w6124), .nC(w6062), .C(w6115), .Q(w5906) );
	vdp_bufif0 g6240 (.A(w6126), .Z(DB[1]), .nE(w6123) );
	vdp_aon222 g6241 (.Z(w6126), .B2(w4408), .B1(w5911), .A1(w5906), .A2(w6063), .C1(w6042), .C2(w6066) );
	vdp_aon22 g6242 (.Z(w6130), .B2(w6056), .B1(w5072), .A1(DB[2]), .A2(w6038) );
	vdp_slatch g6243 (.D(w6127), .nC(w6062), .C(w6115), .Q(w5907) );
	vdp_bufif0 g6244 (.A(w6129), .Z(DB[2]), .nE(w6123) );
	vdp_aon222 g6245 (.Z(w6129), .B2(w4408), .B1(w5830), .A1(w5907), .A2(w6063), .C1(w6043), .C2(w6066) );
	vdp_aon22 g6246 (.Z(w6139), .B2(w6056), .B1(w5039), .A1(DB[3]), .A2(w6038) );
	vdp_slatch g6247 (.D(w6131), .nC(w6062), .C(w6115), .Q(w5912) );
	vdp_bufif0 g6248 (.A(w6138), .Z(DB[3]), .nE(w6123) );
	vdp_aon222 g6249 (.Z(w6138), .B2(w4408), .B1(w5841), .A1(w5912), .A2(w6063), .C1(w6044), .C2(w6066) );
	vdp_aon22 g6250 (.Z(w6136), .B2(w6056), .B1(w4387), .A1(DB[4]), .A2(w6038) );
	vdp_slatch g6251 (.D(w6061), .nC(w6062), .C(w6115), .Q(w5908) );
	vdp_bufif0 g6252 (.A(w6137), .Z(DB[4]), .nE(w6123) );
	vdp_aon222 g6253 (.Z(w6137), .B2(w4408), .B1(w5854), .A1(w5908), .A2(w6063), .C1(w6045), .C2(w6066) );
	vdp_aon22 g6254 (.Z(w6134), .B2(w6056), .B1(w4432), .A1(w6069), .A2(w6038) );
	vdp_slatch g6255 (.D(w6057), .nC(w6062), .C(w6115), .Q(w5909) );
	vdp_bufif0 g6256 (.A(w6135), .Z(w6069), .nE(w6123) );
	vdp_aon222 g6257 (.Z(w6135), .B2(w4408), .B1(w5867), .A1(w5909), .A2(w6063), .C1(w6046), .C2(w6066) );
	vdp_aon22 g6258 (.Z(w6132), .B2(w6056), .B1(w4388), .A1(w6074), .A2(w6038) );
	vdp_slatch g6259 (.D(w6133), .nC(w6062), .C(w6115), .Q(w5954) );
	vdp_bufif0 g6260 (.A(w6155), .Z(w6074), .nE(w6123) );
	vdp_aon222 g6261 (.Z(w6155), .B2(w4408), .B1(w5880), .A1(w5954), .A2(w6063), .C1(w6049), .C2(w6066) );
	vdp_aon22 g6262 (.Z(w6151), .B2(w6056), .B1(w4384), .A1(DB[7]), .A2(w6038) );
	vdp_slatch g6263 (.D(w6152), .nC(w6072), .C(w6153), .Q(w5955) );
	vdp_bufif0 g6264 (.A(w6154), .Z(DB[7]), .nE(w6123) );
	vdp_aon222 g6265 (.Z(w6154), .B2(w4408), .B1(w5879), .A1(w5955), .A2(w6063), .C1(w6048), .C2(w6066) );
	vdp_aon22 g6266 (.Z(w6149), .B2(w6056), .B1(w6116), .A1(DB[8]), .A2(w6038) );
	vdp_slatch g6267 (.D(w6150), .nC(w6072), .C(w6153), .Q(w6034) );
	vdp_bufif0 g6268 (.A(w6420), .Z(DB[8]), .nE(w6123) );
	vdp_aon222 g6269 (.Z(w6420), .B2(w4408), .B1(w5878), .A1(w6034), .A2(w6063), .C1(w6052), .C2(w6066) );
	vdp_aon22 g6270 (.Z(w6147), .B2(w6056), .B1(w6121), .A1(DB[9]), .A2(w6038) );
	vdp_slatch g6271 (.D(w6148), .nC(w6072), .C(w6153), .Q(w6036) );
	vdp_bufif0 g6272 (.A(w6156), .Z(DB[9]), .nE(w6123) );
	vdp_aon222 g6273 (.Z(w6156), .B2(w4408), .B1(1'b0), .A1(w6036), .A2(w6063), .C1(w6051), .C2(w6066) );
	vdp_aon22 g6274 (.Z(w6145), .B2(w6056), .B1(w6120), .A1(DB[10]), .A2(w6038) );
	vdp_slatch g6275 (.D(w6146), .nC(w6072), .C(w6153), .Q(w6035) );
	vdp_bufif0 g6276 (.A(w6157), .Z(DB[10]), .nE(w6123) );
	vdp_aon222 g6277 (.Z(w6157), .B2(w4408), .B1(1'b0), .A1(w6035), .A2(w6063), .C1(w6054), .C2(w6066) );
	vdp_aon22 g6278 (.Z(w6143), .B2(w6056), .B1(w6119), .A1(DB[11]), .A2(w6038) );
	vdp_slatch g6279 (.D(w6144), .nC(w6072), .C(w6153), .Q(w6026) );
	vdp_bufif0 g6280 (.A(w6026), .Z(DB[11]), .nE(w6123) );
	vdp_aon22 g6281 (.Z(w6142), .B2(w6056), .B1(w6118), .A1(DB[12]), .A2(w6038) );
	vdp_slatch g6282 (.D(w6158), .nC(w6072), .C(w6153), .Q(w6024) );
	vdp_bufif0 g6283 (.A(w6024), .Z(DB[12]), .nE(w6123) );
	vdp_aon22 g6284 (.Z(w6140), .B2(w6056), .B1(w6117), .A1(DB[13]), .A2(w6038) );
	vdp_slatch g6285 (.D(w6141), .nC(w6072), .C(w6153), .Q(w6023) );
	vdp_bufif0 g6286 (.A(w6023), .Z(DB[13]), .nE(w6123) );
	vdp_comp_str g6287 (.nZ(w6072), .A(w6037), .Z(w6153) );
	vdp_sr_bit g6288 (.Q(w4544), .D(w119), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6289 (.Q(w4548), .D(VRAMA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6290 (.Q(w6166), .D(w6159), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6291 (.Q(w4537), .D(VRAMA[3]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6292 (.Q(w4539), .D(VRAMA[4]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6293 (.Q(w4540), .D(VRAMA[5]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6294 (.Q(w4541), .D(VRAMA[6]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6295 (.Q(w4542), .D(VRAMA[7]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6296 (.Q(w4543), .D(VRAMA[8]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6297 (.Q(w4484), .D(w6163), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6298 (.Q(w4483), .D(w6164), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_and g6299 (.Z(w6163), .B(w122), .A(w6165) );
	vdp_and g6300 (.Z(w6164), .B(w121), .A(w6165) );
	vdp_sr_bit g6301 (.Q(w6179), .D(RD_DATA[0]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6302 (.Q(w6180), .D(RD_DATA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6303 (.Q(w6182), .D(w321), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6304 (.Q(w6181), .D(RD_DATA[2]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_V_PLA g6305 (.o0(w1812), .o1(w1813), .o2(w1814), .o3(w1815), .o4(w1816), .o5(w1817), .o6(w1818), .o7(w1819), .o8(w1820), .o9(w1821), .o10(w1822), .o11(w6619), .o12(w6620), .o13(w6618), .o14(w1823), .o15(w6539), .o16(w6540), .o17(w6541), .o18(w1824), .o19(w1825), .o20(w1826), .o21(w1827), .o22(w6542), .o23(w1828), .o24(w1904), .o25(w1829), .o26(w1830), .o27(w1905), .o28(w1919), .o29(w1918), .o30(w1939), .o31(w1846), .o32(w1811), .o33(w1810), .o34(w1847), .o35(w1831), .o36(w1848), .o37(w1849), .o38(w1809), .o39(w1808), .o40(w1852), .o41(w1850), .o42(w1851), .o43(w1807), .o44(w1806), .o45(w1805), .o46(w1804), .o47(w6427), .Vcnt0(w1641), .Vcnt1(w1781), .Vcnt2(w1860), .Vcnt3(w1766), .Vcnt4(w1859), .Vcnt5(w1720), .Vcnt6(w1685), .Vcnt7(w1755), .Vcnt8(w1782), .ODD_EVEN(ODD_EVEN), .LS0(LSM0), .PAL(PAL), .nPAL(w1774), .i2(w1773), .i3(w1762), .M5(M5) );
	vdp_not g6306 (.A(w576), .nZ(w6425) );
	vdp_not g6307 (.A(w933), .nZ(w6426) );
	vdp_not g6308 (.nZ(w2368), .A(w6425) );
	vdp_not g6309 (.nZ(w2369), .A(w6426) );
	vdp_cram g6310 (.q8(w2655), .D8(w2660), .q7(w2757), .D7(w2656), .q6(w2654), .D6(w2657), .q5(w2659), .D5(w2658), .q4(w2653), .D4(w2661), .q3(w2662), .D3(w2879), .q2(w2652), .D2(w2663), .q1(w2651), .D1(w2664), .q0(w2649), .D0(w2665), .A0(w2684), .A1(w2688), .CLK(HCLK1), .A2(w2694), .A3(w2704), .A4(w2725), .A5(w2724), .Bi(w2731), .Ai(w2730) );
	vdp_linebuf_ram g6311 (.q0(w5175), .D0(w5525), .q1(w5155), .D1(w5524), .q2(w5117), .D2(w5523), .q3(w5194), .D3(w5538), .q4(w5546), .D4(w5539), .q5(w5553), .D5(w5540), .q6(w5512), .D6(w5541), .q7(w5174), .D7(w5522), .q8(w5158), .D8(w5521), .q9(w5138), .D9(w5520), .q10(w5511), .D10(w5502), .q11(w5513), .D11(w5501), .q12(w5514), .D12(w5534), .q13(w5517), .D13(w5535), .q14(w5173), .D14(w5525), .q15(w5156), .D15(w5524), .q16(w5140), .D16(w5523), .q17(w5186), .D17(w5526), .q18(w5515), .D18(w5533), .q19(w5516), .D19(w5527), .q20(w5529), .D20(w5528), .q21(w5172), .D21(w5522), .q22(w5162), .D22(w5521), .q23(w5135), .D23(w5520), .q24(w5187), .D24(w5508), .q25(w5505), .D25(w5506), .q26(w5510), .D26(w5519), .q27(w5532), .D27(w5518), .CLK(w4369), .A5(w4363), .A4(w4364), .A3(w4365), .A2(w4366), .A1(w4367), .A0(w4368), .Ai(w5531), .Bi(w5500), .Ci(w5499), .Di(w5498) );
	vdp_linebuf_ram g6312 (.q0(w5181), .D0(w5525), .q1(w5152), .D1(w5524), .q2(w5143), .D2(w5523), .q3(w5124), .D3(w5170), .q4(w5123), .D4(w5168), .q5(w5122), .D5(w5169), .q6(w5507), .D6(w6161), .q7(w5176), .D7(w5522), .q8(w5154), .D8(w5521), .q9(w5141), .D9(w5520), .q10(w5191), .D10(w5164), .q11(w5120), .D11(w5165), .q12(w5121), .D12(w5166), .q13(w5504), .D13(w5159), .q14(w5177), .D14(w5525), .q15(w5153), .D15(w5524), .q16(w5144), .D16(w5523), .q17(w5198), .D17(w5133), .q18(w5118), .D18(w5116), .q19(w5119), .D19(w5131), .q20(w5503), .D20(w5132), .q21(w5126), .D21(w5522), .q22(w5125), .D22(w5521), .q23(w5139), .D23(w5520), .q24(w5192), .D24(w6162), .q25(w5536), .D25(w5127), .q26(w5537), .D26(w5128), .q27(w5509), .D27(w5129), .A0(w4368), .CLK(w4369), .A5(w4363), .A3(w4365), .A4(w4364), .A2(w4366), .A1(w4367), .Ai(w5240), .Bi(w5224), .Ci(w5236), .Di(w5226) );
	vdp_att_cashe_ram2 g6313 (.q0(w4561), .D0(FIFOo[0]), .q1(w4560), .D1(FIFOo[1]), .q2(w4559), .D2(FIFOo[2]), .q3(w4558), .D3(FIFOo[3]), .q4(w4534), .D4(FIFOo[4]), .q5(w4533), .D5(FIFOo[5]), .q6(w4528), .D6(FIFOo[6]), .q7(w4704), .D7(w6179), .q8(w4743), .D8(w6180), .q9(w4727), .D9(w6181), .q10(w4724), .D10(w6182), .CLK(HCLK1), .A6(w6186), .A5(w6187), .A1(w6192), .A0(w6191), .A4(w6188), .A3(w6189), .A2(w6190), .Ai(w6183), .Bi(w4546) );
	vdp_att_cashe_ram1 g6314 (.q0(w4593), .D0(FIFOo[0]), .q1(w4596), .D1(FIFOo[1]), .q2(w4589), .D2(FIFOo[2]), .q3(w4590), .D3(FIFOo[3]), .q4(w4572), .D4(FIFOo[4]), .q5(w4564), .D5(FIFOo[5]), .q6(w4565), .D6(FIFOo[6]), .q7(w4563), .D7(FIFOo[7]), .q8(w4562), .D8(w6179), .q9(w4557), .D9(w6180), .CLK(HCLK1), .A0(w6191), .A1(w6192), .A2(w6190), .A3(w6189), .A4(w6188), .A5(w6187), .A6(w6186), .Ai(w6185), .Bi(w6184) );
	vdp_att_temp_ram g6315 (.A4(w4466), .A0(w4470), .A1(w4469), .A2(w4468), .A3(w4467), .q0(w6068), .D0(w6105), .q1(w6112), .D1(w6106), .q2(w6071), .D2(w6108), .q3(w6070), .D3(w6103), .q4(w6078), .D4(w6104), .q5(w6077), .D5(w6107), .q6(w6075), .D6(w6109), .q7(w6076), .D7(w6110), .q8(w6073), .D8(w6111), .q9(w6065), .D9(w6064), .q10(w6082), .D10(w6083), .q11(w6084), .D11(w6085), .q12(w6086), .D12(w6087), .q13(w6088), .D13(w6089), .q14(w6090), .D14(w6091), .q15(w6092), .D15(w6093), .q16(w6094), .D16(w6095), .q17(w6096), .D17(w6097), .q18(w6099), .D18(w6100), .q19(w6098), .D19(w6101), .q20(w6114), .D20(w6125), .q21(w6124), .D21(w6128), .q22(w6127), .D22(w6130), .q23(w6131), .D23(w6139), .q24(w6061), .D24(w6136), .q25(w6057), .D25(w6134), .q26(w6133), .D26(w6132), .q26(w6152), .D26(w6151), .q27(w6150), .D27(w6149), .q28(w6148), .D28(w6147), .q29(w6146), .D29(w6145), .q30(w6144), .D30(w6143), .q31(w6158), .D[31](w6142), .q32(w6141), .D32(w6140), .CLK(HCLK1), .Ai(w4433), .Bi(w4434), .Ci(w4438) );
	vdp_vsram g6316 (.CLK(HCLK1), .D10(w3870), .q10(w3832), .D9(w3874), .q9(w3825), .D8(w3872), .q8(w3847), .D7(w3871), .q7(w3817), .D6(w3859), .q6(w3813), .D5(w3857), .q5(w3805), .D4(w3864), .q4(w3801), .D3(w3866), .q3(w3798), .D2(w3869), .q2(w3852), .D1(w3831), .q1(w3793), .D0(w3845), .q0(w3788), .A1(w3611), .A2(w3583), .A3(w3582), .A4(w3581), .A5(w3580), .A0(w3612), .Ai(w3579), .Bi(w3578) );
	vdp_not g6317 (.nZ(w1756), .A(w6427) );
	vdp_not g6318 (.nZ(PAL), .A(w6428) );
	vdp_H_PLA g6319 (.HPLA0(HPLA0), .HPLA1(HPLA1), .HPLA2(HPLA2), .HPLA3(HPLA3), .HPLA4(HPLA4), .HPLA5(HPLA5), .HPLA7(HPLA7), .HPLA8(HPLA8), .HPLA9(HPLA9), .HPLA6(HPLA6), .HPLA10(HPLA10), .HPLA11(HPLA11), .HPLA16(HPLA16), .HPLA15(HPLA15), .HPLA14(HPLA14), .HPLA13(HPLA13), .HPLA12(HPLA12), .i0(w59), .HPLA17(HPLA17), .HPLA18(HPLA18), .HPLA19(HPLA19), .HPLA20(HPLA20), .HPLA21(HPLA21), .HPLA22(HPLA22), .Hcnt0(w1863), .Hcnt1(w1625), .Hcnt2(w1630), .Hcnt3(w1629), .Hcnt4(w1674), .Hcnt5(w1706), .Hcnt6(w1838), .Hcnt7(w1683), .Hcnt8(w1876), .H40(H40), .M5(M5), .B(w1865), .C(w1609), .A(w1679), .HPLA[23](HPLA23), .HPLA[24](HPLA24), .HPLA[25](HPLA25), .HPLA[26](HPLA26), .HPLA[27](HPLA27), .HPLA[28](HPLA28), .HPLA[29](HPLA29), .HPLA[30](HPLA30), .HPLA[31](HPLA31), .HPLA[32](HPLA32), .HPLA[33](HPLA33), .i3(w1842), .HPLA[35](HPLA35), .HPLA[36](HPLA36), .HPLA[34](HPLA34) );
	vdp_slatch g5073 (.D(S[4]), .nC(w4864), .C(w4865), .Q(w5052) );
endmodule // VDP

// Module Definitions [It is possible to wrap here on your primitives]

module vdp_slatch (  nQ, D, C, nC);

	output wire nQ;
	input wire D;
	input wire C;
	input wire nC;

endmodule // vdp_slatch

module vdp_sr_bit (  D, C2, C1, Q, nC2, nC1);

	input wire D;
	input wire C2;
	input wire C1;
	output wire Q;
	input wire nC2;
	input wire nC1;

endmodule // vdp_sr_bit

module vdp_notif0 (  A, nZ, nE);

	input wire A;
	output wire nZ;
	input wire nE;

endmodule // vdp_notif0

module vdp_aon22 (  Z, A1, A2, B1, B2);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire B1;
	input wire B2;

endmodule // vdp_aon22

module vdp_not (  A, nZ);

	input wire A;
	output wire nZ;

endmodule // vdp_not

module vdp_comp_str (  A, Z, nZ);

	input wire A;
	output wire Z;
	output wire nZ;

endmodule // vdp_comp_str

module vdp_comp_we (  A, Z, nZ);

	input wire A;
	output wire Z;
	output wire nZ;

endmodule // vdp_comp_we

module vdp_and (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_and

module vdp_nand (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_nand

module vdp_and3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_and3

module vdp_fa (  SUM, A, B, CO, CI);

	output wire SUM;
	input wire A;
	input wire B;
	output wire CO;
	input wire CI;

endmodule // vdp_fa

module vdp_comp_dff (  D, C2, C1, Q, nC2, nC1);

	input wire D;
	input wire C2;
	input wire C1;
	output wire Q;
	input wire nC2;
	input wire nC1;

endmodule // vdp_comp_dff

module vdp_or (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_or

module vdp_xor (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_xor

module vdp_aoi21 (  Z, B, A1, A2);

	output wire Z;
	input wire B;
	input wire A1;
	input wire A2;

endmodule // vdp_aoi21

module vdp_nor (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_nor

module vdp_and5 (  Z, A, B, C, D, E);

	output wire Z;
	input wire A;
	input wire B;
	input wire C;
	input wire D;
	input wire E;

endmodule // vdp_and5

module vdp_aon2222 (  C2, B2, A2, C1, B1, A1, Z, D2, D1);

	input wire C2;
	input wire B2;
	input wire A2;
	input wire C1;
	input wire B1;
	input wire A1;
	output wire Z;
	input wire D2;
	input wire D1;

endmodule // vdp_aon2222

module vdp_cnt_bit (  R, Q, C1, C2, nC1, nC2, CI);

	input wire R;
	output wire Q;
	input wire C1;
	input wire C2;
	input wire nC1;
	input wire nC2;
	input wire CI;

endmodule // vdp_cnt_bit

module vdp_oai21 (  A1, Z, A2, B);

	input wire A1;
	output wire Z;
	input wire A2;
	input wire B;

endmodule // vdp_oai21

module vdp_comb1 (  Z, A1, B, A2, C);

	output wire Z;
	input wire A1;
	input wire B;
	input wire A2;
	input wire C;

endmodule // vdp_comb1

module vdp_rs_ff (  Q, R, S);

	output wire Q;
	input wire R;
	input wire S;

endmodule // vdp_rs_ff

module vdp_and4 (  A, Z, B, C, D);

	input wire A;
	output wire Z;
	input wire B;
	input wire C;
	input wire D;

endmodule // vdp_and4

module vdp_or3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_or3

module vdp_bufif0 (  A, Z, nE);

	input wire A;
	output wire Z;
	input wire nE;

endmodule // vdp_bufif0

module vdp_aoi221 (  Z, A2, B1, B2, A1, C);

	output wire Z;
	input wire A2;
	input wire B1;
	input wire B2;
	input wire A1;
	input wire C;

endmodule // vdp_aoi221

module vdp_aon33 (  Z, A2, B1, B2, A1, A3, B3);

	output wire Z;
	input wire A2;
	input wire B1;
	input wire B2;
	input wire A1;
	input wire A3;
	input wire B3;

endmodule // vdp_aon33

module vdp_dlatch_inv (  D, C, Q, nC);

	input wire D;
	input wire C;
	output wire Q;
	input wire nC;

endmodule // vdp_dlatch_inv

module vdp_cnt_bit_load (  D, nL, L, R, Q, C1, C2, nC1, nC2, CI, CO);

	input wire D;
	input wire nL;
	input wire L;
	input wire R;
	output wire Q;
	input wire C1;
	input wire C2;
	input wire nC1;
	input wire nC2;
	input wire CI;
	output wire CO;

endmodule // vdp_cnt_bit_load

module vdp_nand3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_nand3

module vdp_nor3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_nor3

module vdp_dff (  Q, R, C, D);

	output wire Q;
	input wire R;
	input wire C;
	input wire D;

endmodule // vdp_dff

module vdp_ha (  SUM, A, B, CO);

	output wire SUM;
	input wire A;
	input wire B;
	output wire CO;

endmodule // vdp_ha

module vdp_slatch_r (  Q, D, R, C, nC);

	output wire Q;
	input wire D;
	input wire R;
	input wire C;
	input wire nC;

endmodule // vdp_slatch_r

module vdp_or5 (  C, A, B, Z, D, E);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;
	input wire E;

endmodule // vdp_or5

module vdp_2a3oi (  A1, B, Z, A2, C);

	input wire A1;
	input wire B;
	output wire Z;
	input wire A2;
	input wire C;

endmodule // vdp_2a3oi

module vdp_nor5 (  C, A, B, Z, D, E);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;
	input wire E;

endmodule // vdp_nor5

module vdp_or4 (  C, A, B, Z, D);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;

endmodule // vdp_or4

module vdp_aoi22 (  Z, A1, A2, B1, B2);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire B1;
	input wire B2;

endmodule // vdp_aoi22

module vdp_aon222 (  C2, B2, A2, C1, B1, A1, Z);

	input wire C2;
	input wire B2;
	input wire A2;
	input wire C1;
	input wire B1;
	input wire A1;
	output wire Z;

endmodule // vdp_aon222

module vdp_dlatch (  D, C, Q, nC);

	input wire D;
	input wire C;
	output wire Q;
	input wire nC;

endmodule // vdp_dlatch

module vdp_nor4 (  C, A, B, Z, D);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;

endmodule // vdp_nor4

module vdp_and6 (  C, A, B, Z, D, E, F);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;
	input wire E;
	input wire F;

endmodule // vdp_and6

module vdp_n_fet (  Z, A);

	output wire Z;
	input wire A;

endmodule // vdp_n_fet

module vdp_2A3OI (  Z, A1, A2, C, B);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire C;
	input wire B;

endmodule // vdp_2A3OI

module vdp_tff (  C2, C1, nC2, nC1, CI, R, A, Q);

	input wire C2;
	input wire C1;
	input wire nC2;
	input wire nC1;
	input wire CI;
	input wire R;
	input wire A;
	output wire Q;

endmodule // vdp_tff

module vdp_SDELAY8 (  Q, D, nC1, C1, nC2, C2, nC3, C3, nC4, C4, nC5, C5, nC6, C6, nC7, C7, nC8, C8, nC9, C9, nC10, C10, nC11, C11, nC12, C12, nC13, C13, nC14, C14, nC15, C15, nC16, C16);

	output wire Q;
	input wire D;
	input wire nC1;
	input wire C1;
	input wire nC2;
	input wire C2;
	input wire nC3;
	input wire C3;
	input wire nC4;
	input wire C4;
	input wire nC5;
	input wire C5;
	input wire nC6;
	input wire C6;
	input wire nC7;
	input wire C7;
	input wire nC8;
	input wire C8;
	input wire nC9;
	input wire C9;
	input wire nC10;
	input wire C10;
	input wire nC11;
	input wire C11;
	input wire nC12;
	input wire C12;
	input wire nC13;
	input wire C13;
	input wire nC14;
	input wire C14;
	input wire nC15;
	input wire C15;
	input wire nC16;
	input wire C16;

endmodule // vdp_SDELAY8

module vdp_SDELAY7 (  Q, D, C1, nC1, C2, nC2, nC3, C4, nC4, C5, nC5, C6, nC6, C7, nC7, C8, nC8, C9, nC9, C10, nC10, C11, nC11, C12, nC12, C13, nC13, C14, nC14, C3);

	output wire Q;
	input wire D;
	input wire C1;
	input wire nC1;
	input wire C2;
	input wire nC2;
	input wire nC3;
	input wire C4;
	input wire nC4;
	input wire C5;
	input wire nC5;
	input wire C6;
	input wire nC6;
	input wire C7;
	input wire nC7;
	input wire C8;
	input wire nC8;
	input wire C9;
	input wire nC9;
	input wire C10;
	input wire nC10;
	input wire C11;
	input wire nC11;
	input wire C12;
	input wire nC12;
	input wire C13;
	input wire nC13;
	input wire C14;
	input wire nC14;
	input wire C3;

endmodule // vdp_SDELAY7

module vdp_or8 (  Z, A, B, C, D, E, F, G, H);

	output wire Z;
	input wire A;
	input wire B;
	input wire C;
	input wire D;
	input wire E;
	input wire F;
	input wire G;
	input wire H;

endmodule // vdp_or8

module vdp_or7 (  Z, A, B, C, D, E, F, G);

	output wire Z;
	input wire A;
	input wire B;
	input wire C;
	input wire D;
	input wire E;
	input wire F;
	input wire G;

endmodule // vdp_or7

module vdp_clkgen (  PH, CLK1, nCLK1, CLK2, nCLK2);

	input wire PH;
	output wire CLK1;
	output wire nCLK1;
	output wire CLK2;
	output wire nCLK2;

endmodule // vdp_clkgen

module vdp_cgi2a (  Z, A, C, B);

	output wire Z;
	input wire A;
	input wire C;
	input wire B;

endmodule // vdp_cgi2a

module vdp_nand4 (  Z, A, B, D, C);

	output wire Z;
	input wire A;
	input wire B;
	input wire D;
	input wire C;

endmodule // vdp_nand4

module vdp_lfsr_bit (  Q, A, C2, C1, nC2, nC1, C, B);

	output wire Q;
	input wire A;
	input wire C2;
	input wire C1;
	input wire nC2;
	input wire nC1;
	input wire C;
	input wire B;

endmodule // vdp_lfsr_bit

module vdp_aoi222 (  Z, A1, B1, B2, A2, C1, C2);

	output wire Z;
	input wire A1;
	input wire B1;
	input wire B2;
	input wire A2;
	input wire C1;
	input wire C2;

endmodule // vdp_aoi222

module vdp_aon333 (  Z, A1, A2, A3, B1, B2, B3, C1, C2, C3);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire A3;
	input wire B1;
	input wire B2;
	input wire B3;
	input wire C1;
	input wire C2;
	input wire C3;

endmodule // vdp_aon333

module vdp_aoi33 (  Z, A1, A2, A3, B1, B2, B3);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire A3;
	input wire B1;
	input wire B2;
	input wire B3;

endmodule // vdp_aoi33

module vdp_comp_strong (  nZ, Z, A);

	output wire nZ;
	output wire Z;
	input wire A;

endmodule // vdp_comp_strong

module vdp_neg_dff (  Q, C, D, R);

	output wire Q;
	input wire C;
	input wire D;
	input wire R;

endmodule // vdp_neg_dff

module vdp_aon2x8 (  Z, A1, B1, C1, D2, A2, B2, C2, D1, E2, F1, E1, F2, G1, H2, G2, H1);

	output wire Z;
	input wire A1;
	input wire B1;
	input wire C1;
	input wire D2;
	input wire A2;
	input wire B2;
	input wire C2;
	input wire D1;
	input wire E2;
	input wire F1;
	input wire E1;
	input wire F2;
	input wire G1;
	input wire H2;
	input wire G2;
	input wire H1;

endmodule // vdp_aon2x8

module vdp_xnor (  Z, A, B);

	output wire Z;
	input wire A;
	input wire B;

endmodule // vdp_xnor

module vdp_oai211 (  Z, A1, A2, B, C);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire B;
	input wire C;

endmodule // vdp_oai211

module vdp_aoi31 (  Z, B3, B2, B1, A);

	output wire Z;
	input wire B3;
	input wire B2;
	input wire B1;
	input wire A;

endmodule // vdp_aoi31

module vdp_AOI222 (  Z, B1, A1, B2, A2, C1, C2);

	output wire Z;
	input wire B1;
	input wire A1;
	input wire B2;
	input wire A2;
	input wire C1;
	input wire C2;

endmodule // vdp_AOI222

module vdp_cnt_bit_rev (  nC2, nC1, C2, C1, Q, CI, B, A);

	input wire nC2;
	input wire nC1;
	input wire C2;
	input wire C1;
	output wire Q;
	input wire CI;
	input wire B;
	input wire A;

endmodule // vdp_cnt_bit_rev

module vdp_2x_sr_bit (  Q, D, nC2, nC1, C2, C1, nC4, nC3, C4, C3);

	output wire Q;
	input wire D;
	input wire nC2;
	input wire nC1;
	input wire C2;
	input wire C1;
	input wire nC4;
	input wire nC3;
	input wire C4;
	input wire C3;

endmodule // vdp_2x_sr_bit

module vdp_and9 (  Z, B, A, C, D, F, E, G, H, I);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;
	input wire I;

endmodule // vdp_and9

module vdp_nor12 (  Z, B, A, C, D, F, E, G, H, J, I, K, L);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;
	input wire J;
	input wire I;
	input wire K;
	input wire L;

endmodule // vdp_nor12

module vdp_nor8 (  Z, B, A, C, D, F, E, G, H);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;

endmodule // vdp_nor8

module vdp_aon21_sr (  Q, A1, A2, B, nC2, nC1, C2, C1);

	output wire Q;
	input wire A1;
	input wire A2;
	input wire B;
	input wire nC2;
	input wire nC1;
	input wire C2;
	input wire C1;

endmodule // vdp_aon21_sr

module vdp_or9 (  Z, B, A, C, D, F, E, G, H, I);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;
	input wire I;

endmodule // vdp_or9

module vdp_V_PLA (  o0, o1, o2, o3, o4, o5, o6, o7, o8, o9, o10, o11, o12, o13, o14, o15, o16, o17, o18, o19, o20, o21, o22, o23, o24, o25, o26, o27, o28, o29, o30, o31, o32, o33, o34, o35, o36, o37, o38, o39, o40, o41, o42, o43, o44, o45, o46, o47, Vcnt0, Vcnt1, Vcnt2, Vcnt3, Vcnt4, Vcnt5, Vcnt6, Vcnt7, Vcnt8, ODD_EVEN, LS0, PAL, nPAL, i2, i3, M5);

	output wire o0;
	output wire o1;
	output wire o2;
	output wire o3;
	output wire o4;
	output wire o5;
	output wire o6;
	output wire o7;
	output wire o8;
	output wire o9;
	output wire o10;
	output wire o11;
	output wire o12;
	output wire o13;
	output wire o14;
	output wire o15;
	output wire o16;
	output wire o17;
	output wire o18;
	output wire o19;
	output wire o20;
	output wire o21;
	output wire o22;
	output wire o23;
	output wire o24;
	output wire o25;
	output wire o26;
	output wire o27;
	output wire o28;
	output wire o29;
	output wire o30;
	output wire o31;
	output wire o32;
	output wire o33;
	output wire o34;
	output wire o35;
	output wire o36;
	output wire o37;
	output wire o38;
	output wire o39;
	output wire o40;
	output wire o41;
	output wire o42;
	output wire o43;
	output wire o44;
	output wire o45;
	output wire o46;
	output wire o47;
	input wire Vcnt0;
	input wire Vcnt1;
	input wire Vcnt2;
	input wire Vcnt3;
	input wire Vcnt4;
	input wire Vcnt5;
	input wire Vcnt6;
	input wire Vcnt7;
	input wire Vcnt8;
	input wire ODD_EVEN;
	input wire LS0;
	input wire PAL;
	input wire nPAL;
	input wire i2;
	input wire i3;
	input wire M5;

endmodule // vdp_V_PLA

module vdp_cram (  q8, D8, q7, D7, q6, D6, q5, D5, q4, D4, q3, D3, q2, D2, q1, D1, q0, D0, A0, A1, CLK, A2, A3, A4, A5, Bi, Ai);

	output wire q8;
	input wire D8;
	output wire q7;
	input wire D7;
	output wire q6;
	input wire D6;
	output wire q5;
	input wire D5;
	output wire q4;
	input wire D4;
	output wire q3;
	input wire D3;
	output wire q2;
	input wire D2;
	output wire q1;
	input wire D1;
	output wire q0;
	input wire D0;
	input wire A0;
	input wire A1;
	input wire CLK;
	input wire A2;
	input wire A3;
	input wire A4;
	input wire A5;
	input wire Bi;
	input wire Ai;

endmodule // vdp_cram

module vdp_linebuf_ram (  q0, D0, q1, D1, q2, D2, q3, D3, q4, D4, q5, D5, q6, D6, q7, D7, q8, D8, q9, D9, q10, D10, q11, D11, q12, D12, q13, D13, q14, D14, q15, D15, q16, D16, q17, D17, q18, D18, q19, D19, q20, D20, q21, D21, q22, D22, q23, D23, q24, D24, q25, D25, q26, D26, q27, D27, CLK, A5, A4, A3, A2, A1, A0, Ai, Bi, Ci, Di);

	output wire q0;
	input wire D0;
	output wire q1;
	input wire D1;
	output wire q2;
	input wire D2;
	output wire q3;
	input wire D3;
	output wire q4;
	input wire D4;
	output wire q5;
	input wire D5;
	output wire q6;
	input wire D6;
	output wire q7;
	input wire D7;
	output wire q8;
	input wire D8;
	output wire q9;
	input wire D9;
	output wire q10;
	input wire D10;
	output wire q11;
	input wire D11;
	output wire q12;
	input wire D12;
	output wire q13;
	input wire D13;
	output wire q14;
	input wire D14;
	output wire q15;
	input wire D15;
	output wire q16;
	input wire D16;
	output wire q17;
	input wire D17;
	output wire q18;
	input wire D18;
	output wire q19;
	input wire D19;
	output wire q20;
	input wire D20;
	output wire q21;
	input wire D21;
	output wire q22;
	input wire D22;
	output wire q23;
	input wire D23;
	output wire q24;
	input wire D24;
	output wire q25;
	input wire D25;
	output wire q26;
	input wire D26;
	output wire q27;
	input wire D27;
	input wire CLK;
	input wire A5;
	input wire A4;
	input wire A3;
	input wire A2;
	input wire A1;
	input wire A0;
	input wire Ai;
	input wire Bi;
	input wire Ci;
	input wire Di;

endmodule // vdp_linebuf_ram

module vdp_att_cashe_ram2 (  q0, D0, q1, D1, q2, D2, q3, D3, q4, D4, q5, D5, q6, D6, q7, D7, q8, D8, q9, D9, q10, D10, CLK, A6, A5, A1, A0, A4, A3, A2, Ai, Bi);

	output wire q0;
	input wire D0;
	output wire q1;
	input wire D1;
	output wire q2;
	input wire D2;
	output wire q3;
	input wire D3;
	output wire q4;
	input wire D4;
	output wire q5;
	input wire D5;
	output wire q6;
	input wire D6;
	output wire q7;
	input wire D7;
	output wire q8;
	input wire D8;
	output wire q9;
	input wire D9;
	output wire q10;
	input wire D10;
	input wire CLK;
	input wire A6;
	input wire A5;
	input wire A1;
	input wire A0;
	input wire A4;
	input wire A3;
	input wire A2;
	input wire Ai;
	input wire Bi;

endmodule // vdp_att_cashe_ram2

module vdp_att_cashe_ram1 (  q0, D0, q1, D1, q2, D2, q3, D3, q4, D4, q5, D5, q6, D6, q7, D7, q8, D8, q9, D9, CLK, A0, A1, A2, A3, A4, A5, A6, Ai, Bi);

	output wire q0;
	input wire D0;
	output wire q1;
	input wire D1;
	output wire q2;
	input wire D2;
	output wire q3;
	input wire D3;
	output wire q4;
	input wire D4;
	output wire q5;
	input wire D5;
	output wire q6;
	input wire D6;
	output wire q7;
	input wire D7;
	output wire q8;
	input wire D8;
	output wire q9;
	input wire D9;
	input wire CLK;
	input wire A0;
	input wire A1;
	input wire A2;
	input wire A3;
	input wire A4;
	input wire A5;
	input wire A6;
	input wire Ai;
	input wire Bi;

endmodule // vdp_att_cashe_ram1

module vdp_att_temp_ram (  A4, A0, A1, A2, A3, q0, D0, q1, D1, q2, D2, q3, D3, q4, D4, q5, D5, q6, D6, q7, D7, q8, D8, q9, D9, q10, D10, q11, D11, q12, D12, q13, D13, q14, D14, q15, D15, q16, D16, q17, D17, q18, D18, q19, D19, q20, D20, q21, D21, q22, D22, q23, D23, q24, D24, q25, D25, q26, D26, q26, D26, q27, D27, q28, D28, q29, D29, q30, D30, q31, D[31], q32, D32, CLK, Ai, Bi, Ci);

	input wire A4;
	input wire A0;
	input wire A1;
	input wire A2;
	input wire A3;
	output wire q0;
	input wire D0;
	output wire q1;
	input wire D1;
	output wire q2;
	input wire D2;
	output wire q3;
	input wire D3;
	output wire q4;
	input wire D4;
	output wire q5;
	input wire D5;
	output wire q6;
	input wire D6;
	output wire q7;
	input wire D7;
	output wire q8;
	input wire D8;
	output wire q9;
	input wire D9;
	output wire q10;
	input wire D10;
	output wire q11;
	input wire D11;
	output wire q12;
	input wire D12;
	output wire q13;
	input wire D13;
	output wire q14;
	input wire D14;
	output wire q15;
	input wire D15;
	output wire q16;
	input wire D16;
	output wire q17;
	input wire D17;
	output wire q18;
	input wire D18;
	output wire q19;
	input wire D19;
	output wire q20;
	input wire D20;
	output wire q21;
	input wire D21;
	output wire q22;
	input wire D22;
	output wire q23;
	input wire D23;
	output wire q24;
	input wire D24;
	output wire q25;
	input wire D25;
	output wire q26;
	input wire D26;
	output wire q26;
	input wire D26;
	output wire q27;
	input wire D27;
	output wire q28;
	input wire D28;
	output wire q29;
	input wire D29;
	output wire q30;
	input wire D30;
	output wire q31;
	input wire D[31];
	output wire q32;
	input wire D32;
	input wire CLK;
	input wire Ai;
	input wire Bi;
	input wire Ci;

endmodule // vdp_att_temp_ram

module vdp_vsram (  CLK, D10, q10, D9, q9, D8, q8, D7, q7, D6, q6, D5, q5, D4, q4, D3, q3, D2, q2, D1, q1, D0, q0, A1, A2, A3, A4, A5, A0, Ai, Bi);

	input wire CLK;
	input wire D10;
	output wire q10;
	input wire D9;
	output wire q9;
	input wire D8;
	output wire q8;
	input wire D7;
	output wire q7;
	input wire D6;
	output wire q6;
	input wire D5;
	output wire q5;
	input wire D4;
	output wire q4;
	input wire D3;
	output wire q3;
	input wire D2;
	output wire q2;
	input wire D1;
	output wire q1;
	input wire D0;
	output wire q0;
	input wire A1;
	input wire A2;
	input wire A3;
	input wire A4;
	input wire A5;
	input wire A0;
	input wire Ai;
	input wire Bi;

endmodule // vdp_vsram

module vdp_H_PLA (  HPLA0, HPLA1, HPLA2, HPLA3, HPLA4, HPLA5, HPLA7, HPLA8, HPLA9, HPLA6, HPLA10, HPLA11, HPLA16, HPLA15, HPLA14, HPLA13, HPLA12, i0, HPLA17, HPLA18, HPLA19, HPLA20, HPLA21, HPLA22, Hcnt0, Hcnt1, Hcnt2, Hcnt3, Hcnt4, Hcnt5, Hcnt6, Hcnt7, Hcnt8, H40, M5, B, C, A, HPLA[23], HPLA[24], HPLA[25], HPLA[26], HPLA[27], HPLA[28], HPLA[29], HPLA[30], HPLA[31], HPLA[32], HPLA[33], i3, HPLA[35], HPLA[36], HPLA[34]);

	output wire HPLA0;
	output wire HPLA1;
	output wire HPLA2;
	output wire HPLA3;
	output wire HPLA4;
	output wire HPLA5;
	output wire HPLA7;
	output wire HPLA8;
	output wire HPLA9;
	output wire HPLA6;
	output wire HPLA10;
	output wire HPLA11;
	output wire HPLA16;
	output wire HPLA15;
	output wire HPLA14;
	output wire HPLA13;
	output wire HPLA12;
	input wire i0;
	output wire HPLA17;
	output wire HPLA18;
	output wire HPLA19;
	output wire HPLA20;
	output wire HPLA21;
	output wire HPLA22;
	input wire Hcnt0;
	input wire Hcnt1;
	input wire Hcnt2;
	input wire Hcnt3;
	input wire Hcnt4;
	input wire Hcnt5;
	input wire Hcnt6;
	input wire Hcnt7;
	input wire Hcnt8;
	input wire H40;
	input wire M5;
	input wire B;
	input wire C;
	input wire A;
	output wire HPLA[23];
	output wire HPLA[24];
	output wire HPLA[25];
	output wire HPLA[26];
	output wire HPLA[27];
	output wire HPLA[28];
	output wire HPLA[29];
	output wire HPLA[30];
	output wire HPLA[31];
	output wire HPLA[32];
	output wire HPLA[33];
	input wire i3;
	output wire HPLA[35];
	output wire HPLA[36];
	output wire HPLA[34];

endmodule // vdp_H_PLA



// ERROR: conflicting wire AD_DATA[7]
// ERROR: conflicting wire AD_DATA[6]
// ERROR: conflicting wire AD_DATA[4]
// ERROR: conflicting wire RD_DATA[2]
// ERROR: conflicting wire RD_DATA[1]
// ERROR: conflicting wire RD_DATA[0]
// ERROR: conflicting wire AD_DATA[5]
// ERROR: conflicting wire DB[0]
// ERROR: conflicting wire DB[1]
// ERROR: conflicting wire DB[2]
// ERROR: conflicting wire DB[3]
// ERROR: conflicting wire DB[4]
// ERROR: conflicting wire DB[5]
// ERROR: conflicting wire DB[6]
// ERROR: conflicting wire DB[7]
// ERROR: conflicting wire DB[8]
// ERROR: conflicting wire DB[9]
// ERROR: conflicting wire AD_DATA[3]
// ERROR: conflicting wire AD_DATA[2]
// ERROR: conflicting wire AD_DATA[1]
// ERROR: conflicting wire AD_DATA[0]
// ERROR: conflicting wire DB[14]
// ERROR: conflicting wire DB[13]
// ERROR: conflicting wire DB[12]
// ERROR: conflicting wire DB[11]
// ERROR: conflicting wire DB[10]
// ERROR: floating wire w188
// ERROR: conflicting wire RD_DATA[4]
// ERROR: floating wire w219
// ERROR: conflicting wire RD_DATA[6]
// ERROR: floating wire w235
// ERROR: conflicting wire w237
// ERROR: conflicting wire w245
// ERROR: conflicting wire w254
// ERROR: conflicting wire w262
// ERROR: conflicting wire w279
// ERROR: conflicting wire w288
// ERROR: conflicting wire w297
// ERROR: conflicting wire w305
// ERROR: conflicting wire w321
// ERROR: floating wire w334
// ERROR: conflicting wire RD_DATA[5]
// ERROR: floating wire w350
// ERROR: conflicting wire DB[15]
// ERROR: conflicting wire w355
// ERROR: floating wire w449
// ERROR: conflicting wire VRAMA[0]
// ERROR: floating wire w561
// ERROR: conflicting wire VRAMA[8]
// ERROR: conflicting wire VRAMA[7]
// ERROR: conflicting wire VRAMA[9]
// ERROR: conflicting wire VRAMA[10]
// ERROR: conflicting wire VRAMA[6]
// ERROR: conflicting wire VRAMA[5]
// ERROR: conflicting wire VRAMA[11]
// ERROR: conflicting wire VRAMA[12]
// ERROR: conflicting wire VRAMA[4]
// ERROR: conflicting wire VRAMA[13]
// ERROR: conflicting wire VRAMA[3]
// ERROR: conflicting wire VRAMA[14]
// ERROR: conflicting wire VRAMA[2]
// ERROR: conflicting wire VRAMA[15]
// ERROR: conflicting wire VRAMA[1]
// ERROR: conflicting wire VRAMA[16]
// ERROR: floating wire w774
// ERROR: floating wire w776
// ERROR: floating wire w789
// ERROR: floating wire w790
// ERROR: floating wire w1040
// ERROR: conflicting wire COL[1]
// ERROR: conflicting wire COL[0]
// ERROR: conflicting wire COL[2]
// ERROR: conflicting wire COL[3]
// ERROR: conflicting wire COL[4]
// ERROR: conflicting wire COL[6]
// ERROR: conflicting wire COL[5]
// ERROR: floating wire w1060
// ERROR: floating wire w1061
// ERROR: floating wire w1183
// ERROR: floating wire w1254
// ERROR: floating wire w1261
// ERROR: floating wire w1269
// ERROR: floating wire w1285
// ERROR: floating wire w1314
// ERROR: floating wire w1338
// ERROR: floating wire w1555
// ERROR: floating wire w1623
// ERROR: floating wire w1722
// ERROR: floating wire w1752
// ERROR: floating wire w1765
// ERROR: floating wire w1775
// ERROR: floating wire w1908
// ERROR: floating wire w1999
// ERROR: floating wire w2185
// ERROR: floating wire w2220
// ERROR: floating wire w2397
// ERROR: floating wire w2541
// ERROR: floating wire w2547
// ERROR: floating wire w2701
// ERROR: floating wire w3004
// ERROR: floating wire w3014
// ERROR: floating wire w3350
// ERROR: floating wire w3408
// ERROR: floating wire w3488
// ERROR: floating wire w3544
// ERROR: floating wire w3585
// ERROR: floating wire w3626
// ERROR: floating wire w3631
// ERROR: floating wire w3685
// ERROR: floating wire w3687
// ERROR: floating wire w3760
// ERROR: floating wire con0
// ERROR: floating wire w3837
// ERROR: floating wire w3951
// ERROR: floating wire w4282
// ERROR: floating wire w4291
// ERROR: floating wire w4443
// ERROR: floating wire w4505
// ERROR: floating wire w4510
// ERROR: floating wire w4547
// ERROR: floating wire w4606
// ERROR: floating wire w4611
// ERROR: floating wire w4640
// ERROR: floating wire w4685
// ERROR: floating wire w4744
// ERROR: floating wire w4751
// ERROR: floating wire w4796
// ERROR: floating wire w4981
// ERROR: floating wire w5036
// ERROR: floating wire w5163
// ERROR: floating wire w5171
// ERROR: floating wire w5185
// ERROR: floating wire w5331
// ERROR: floating wire w5379
// ERROR: floating wire w5565
// ERROR: floating wire w5702
// ERROR: floating wire w5704
// ERROR: floating wire w5799
// ERROR: floating wire w5941
// ERROR: floating wire w5956
// ERROR: floating wire w5987
// ERROR: floating wire w6032
// ERROR: floating wire w6079
// ERROR: floating wire w6080
// ERROR: floating wire w6324
// ERROR: floating wire w6439
// ERROR: floating wire w6441
// ERROR: floating wire w6442
// ERROR: floating wire w6537
// ERROR: floating wire w6589
// WARNING: Cell vdp_fa:g385 port CO not connected.
// WARNING: Cell vdp_and:g527 port Z not connected.
// WARNING: Cell vdp_cnt_bit_load:g871 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g873 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g1405 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g1406 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1407 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1408 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1409 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1410 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1411 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1412 port Q not connected.
// WARNING: Cell vdp_or:g1576 port Z not connected.
// WARNING: Cell vdp_cnt_bit_load:g1959 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g1960 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2145 port CO not connected.
// WARNING: Cell vdp_ha:g2278 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2280 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2282 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2284 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2286 port CO not connected.
// WARNING: Cell vdp_rs_ff:g2380 port nQ not connected.
// WARNING: Cell vdp_rs_ff:g2381 port nQ not connected.
// WARNING: Cell vdp_comp_we:g2612 port nZ not connected.
// WARNING: Cell vdp_comp_we:g2701 port nZ not connected.
// WARNING: Cell vdp_fa:g3842 port CO not connected.
// WARNING: Cell vdp_fa:g4058 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g4437 port CO not connected.
// WARNING: Cell vdp_fa:g4453 port CO not connected.
// WARNING: Cell vdp_fa:g4463 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g5851 port CO not connected.
// WARNING: Cell vdp_fa:g5862 port CO not connected.
// WARNING: Cell vdp_fa:g5888 port CO not connected.
// WARNING: Cell vdp_fa:g5892 port CO not connected.
// WARNING: Cell vdp_fa:g6086 port CO not connected.
// WARNING: Cell vdp_ha:g6137 port CO not connected.
// WARNING: Cell vdp_sr_bit:g6146 port Q not connected.
// WARNING: Cell vdp_fa:g6150 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g6216 port CO not connected.
