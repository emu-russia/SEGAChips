module VDP (  CH0_EN, CH0VOL[0], CH0VOL[1], CH1_EN, CH1VOL[0], CH1VOL[1], CH2_EN, CH2VOL[0], CH2VOL[1], CH3_EN, CH3VOL[0], CH3VOL[1], PSGDAC0[0], PSGDAC0[1], PSGDAC0[2], PSGDAC0[3], PSGDAC0[4], PSGDAC0[5], PSGDAC0[6], PSGDAC0[7], PSGDAC1[0], PSGDAC1[1], PSGDAC1[2], PSGDAC1[3], PSGDAC1[4], PSGDAC1[5], PSGDAC1[6], PSGDAC1[7], PSGDAC2[0], PSGDAC2[1], PSGDAC2[2], PSGDAC2[3], PSGDAC2[4], PSGDAC2[5], PSGDAC2[6], PSGDAC2[7], PSGDAC3[0], PSGDAC3[1], PSGDAC3[2], PSGDAC3[3], PSGDAC3[4], PSGDAC3[5], PSGDAC3[6], PSGDAC3[7], CAi[22], CAo[22], CA[19], DTACK_OUT, Z80_INT, RA[7], RA[6], RA[5], RA[4], RA[2], RA[1], RA[0], nRAS0, RA[3], nCAS0, nOE0, nLWR, nUWR, DTACK_IN, RnW, nLDS, nUDS, nAS, nM1, nWR, nRD, nIORQ, nILP2, nILP1, nINTAK, nMREQ, nBG, BGACK_OUT, BGACK_IN, nBR, VSYNC, nCSYNC, nCSYNC_IN, nHSYNC, nHSYNC_IN, DB[15], DB[14], DB[13], DB[12], DB[11], DB[10], DB[9], DB[8], DB[7], DB[6], DB[5], DB[4], DB[3], DB[2], DB[1], DB[0], CA[0], CA[1], CA[2], CA[3], CA[4], CA[5], CA[6], CA[7], CA[8], CA[9], CA[10], CA[11], CA[12], CA[13], CA[14], CA[15], CA[16], CA[17], CA[18], CA[20], CA[21], R_DAC[0], R_DAC[1], R_DAC[2], R_DAC[3], R_DAC[4], R_DAC[5], R_DAC[6], R_DAC[7], R_DAC[8], G_DAC[0], G_DAC[1], G_DAC[2], G_DAC[3], G_DAC[4], G_DAC[5], G_DAC[6], G_DAC[7], G_DAC[8], R_DAC[9], R_DAC[10], R_DAC[11], R_DAC[12], R_DAC[13], R_DAC[14], R_DAC[15], R_DAC[16], B_DAC[0], B_DAC[1], B_DAC[2], B_DAC[3], B_DAC[4], B_DAC[5], B_DAC[6], B_DAC[7], B_DAC[8], G_DAC[9], G_DAC[10], G_DAC[11], G_DAC[12], G_DAC[13], G_DAC[14], G_DAC[15], G_DAC[16], B_DAC[9], B_DAC[10], B_DAC[11], B_DAC[12], B_DAC[13], B_DAC[14], B_DAC[15], B_DAC[16], nOE1, nWE0, nWE1, nCAS1, nRAS1, AD_RD_DIR, nYS, nSC, nSE0_1, ADo[7], ADo[6], ADo[5], ADo[4], ADo[3], ADo[2], ADo[1], ADo[0], RDo[6], RDo[5], RDo[4], RDo[3], RDo[2], RDo[1], RDo[0], RDi[6], RDi[7], RDi[4], RDi[5], RDi[2], RDi[3], RDi[0], RDi[1], ADi[6], ADi[7], ADi[4], ADi[5], ADi[2], ADi[3], ADi[0], ADi[1], RDo[7], SD[7], SD[6], SD[5], SD[4], SD[3], SD[2], SD[1], SD[0], CLK1, CLK0, EDCLKi, EDCLKo, MCLK, SUB_CLK, nRES_PAD, M68kCLKi, EDCLKd, CA_PAD_DIR, DB_PAD_DIR, nSEL0_M3, nPAL, nHL, SPA_Bo, SPA_Bi);

	output wire CH0_EN;
	output wire CH0VOL[0];
	output wire CH0VOL[1];
	output wire CH1_EN;
	output wire CH1VOL[0];
	output wire CH1VOL[1];
	output wire CH2_EN;
	output wire CH2VOL[0];
	output wire CH2VOL[1];
	output wire CH3_EN;
	output wire CH3VOL[0];
	output wire CH3VOL[1];
	output wire PSGDAC0[0];
	output wire PSGDAC0[1];
	output wire PSGDAC0[2];
	output wire PSGDAC0[3];
	output wire PSGDAC0[4];
	output wire PSGDAC0[5];
	output wire PSGDAC0[6];
	output wire PSGDAC0[7];
	output wire PSGDAC1[0];
	output wire PSGDAC1[1];
	output wire PSGDAC1[2];
	output wire PSGDAC1[3];
	output wire PSGDAC1[4];
	output wire PSGDAC1[5];
	output wire PSGDAC1[6];
	output wire PSGDAC1[7];
	output wire PSGDAC2[0];
	output wire PSGDAC2[1];
	output wire PSGDAC2[2];
	output wire PSGDAC2[3];
	output wire PSGDAC2[4];
	output wire PSGDAC2[5];
	output wire PSGDAC2[6];
	output wire PSGDAC2[7];
	output wire PSGDAC3[0];
	output wire PSGDAC3[1];
	output wire PSGDAC3[2];
	output wire PSGDAC3[3];
	output wire PSGDAC3[4];
	output wire PSGDAC3[5];
	output wire PSGDAC3[6];
	output wire PSGDAC3[7];
	input wire CAi[22];
	output wire CAo[22];
	output wire CA[19];
	output wire DTACK_OUT;
	output wire Z80_INT;
	output wire RA[7];
	output wire RA[6];
	output wire RA[5];
	output wire RA[4];
	output wire RA[2];
	output wire RA[1];
	output wire RA[0];
	output wire nRAS0;
	output wire RA[3];
	output wire nCAS0;
	output wire nOE0;
	output wire nLWR;
	output wire nUWR;
	input wire DTACK_IN;
	input wire RnW;
	input wire nLDS;
	input wire nUDS;
	input wire nAS;
	input wire nM1;
	input wire nWR;
	input wire nRD;
	input wire nIORQ;
	output wire nILP2;
	output wire nILP1;
	input wire nINTAK;
	input wire nMREQ;
	input wire nBG;
	output wire BGACK_OUT;
	input wire BGACK_IN;
	output wire nBR;
	output wire VSYNC;
	output wire nCSYNC;
	input wire nCSYNC_IN;
	output wire nHSYNC;
	input wire nHSYNC_IN;
	inout wire DB[15];
	inout wire DB[14];
	inout wire DB[13];
	inout wire DB[12];
	inout wire DB[11];
	inout wire DB[10];
	inout wire DB[9];
	inout wire DB[8];
	inout wire DB[7];
	inout wire DB[6];
	inout wire DB[5];
	inout wire DB[4];
	inout wire DB[3];
	inout wire DB[2];
	inout wire DB[1];
	inout wire DB[0];
	inout wire CA[0];
	inout wire CA[1];
	inout wire CA[2];
	inout wire CA[3];
	inout wire CA[4];
	inout wire CA[5];
	inout wire CA[6];
	inout wire CA[7];
	inout wire CA[8];
	inout wire CA[9];
	inout wire CA[10];
	inout wire CA[11];
	inout wire CA[12];
	inout wire CA[13];
	inout wire CA[14];
	inout wire CA[15];
	inout wire CA[16];
	inout wire CA[17];
	output wire CA[18];
	inout wire CA[20];
	inout wire CA[21];
	output wire R_DAC[0];
	output wire R_DAC[1];
	output wire R_DAC[2];
	output wire R_DAC[3];
	output wire R_DAC[4];
	output wire R_DAC[5];
	output wire R_DAC[6];
	output wire R_DAC[7];
	output wire R_DAC[8];
	output wire G_DAC[0];
	output wire G_DAC[1];
	output wire G_DAC[2];
	output wire G_DAC[3];
	output wire G_DAC[4];
	output wire G_DAC[5];
	output wire G_DAC[6];
	output wire G_DAC[7];
	output wire G_DAC[8];
	output wire R_DAC[9];
	output wire R_DAC[10];
	output wire R_DAC[11];
	output wire R_DAC[12];
	output wire R_DAC[13];
	output wire R_DAC[14];
	output wire R_DAC[15];
	output wire R_DAC[16];
	output wire B_DAC[0];
	output wire B_DAC[1];
	output wire B_DAC[2];
	output wire B_DAC[3];
	output wire B_DAC[4];
	output wire B_DAC[5];
	output wire B_DAC[6];
	output wire B_DAC[7];
	output wire B_DAC[8];
	output wire G_DAC[9];
	output wire G_DAC[10];
	output wire G_DAC[11];
	output wire G_DAC[12];
	output wire G_DAC[13];
	output wire G_DAC[14];
	output wire G_DAC[15];
	output wire G_DAC[16];
	output wire B_DAC[9];
	output wire B_DAC[10];
	output wire B_DAC[11];
	output wire B_DAC[12];
	output wire B_DAC[13];
	output wire B_DAC[14];
	output wire B_DAC[15];
	output wire B_DAC[16];
	output wire nOE1;
	output wire nWE0;
	output wire nWE1;
	output wire nCAS1;
	output wire nRAS1;
	output wire AD_RD_DIR;
	output wire nYS;
	output wire nSC;
	output wire nSE0_1;
	output wire ADo[7];
	output wire ADo[6];
	output wire ADo[5];
	output wire ADo[4];
	output wire ADo[3];
	output wire ADo[2];
	output wire ADo[1];
	output wire ADo[0];
	output wire RDo[6];
	output wire RDo[5];
	output wire RDo[4];
	output wire RDo[3];
	output wire RDo[2];
	output wire RDo[1];
	output wire RDo[0];
	input wire RDi[6];
	input wire RDi[7];
	input wire RDi[4];
	input wire RDi[5];
	input wire RDi[2];
	input wire RDi[3];
	input wire RDi[0];
	input wire RDi[1];
	input wire ADi[6];
	input wire ADi[7];
	input wire ADi[4];
	input wire ADi[5];
	input wire ADi[2];
	input wire ADi[3];
	input wire ADi[0];
	input wire ADi[1];
	output wire RDo[7];
	input wire SD[7];
	input wire SD[6];
	input wire SD[5];
	input wire SD[4];
	input wire SD[3];
	input wire SD[2];
	input wire SD[1];
	input wire SD[0];
	output wire CLK1;
	output wire CLK0;
	input wire EDCLKi;
	output wire EDCLKo;
	input wire MCLK;
	output wire SUB_CLK;
	input wire nRES_PAD;
	input wire M68kCLKi;
	output wire EDCLKd;
	output wire CA_PAD_DIR;
	output wire DB_PAD_DIR;
	input wire nSEL0_M3;
	input wire nPAL;
	input wire nHL;
	output wire SPA_Bo;
	input wire SPA_Bi;

	// Wires

	wire w1;
	wire H40;
	wire w3;
	wire w4;
	wire w5;
	wire w6;
	wire w7;
	wire w8;
	wire w9;
	wire w10;
	wire w11;
	wire w12;
	wire w13;
	wire w14;
	wire w15;
	wire w16;
	wire w17;
	wire w18;
	wire w19;
	wire w20;
	wire w21;
	wire w22;
	wire w23;
	wire w24;
	wire w25;
	wire w26;
	wire w27;
	wire w28;
	wire w29;
	wire w30;
	wire w31;
	wire w32;
	wire w33;
	wire w34;
	wire w35;
	wire w36;
	wire w37;
	wire w38;
	wire w39;
	wire w40;
	wire VSCR;
	wire w42;
	wire w43;
	wire w44;
	wire w45;
	wire ODD_EVEN;
	wire w47;
	wire w48;
	wire w49;
	wire w50;
	wire w51;
	wire w52;
	wire w53;
	wire w54;
	wire w55;
	wire w56;
	wire FIFOo[7];
	wire FIFOo[6];
	wire FIFOo[5];
	wire FIFOo[4];
	wire FIFOo[3];
	wire FIFOo[2];
	wire FIFOo[1];
	wire FIFOo[0];
	wire w65;
	wire w66;
	wire w67;
	wire w68;
	wire w69;
	wire w70;
	wire w71;
	wire w72;
	wire w73;
	wire S_TE;
	wire w75;
	wire LSCR;
	wire w77;
	wire HSCR;
	wire w79;
	wire w80;
	wire w81;
	wire w82;
	wire w83;
	wire w84;
	wire w85;
	wire w86;
	wire VPOS[9];
	wire w88;
	wire w89;
	wire w90;
	wire w91;
	wire HPOS[0];
	wire w93;
	wire w94;
	wire w95;
	wire V_INT_HAPPENED;
	wire w97;
	wire w98;
	wire w99;
	wire w100;
	wire VPOS[8];
	wire w102;
	wire COLLISION;
	wire w104;
	wire w105;
	wire w106;
	wire w107;
	wire w108;
	wire w109;
	wire SPRITE_OVF;
	wire w111;
	wire w112;
	wire w113;
	wire w114;
	wire COL[7];
	wire w116;
	wire w117;
	wire w118;
	wire w119;
	wire AD_DATA[7];
	wire AD_DATA[6];
	wire AD_DATA[4];
	wire RD_DATA[2];
	wire RD_DATA[1];
	wire RD_DATA[0];
	wire AD_DATA[5];
	wire DCLK1;
	wire DCLK2;
	wire nDCLK1;
	wire nDCLK2;
	wire HCLK1;
	wire HCLK2;
	wire nHCLK1;
	wire nHCLK2;
	wire SYSRES;
	wire DB[0];
	wire DB[1];
	wire DB[2];
	wire DB[3];
	wire DB[4];
	wire DB[5];
	wire DB[6];
	wire DB[7];
	wire DB[8];
	wire DB[9];
	wire AD_DATA[3];
	wire AD_DATA[2];
	wire AD_DATA[1];
	wire AD_DATA[0];
	wire DB[14];
	wire DB[13];
	wire DB[12];
	wire DB[11];
	wire DB[10];
	wire M5;
	wire w156;
	wire w157;
	wire VPOS_80;
	wire w159;
	wire HPOS[1];
	wire w161;
	wire w162;
	wire w163;
	wire w164;
	wire w165;
	wire w166;
	wire w167;
	wire w168;
	wire w169;
	wire w170;
	wire w171;
	wire w172;
	wire VPOS[2];
	wire w174;
	wire HPOS[3];
	wire w176;
	wire w177;
	wire w178;
	wire w179;
	wire w180;
	wire w181;
	wire w182;
	wire w183;
	wire w184;
	wire w185;
	wire w186;
	wire w187;
	wire VPOS[4];
	wire w189;
	wire RD_DATA[4];
	wire HPOS[5];
	wire w192;
	wire w193;
	wire w194;
	wire w195;
	wire w196;
	wire w197;
	wire w198;
	wire w199;
	wire w200;
	wire w201;
	wire w202;
	wire w203;
	wire w204;
	wire RD_DATA[6];
	wire HPOS[7];
	wire w207;
	wire w208;
	wire w209;
	wire w210;
	wire w211;
	wire w212;
	wire w213;
	wire w214;
	wire w215;
	wire w216;
	wire w217;
	wire w218;
	wire w219;
	wire w220;
	wire w221;
	wire w222;
	wire w223;
	wire w224;
	wire w225;
	wire w226;
	wire w227;
	wire w228;
	wire w229;
	wire w230;
	wire w231;
	wire w232;
	wire w233;
	wire w234;
	wire w235;
	wire w236;
	wire w237;
	wire w238;
	wire w239;
	wire w240;
	wire w241;
	wire w242;
	wire w243;
	wire w244;
	wire w245;
	wire w246;
	wire w247;
	wire w248;
	wire w249;
	wire w250;
	wire w251;
	wire w252;
	wire w253;
	wire w254;
	wire w255;
	wire w256;
	wire w257;
	wire w258;
	wire w259;
	wire w260;
	wire w261;
	wire w262;
	wire w263;
	wire w264;
	wire w265;
	wire w266;
	wire w267;
	wire w268;
	wire w269;
	wire w270;
	wire w271;
	wire w272;
	wire w273;
	wire w274;
	wire w275;
	wire w276;
	wire w277;
	wire w278;
	wire w279;
	wire w280;
	wire w281;
	wire w282;
	wire w283;
	wire w284;
	wire w285;
	wire VPOS[1];
	wire HPOS[2];
	wire w288;
	wire w289;
	wire w290;
	wire w291;
	wire w292;
	wire w293;
	wire w294;
	wire w295;
	wire w296;
	wire w297;
	wire w298;
	wire VPOS[3];
	wire w300;
	wire HPOS[4];
	wire w302;
	wire w303;
	wire w304;
	wire w305;
	wire w306;
	wire w307;
	wire w308;
	wire w309;
	wire w310;
	wire w311;
	wire w312;
	wire w313;
	wire w314;
	wire VPOS[5];
	wire RD_DATA[5];
	wire HPOS[6];
	wire w318;
	wire w319;
	wire w320;
	wire w321;
	wire w322;
	wire w323;
	wire w324;
	wire w325;
	wire w326;
	wire w327;
	wire w328;
	wire w329;
	wire w330;
	wire VPOS[7];
	wire DB[15];
	wire HPOS[8];
	wire w334;
	wire w335;
	wire w336;
	wire w337;
	wire w338;
	wire w339;
	wire w340;
	wire w341;
	wire w342;
	wire w343;
	wire w344;
	wire w345;
	wire w346;
	wire w347;
	wire w348;
	wire w349;
	wire w350;
	wire w351;
	wire w352;
	wire w353;
	wire w354;
	wire w355;
	wire w356;
	wire w357;
	wire w358;
	wire w359;
	wire w360;
	wire w361;
	wire w362;
	wire w363;
	wire w364;
	wire w365;
	wire w366;
	wire w367;
	wire w368;
	wire w369;
	wire w370;
	wire w371;
	wire w372;
	wire w373;
	wire nSEL0_M3;
	wire w375;
	wire w376;
	wire w377;
	wire w378;
	wire w379;
	wire w380;
	wire w381;
	wire w382;
	wire w383;
	wire w384;
	wire w385;
	wire w386;
	wire w387;
	wire w388;
	wire w389;
	wire w390;
	wire w391;
	wire w392;
	wire w393;
	wire w394;
	wire w395;
	wire w396;
	wire w397;
	wire w398;
	wire w399;
	wire w400;
	wire w401;
	wire w402;
	wire VRAM128k;
	wire w404;
	wire w405;
	wire w406;
	wire w407;
	wire w408;
	wire w409;
	wire w410;
	wire w411;
	wire w412;
	wire w413;
	wire w414;
	wire w415;
	wire w416;
	wire w417;
	wire w418;
	wire w419;
	wire w420;
	wire w421;
	wire w422;
	wire w423;
	wire w424;
	wire w425;
	wire w426;
	wire w427;
	wire w428;
	wire w429;
	wire w430;
	wire w431;
	wire w432;
	wire w433;
	wire w434;
	wire CD[2];
	wire CD[3];
	wire w437;
	wire w438;
	wire CA[0];
	wire w440;
	wire M3;
	wire w442;
	wire w443;
	wire w444;
	wire w445;
	wire w446;
	wire w447;
	wire w448;
	wire w449;
	wire w450;
	wire w451;
	wire w452;
	wire w453;
	wire w454;
	wire w455;
	wire w456;
	wire w457;
	wire w458;
	wire w459;
	wire w460;
	wire w461;
	wire CD[1];
	wire w463;
	wire w464;
	wire w465;
	wire w466;
	wire w467;
	wire w468;
	wire w469;
	wire w470;
	wire w471;
	wire w472;
	wire w473;
	wire w474;
	wire w475;
	wire CD[0];
	wire w477;
	wire w478;
	wire w479;
	wire w480;
	wire w481;
	wire w482;
	wire w483;
	wire w484;
	wire w485;
	wire w486;
	wire w487;
	wire w488;
	wire w489;
	wire w490;
	wire w491;
	wire w492;
	wire w493;
	wire w494;
	wire w495;
	wire w496;
	wire w497;
	wire w498;
	wire w499;
	wire w500;
	wire w501;
	wire w502;
	wire w503;
	wire w504;
	wire w505;
	wire w506;
	wire w507;
	wire w508;
	wire w509;
	wire w510;
	wire w511;
	wire w512;
	wire w513;
	wire w514;
	wire w515;
	wire w516;
	wire w517;
	wire w518;
	wire w519;
	wire w520;
	wire w521;
	wire w522;
	wire w523;
	wire w524;
	wire w525;
	wire w526;
	wire w527;
	wire w528;
	wire VRAMA[0];
	wire w530;
	wire w531;
	wire w532;
	wire w533;
	wire w534;
	wire w535;
	wire w536;
	wire w537;
	wire w538;
	wire w539;
	wire w540;
	wire w541;
	wire w542;
	wire w543;
	wire w544;
	wire w545;
	wire w546;
	wire w547;
	wire w548;
	wire w549;
	wire w550;
	wire w551;
	wire w552;
	wire w553;
	wire FIFO_EMPTY;
	wire w555;
	wire w556;
	wire w557;
	wire w558;
	wire w559;
	wire w560;
	wire w561;
	wire w562;
	wire w563;
	wire DMA_BUSY;
	wire w565;
	wire w566;
	wire w567;
	wire w568;
	wire w569;
	wire w570;
	wire w571;
	wire REG_BUS[0];
	wire w573;
	wire w574;
	wire w575;
	wire w576;
	wire w577;
	wire w578;
	wire w579;
	wire w580;
	wire w581;
	wire w582;
	wire w583;
	wire REG_BUS[7];
	wire w585;
	wire w586;
	wire w587;
	wire w588;
	wire w589;
	wire w590;
	wire w591;
	wire w592;
	wire w593;
	wire w594;
	wire w595;
	wire w596;
	wire VRAMA[8];
	wire w598;
	wire w599;
	wire w600;
	wire w601;
	wire CA[8];
	wire CA[7];
	wire w604;
	wire w605;
	wire w606;
	wire w607;
	wire w608;
	wire w609;
	wire w610;
	wire w611;
	wire w612;
	wire w613;
	wire w614;
	wire w615;
	wire CA[9];
	wire w617;
	wire VRAMA[7];
	wire w619;
	wire REG_BUS[6];
	wire VRAMA[9];
	wire w622;
	wire CA[6];
	wire w624;
	wire w625;
	wire w626;
	wire w627;
	wire w628;
	wire w629;
	wire w630;
	wire w631;
	wire w632;
	wire w633;
	wire w634;
	wire w635;
	wire w636;
	wire w637;
	wire REG_BUS[5];
	wire VRAMA[10];
	wire VRAMA[6];
	wire w641;
	wire REG_BUS[1];
	wire w643;
	wire w644;
	wire w645;
	wire w646;
	wire CA[10];
	wire w648;
	wire w649;
	wire w650;
	wire w651;
	wire w652;
	wire w653;
	wire REG_BUS[2];
	wire w655;
	wire CA[11];
	wire w657;
	wire w658;
	wire w659;
	wire w660;
	wire w661;
	wire w662;
	wire w663;
	wire w664;
	wire w665;
	wire VRAMA[5];
	wire w667;
	wire w668;
	wire VRAMA[11];
	wire CA[5];
	wire w671;
	wire w672;
	wire w673;
	wire REG_BUS[3];
	wire VRAMA[12];
	wire VRAMA[4];
	wire w677;
	wire w678;
	wire w679;
	wire REG_BUS[4];
	wire w681;
	wire CA[12];
	wire w683;
	wire w684;
	wire CA[4];
	wire w686;
	wire w687;
	wire w688;
	wire w689;
	wire CA[19];
	wire w691;
	wire w692;
	wire w693;
	wire w694;
	wire VRAMA[13];
	wire w696;
	wire w697;
	wire w698;
	wire VRAMA[3];
	wire CA[3];
	wire w701;
	wire w702;
	wire CA[13];
	wire CA[20];
	wire w705;
	wire w706;
	wire w707;
	wire w708;
	wire w709;
	wire VRAMA[14];
	wire VRAMA[2];
	wire w712;
	wire w713;
	wire w714;
	wire w715;
	wire w716;
	wire CA[2];
	wire w718;
	wire CA[21];
	wire w720;
	wire w721;
	wire w722;
	wire w723;
	wire w724;
	wire CA[14];
	wire w726;
	wire w727;
	wire VRAMA[15];
	wire CA[15];
	wire VRAMA[1];
	wire w731;
	wire w732;
	wire w733;
	wire w734;
	wire w735;
	wire w736;
	wire w737;
	wire w738;
	wire w739;
	wire w740;
	wire w741;
	wire CA[17];
	wire CA[1];
	wire VRAMA[16];
	wire w745;
	wire w746;
	wire CA[16];
	wire w748;
	wire w749;
	wire w750;
	wire w751;
	wire w752;
	wire w753;
	wire w754;
	wire w755;
	wire w756;
	wire w757;
	wire w758;
	wire w759;
	wire w760;
	wire w761;
	wire w762;
	wire w763;
	wire w764;
	wire w765;
	wire w766;
	wire w767;
	wire w768;
	wire w769;
	wire w770;
	wire w771;
	wire w772;
	wire w773;
	wire w774;
	wire w775;
	wire w776;
	wire w777;
	wire w778;
	wire w779;
	wire w780;
	wire w781;
	wire w782;
	wire w783;
	wire w784;
	wire w785;
	wire w786;
	wire w787;
	wire w788;
	wire w789;
	wire w790;
	wire w791;
	wire w792;
	wire w793;
	wire w794;
	wire w795;
	wire w796;
	wire w797;
	wire w798;
	wire w799;
	wire w800;
	wire w801;
	wire w802;
	wire w803;
	wire w804;
	wire w805;
	wire w806;
	wire w807;
	wire w808;
	wire w809;
	wire w810;
	wire w811;
	wire w812;
	wire w813;
	wire w814;
	wire w815;
	wire w816;
	wire w817;
	wire w818;
	wire w819;
	wire w820;
	wire w821;
	wire w822;
	wire w823;
	wire w824;
	wire w825;
	wire w826;
	wire w827;
	wire w828;
	wire w829;
	wire w830;
	wire w831;
	wire w832;
	wire w833;
	wire w834;
	wire w835;
	wire w836;
	wire w837;
	wire w838;
	wire w839;
	wire w840;
	wire w841;
	wire w842;
	wire w843;
	wire w844;
	wire w845;
	wire w846;
	wire w847;
	wire w848;
	wire w849;
	wire w850;
	wire w851;
	wire w852;
	wire w853;
	wire w854;
	wire w855;
	wire w856;
	wire w857;
	wire w858;
	wire w859;
	wire w860;
	wire w861;
	wire w862;
	wire w863;
	wire w864;
	wire w865;
	wire w866;
	wire w867;
	wire w868;
	wire w869;
	wire w870;
	wire w871;
	wire w872;
	wire w873;
	wire w874;
	wire w875;
	wire w876;
	wire w877;
	wire w878;
	wire w879;
	wire w880;
	wire w881;
	wire w882;
	wire w883;
	wire w884;
	wire w885;
	wire w886;
	wire w887;
	wire w888;
	wire w889;
	wire w890;
	wire w891;
	wire w892;
	wire w893;
	wire w894;
	wire w895;
	wire w896;
	wire w897;
	wire w898;
	wire w899;
	wire w900;
	wire w901;
	wire w902;
	wire w903;
	wire w904;
	wire w905;
	wire w906;
	wire w907;
	wire w908;
	wire w909;
	wire w910;
	wire w911;
	wire w912;
	wire w913;
	wire w914;
	wire w915;
	wire w916;
	wire w917;
	wire w918;
	wire w919;
	wire w920;
	wire w921;
	wire w922;
	wire w923;
	wire w924;
	wire w925;
	wire w926;
	wire w927;
	wire w928;
	wire w929;
	wire w930;
	wire w931;
	wire w932;
	wire w933;
	wire w934;
	wire w935;
	wire w936;
	wire w937;
	wire w938;
	wire w939;
	wire w940;
	wire w941;
	wire w942;
	wire CD[4];
	wire w944;
	wire w945;
	wire w946;
	wire w947;
	wire w948;
	wire w949;
	wire w950;
	wire w951;
	wire w952;
	wire w953;
	wire w954;
	wire w955;
	wire w956;
	wire w957;
	wire w958;
	wire w959;
	wire w960;
	wire w961;
	wire w962;
	wire w963;
	wire w964;
	wire w965;
	wire w966;
	wire w967;
	wire w968;
	wire w969;
	wire w970;
	wire w971;
	wire w972;
	wire w973;
	wire w974;
	wire w975;
	wire w976;
	wire w977;
	wire w978;
	wire w979;
	wire w980;
	wire w981;
	wire w982;
	wire w983;
	wire w984;
	wire w985;
	wire w986;
	wire w987;
	wire w988;
	wire w989;
	wire w990;
	wire w991;
	wire w992;
	wire w993;
	wire FIFO_FULL;
	wire w995;
	wire w996;
	wire w997;
	wire w998;
	wire w999;
	wire w1000;
	wire w1001;
	wire w1002;
	wire w1003;
	wire w1004;
	wire w1005;
	wire w1006;
	wire w1007;
	wire w1008;
	wire w1009;
	wire w1010;
	wire w1011;
	wire w1012;
	wire w1013;
	wire w1014;
	wire PSG_Z80_CLK;
	wire w1016;
	wire w1017;
	wire VPOS[0];
	wire w1019;
	wire w1020;
	wire w1021;
	wire w1022;
	wire w1023;
	wire w1024;
	wire nPSGWRITE;
	wire w1026;
	wire w1027;
	wire w1028;
	wire w1029;
	wire w1030;
	wire w1031;
	wire w1032;
	wire w1033;
	wire w1034;
	wire w1035;
	wire w1036;
	wire w1037;
	wire COL[1];
	wire COL[0];
	wire COL[2];
	wire COL[3];
	wire COL[4];
	wire COL[6];
	wire w1044;
	wire w1045;
	wire w1046;
	wire w1047;
	wire COL[5];
	wire w1049;
	wire w1050;
	wire w1051;
	wire w1052;
	wire w1053;
	wire w1054;
	wire w1055;
	wire w1056;
	wire w1057;
	wire w1058;
	wire w1059;
	wire w1060;
	wire w1061;
	wire DISP;
	wire w1063;
	wire w1064;
	wire w1065;
	wire w1066;
	wire w1067;
	wire w1068;
	wire LSM0;
	wire w1070;
	wire M2;
	wire w1072;
	wire w1073;
	wire w1074;
	wire w1075;
	wire w1076;
	wire w1077;
	wire w1078;
	wire w1079;
	wire w1080;
	wire w1081;
	wire w1082;
	wire LSM1;
	wire w1084;
	wire w1085;
	wire w1086;
	wire w1087;
	wire w1088;
	wire w1089;
	wire w1090;
	wire w1091;
	wire w1092;
	wire w1093;
	wire w1094;
	wire w1095;
	wire w1096;
	wire w1097;
	wire IE2;
	wire IE0;
	wire M1;
	wire w1101;
	wire RS0;
	wire PSG_TEST_OE;
	wire w1104;
	wire w1105;
	wire w1106;
	wire w1107;
	wire w1108;
	wire w1109;
	wire w1110;
	wire w1111;
	wire w1112;
	wire w1113;
	wire PSG_TEST9;
	wire PSG_TEST10;
	wire PSG_TEST11;
	wire w1117;
	wire w1118;
	wire w1119;
	wire w1120;
	wire w1121;
	wire w1122;
	wire w1123;
	wire w1124;
	wire w1125;
	wire w1126;
	wire w1127;
	wire w1128;
	wire w1129;
	wire w1130;
	wire w1131;
	wire w1132;
	wire w1133;
	wire w1134;
	wire w1135;
	wire w1136;
	wire w1137;
	wire w1138;
	wire w1139;
	wire w1140;
	wire w1141;
	wire w1142;
	wire w1143;
	wire w1144;
	wire w1145;
	wire w1146;
	wire w1147;
	wire w1148;
	wire w1149;
	wire w1150;
	wire PAL;
	wire w1152;
	wire w1153;
	wire HIT[0];
	wire w1155;
	wire w1156;
	wire HIT[5];
	wire HIT[6];
	wire HIT[7];
	wire w1160;
	wire w1161;
	wire w1162;
	wire w1163;
	wire HIT[2];
	wire HIT[3];
	wire HIT[4];
	wire w1167;
	wire w1168;
	wire w1169;
	wire HIT[1];
	wire w1171;
	wire w1172;
	wire w1173;
	wire w1174;
	wire w1175;
	wire w1176;
	wire w1177;
	wire w1178;
	wire w1179;
	wire w1180;
	wire w1181;
	wire w1182;
	wire w1183;
	wire w1184;
	wire w1185;
	wire w1186;
	wire w1187;
	wire w1188;
	wire w1189;
	wire w1190;
	wire w1191;
	wire w1192;
	wire w1193;
	wire w1194;
	wire w1195;
	wire w1196;
	wire w1197;
	wire w1198;
	wire w1199;
	wire w1200;
	wire w1201;
	wire w1202;
	wire w1203;
	wire w1204;
	wire w1205;
	wire w1206;
	wire w1207;
	wire w1208;
	wire w1209;
	wire w1210;
	wire w1211;
	wire w1212;
	wire w1213;
	wire w1214;
	wire w1215;
	wire w1216;
	wire w1217;
	wire w1218;
	wire w1219;
	wire w1220;
	wire w1221;
	wire w1222;
	wire w1223;
	wire w1224;
	wire w1225;
	wire w1226;
	wire w1227;
	wire w1228;
	wire w1229;
	wire w1230;
	wire w1231;
	wire w1232;
	wire w1233;
	wire w1234;
	wire w1235;
	wire w1236;
	wire w1237;
	wire w1238;
	wire w1239;
	wire w1240;
	wire w1241;
	wire w1242;
	wire w1243;
	wire w1244;
	wire w1245;
	wire w1246;
	wire w1247;
	wire w1248;
	wire w1249;
	wire w1250;
	wire w1251;
	wire w1252;
	wire w1253;
	wire w1254;
	wire w1255;
	wire w1256;
	wire w1257;
	wire w1258;
	wire w1259;
	wire w1260;
	wire w1261;
	wire w1262;
	wire w1263;
	wire w1264;
	wire w1265;
	wire w1266;
	wire w1267;
	wire w1268;
	wire w1269;
	wire w1270;
	wire w1271;
	wire w1272;
	wire w1273;
	wire w1274;
	wire w1275;
	wire w1276;
	wire w1277;
	wire w1278;
	wire w1279;
	wire w1280;
	wire w1281;
	wire w1282;
	wire w1283;
	wire w1284;
	wire w1285;
	wire w1286;
	wire w1287;
	wire w1288;
	wire w1289;
	wire w1290;
	wire w1291;
	wire w1292;
	wire w1293;
	wire w1294;
	wire w1295;
	wire w1296;
	wire w1297;
	wire w1298;
	wire w1299;
	wire w1300;
	wire w1301;
	wire w1302;
	wire w1303;
	wire w1304;
	wire w1305;
	wire w1306;
	wire w1307;
	wire w1308;
	wire w1309;
	wire w1310;
	wire w1311;
	wire w1312;
	wire w1313;
	wire w1314;
	wire w1315;
	wire w1316;
	wire w1317;
	wire w1318;
	wire w1319;
	wire w1320;
	wire w1321;
	wire w1322;
	wire w1323;
	wire w1324;
	wire w1325;
	wire w1326;
	wire w1327;
	wire w1328;
	wire VRAM_REFRESH;
	wire w1330;
	wire w1331;
	wire w1332;
	wire w1333;
	wire w1334;
	wire w1335;
	wire w1336;
	wire w1337;
	wire w1338;
	wire w1339;
	wire w1340;
	wire w1341;
	wire w1342;
	wire w1343;
	wire w1344;
	wire w1345;
	wire w1346;
	wire w1347;
	wire w1348;
	wire w1349;
	wire w1350;
	wire w1351;
	wire w1352;
	wire w1353;
	wire w1354;
	wire w1355;
	wire w1356;
	wire w1357;
	wire w1358;
	wire w1359;
	wire w1360;
	wire w1361;
	wire w1362;
	wire w1363;
	wire w1364;
	wire w1365;
	wire w1366;
	wire IE1;
	wire w1368;
	wire w1369;
	wire w1370;
	wire w1371;
	wire w1372;
	wire w1373;
	wire w1374;
	wire w1375;
	wire w1376;
	wire w1377;
	wire w1378;
	wire w1379;
	wire w1380;
	wire w1381;
	wire w1382;
	wire w1383;
	wire w1384;
	wire w1385;
	wire w1386;
	wire w1387;
	wire w1388;
	wire w1389;
	wire w1390;
	wire w1391;
	wire w1392;
	wire w1393;
	wire w1394;
	wire w1395;
	wire w1396;
	wire w1397;
	wire w1398;
	wire w1399;
	wire w1400;
	wire w1401;
	wire w1402;
	wire w1403;
	wire w1404;
	wire w1405;
	wire w1406;
	wire w1407;
	wire w1408;
	wire w1409;
	wire w1410;
	wire w1411;
	wire w1412;
	wire w1413;
	wire w1414;
	wire w1415;
	wire w1416;
	wire w1417;
	wire w1418;
	wire w1419;
	wire w1420;
	wire w1421;
	wire w1422;
	wire w1423;
	wire w1424;
	wire w1425;
	wire w1426;
	wire w1427;
	wire w1428;
	wire w1429;
	wire w1430;
	wire w1431;
	wire w1432;
	wire M2;
	wire w1434;
	wire w1435;
	wire w1436;
	wire w1437;
	wire w1438;
	wire w1439;
	wire w1440;
	wire w1441;
	wire w1442;
	wire w1443;
	wire w1444;
	wire w1445;
	wire w1446;
	wire w1447;
	wire CA[18];
	wire w1449;
	wire w1450;
	wire w1451;
	wire w1452;
	wire w1453;
	wire w1454;
	wire w1455;
	wire w1456;
	wire w1457;
	wire w1458;
	wire w1459;
	wire w1460;
	wire w1461;
	wire w1462;
	wire w1463;
	wire w1464;
	wire w1465;
	wire w1466;
	wire w1467;
	wire w1468;
	wire w1469;
	wire w1470;
	wire w1471;
	wire w1472;
	wire w1473;
	wire w1474;
	wire w1475;
	wire w1476;
	wire w1477;
	wire w1478;
	wire w1479;
	wire w1480;
	wire w1481;
	wire w1482;
	wire w1483;
	wire w1484;
	wire w1485;
	wire w1486;
	wire w1487;
	wire w1488;
	wire w1489;
	wire w1490;
	wire w1491;
	wire w1492;
	wire w1493;
	wire w1494;
	wire w1495;
	wire w1496;
	wire w1497;
	wire w1498;
	wire w1499;
	wire w1500;
	wire w1501;
	wire w1502;
	wire w1503;
	wire w1504;
	wire w1505;
	wire w1506;
	wire w1507;
	wire w1508;
	wire w1509;
	wire w1510;
	wire w1511;
	wire w1512;
	wire VPOS[6];
	wire w1514;
	wire w1515;
	wire w1516;
	wire w1517;
	wire w1518;
	wire w1519;
	wire w1520;
	wire w1521;
	wire w1522;
	wire w1523;
	wire w1524;
	wire w1525;
	wire w1526;
	wire w1527;
	wire w1528;
	wire w1529;
	wire w1530;
	wire w1531;
	wire w1532;
	wire w1533;
	wire w1534;
	wire w1535;
	wire w1536;
	wire w1537;
	wire w1538;
	wire w1539;
	wire w1540;
	wire w1541;
	wire w1542;
	wire w1543;
	wire w1544;
	wire w1545;
	wire w1546;
	wire w1547;
	wire w1548;
	wire w1549;
	wire w1550;
	wire w1551;
	wire w1552;
	wire w1553;
	wire w1554;
	wire w1555;
	wire w1556;
	wire w1557;
	wire w1558;
	wire w1559;
	wire w1560;
	wire w1561;
	wire w1562;
	wire w1563;
	wire w1564;
	wire w1565;
	wire w1566;
	wire w1567;
	wire w1568;
	wire w1569;
	wire w1570;
	wire w1571;
	wire w1572;
	wire w1573;
	wire w1574;
	wire w1575;
	wire w1576;
	wire w1577;
	wire w1578;
	wire w1579;
	wire w1580;
	wire w1581;
	wire w1582;
	wire w1583;
	wire w1584;
	wire w1585;
	wire w1586;
	wire w1587;
	wire w1588;
	wire w1589;
	wire w1590;
	wire w1591;
	wire w1592;
	wire w1593;
	wire w1594;
	wire w1595;
	wire VPLA1;
	wire w1597;
	wire w1598;
	wire w1599;
	wire w1600;
	wire w1601;
	wire w1602;
	wire w1603;
	wire w1604;
	wire w1605;
	wire w1606;
	wire HPLA29;
	wire w1608;
	wire w1609;
	wire w1610;
	wire w1611;
	wire w1612;
	wire w1613;
	wire w1614;
	wire w1615;
	wire w1616;
	wire w1617;
	wire w1618;
	wire w1619;
	wire HPLA26;
	wire HPLA24;
	wire HPLA25;
	wire HPLA23;
	wire w1624;
	wire w1625;
	wire w1626;
	wire w1627;
	wire w1628;
	wire w1629;
	wire w1630;
	wire w1631;
	wire w1632;
	wire w1633;
	wire w1634;
	wire w1635;
	wire w1636;
	wire w1637;
	wire w1638;
	wire w1639;
	wire w1640;
	wire w1641;
	wire w1642;
	wire w1643;
	wire w1644;
	wire w1645;
	wire w1646;
	wire w1647;
	wire w1648;
	wire w1649;
	wire w1650;
	wire w1651;
	wire w1652;
	wire w1653;
	wire w1654;
	wire w1655;
	wire w1656;
	wire HPLA30;
	wire w1658;
	wire w1659;
	wire w1660;
	wire w1661;
	wire w1662;
	wire w1663;
	wire w1664;
	wire w1665;
	wire w1666;
	wire w1667;
	wire w1668;
	wire w1669;
	wire w1670;
	wire w1671;
	wire w1672;
	wire w1673;
	wire w1674;
	wire w1675;
	wire w1676;
	wire w1677;
	wire HPLA31;
	wire w1679;
	wire w1680;
	wire HPLA3;
	wire HPLA7;
	wire HPLA6;
	wire w1684;
	wire w1685;
	wire w1686;
	wire w1687;
	wire w1688;
	wire w1689;
	wire w1690;
	wire w1691;
	wire w1692;
	wire w1693;
	wire w1694;
	wire w1695;
	wire HPLA36;
	wire w1697;
	wire HPLA33;
	wire w1699;
	wire w1700;
	wire w1701;
	wire HPLA8;
	wire HPLA18;
	wire HPLA17;
	wire w1705;
	wire w1706;
	wire w1707;
	wire w1708;
	wire w1709;
	wire w1710;
	wire w1711;
	wire w1712;
	wire w1713;
	wire w1714;
	wire w1715;
	wire w1716;
	wire w1717;
	wire w1718;
	wire w1719;
	wire w1720;
	wire w1721;
	wire w1722;
	wire w1723;
	wire w1724;
	wire w1725;
	wire w1726;
	wire w1727;
	wire w1728;
	wire w1729;
	wire w1730;
	wire HPLA35;
	wire w1732;
	wire w1733;
	wire w1734;
	wire w1735;
	wire w1736;
	wire w1737;
	wire w1738;
	wire w1739;
	wire w1740;
	wire w1741;
	wire w1742;
	wire w1743;
	wire w1744;
	wire w1745;
	wire w1746;
	wire w1747;
	wire w1748;
	wire w1749;
	wire w1750;
	wire VPLA0;
	wire VPLA2;
	wire VPLA3;
	wire w1754;
	wire w1755;
	wire w1756;
	wire w1757;
	wire w1758;
	wire w1759;
	wire w1760;
	wire VPLA7;
	wire VPLA6;
	wire VPLA5;
	wire VPLA4;
	wire w1765;
	wire w1766;
	wire w1767;
	wire w1768;
	wire w1769;
	wire w1770;
	wire w1771;
	wire w1772;
	wire w1773;
	wire w1774;
	wire w1775;
	wire w1776;
	wire w1777;
	wire w1778;
	wire w1779;
	wire w1780;
	wire w1781;
	wire w1782;
	wire w1783;
	wire w1784;
	wire w1785;
	wire w1786;
	wire w1787;
	wire w1788;
	wire w1789;
	wire HPLA28;
	wire w1791;
	wire HPLA9;
	wire HPLA20;
	wire HPLA19;
	wire HPLA10;
	wire HPLA16;
	wire HPLA27;
	wire w1798;
	wire w1799;
	wire w1800;
	wire w1801;
	wire w1802;
	wire w1803;
	wire w1804;
	wire w1805;
	wire w1806;
	wire w1807;
	wire w1808;
	wire w1809;
	wire w1810;
	wire w1811;
	wire w1812;
	wire w1813;
	wire w1814;
	wire w1815;
	wire w1816;
	wire w1817;
	wire w1818;
	wire w1819;
	wire w1820;
	wire w1821;
	wire w1822;
	wire w1823;
	wire w1824;
	wire w1825;
	wire w1826;
	wire HPLA22;
	wire HPLA4;
	wire HPLA32;
	wire HPLA2;
	wire HPLA5;
	wire HPLA21;
	wire w1833;
	wire HPLA11;
	wire HPLA14;
	wire HPLA15;
	wire w1837;
	wire HPLA1;
	wire HPLA13;
	wire HPLA12;
	wire w1841;
	wire w1842;
	wire w1843;
	wire w1844;
	wire w1845;
	wire w1846;
	wire w1847;
	wire w1848;
	wire w1849;
	wire w1850;
	wire w1851;
	wire w1852;
	wire w1853;
	wire w1854;
	wire w1855;
	wire w1856;
	wire w1857;
	wire w1858;
	wire HPLA0;
	wire w1860;
	wire HPLA34;
	wire w1862;
	wire w1863;
	wire w1864;
	wire w1865;
	wire w1866;
	wire w1867;
	wire w1868;
	wire w1869;
	wire w1870;
	wire w1871;
	wire w1872;
	wire w1873;
	wire w1874;
	wire w1875;
	wire w1876;
	wire w1877;
	wire w1878;
	wire w1879;
	wire w1880;
	wire w1881;
	wire w1882;
	wire w1883;
	wire w1884;
	wire w1885;
	wire w1886;
	wire w1887;
	wire w1888;
	wire w1889;
	wire w1890;
	wire w1891;
	wire w1892;
	wire w1893;
	wire w1894;
	wire w1895;
	wire w1896;
	wire w1897;
	wire w1898;
	wire w1899;
	wire w1900;
	wire w1901;
	wire w1902;
	wire w1903;
	wire w1904;
	wire w1905;
	wire w1906;
	wire w1907;
	wire w1908;
	wire w1909;
	wire w1910;
	wire w1911;
	wire w1912;
	wire w1913;
	wire w1914;
	wire w1915;
	wire w1916;
	wire w1917;
	wire w1918;
	wire w1919;
	wire w1920;
	wire w1921;
	wire w1922;
	wire w1923;
	wire w1924;
	wire w1925;
	wire w1926;
	wire w1927;
	wire w1928;
	wire w1929;
	wire w1930;
	wire w1931;
	wire w1932;
	wire w1933;
	wire w1934;
	wire w1935;
	wire w1936;
	wire w1937;
	wire w1938;
	wire w1939;
	wire w1940;
	wire w1941;
	wire w1942;
	wire w1943;
	wire w1944;
	wire w1945;
	wire w1946;
	wire w1947;
	wire w1948;
	wire w1949;
	wire w1950;
	wire w1951;
	wire w1952;
	wire w1953;
	wire w1954;
	wire w1955;
	wire w1956;
	wire w1957;
	wire w1958;
	wire w1959;
	wire w1960;
	wire w1961;
	wire w1962;
	wire w1963;
	wire w1964;
	wire w1965;
	wire w1966;
	wire w1967;
	wire w1968;
	wire w1969;
	wire w1970;
	wire w1971;
	wire w1972;
	wire w1973;
	wire w1974;
	wire w1975;
	wire w1976;
	wire w1977;
	wire w1978;
	wire w1979;
	wire w1980;
	wire w1981;
	wire w1982;
	wire w1983;
	wire w1984;
	wire w1985;
	wire w1986;
	wire w1987;
	wire w1988;
	wire w1989;
	wire w1990;
	wire w1991;
	wire w1992;
	wire w1993;
	wire w1994;
	wire w1995;
	wire w1996;
	wire w1997;
	wire w1998;
	wire w1999;
	wire w2000;
	wire w2001;
	wire w2002;
	wire w2003;
	wire w2004;
	wire w2005;
	wire w2006;
	wire w2007;
	wire w2008;
	wire w2009;
	wire w2010;
	wire w2011;
	wire w2012;
	wire w2013;
	wire w2014;
	wire w2015;
	wire w2016;
	wire w2017;
	wire w2018;
	wire w2019;
	wire w2020;
	wire w2021;
	wire w2022;
	wire w2023;
	wire w2024;
	wire w2025;
	wire w2026;
	wire w2027;
	wire w2028;
	wire w2029;
	wire w2030;
	wire w2031;
	wire w2032;
	wire w2033;
	wire w2034;
	wire w2035;
	wire w2036;
	wire w2037;
	wire w2038;
	wire w2039;
	wire w2040;
	wire w2041;
	wire w2042;
	wire w2043;
	wire w2044;
	wire w2045;
	wire w2046;
	wire w2047;
	wire w2048;
	wire w2049;
	wire w2050;
	wire w2051;
	wire w2052;
	wire w2053;
	wire w2054;
	wire w2055;
	wire w2056;
	wire w2057;
	wire w2058;
	wire w2059;
	wire w2060;
	wire w2061;
	wire w2062;
	wire w2063;
	wire w2064;
	wire w2065;
	wire w2066;
	wire w2067;
	wire w2068;
	wire w2069;
	wire w2070;
	wire w2071;
	wire w2072;
	wire w2073;
	wire w2074;
	wire w2075;
	wire w2076;
	wire w2077;
	wire w2078;
	wire w2079;
	wire w2080;
	wire w2081;
	wire w2082;
	wire w2083;
	wire w2084;
	wire w2085;
	wire w2086;
	wire w2087;
	wire w2088;
	wire w2089;
	wire w2090;
	wire w2091;
	wire w2092;
	wire w2093;
	wire w2094;
	wire w2095;
	wire w2096;
	wire w2097;
	wire w2098;
	wire w2099;
	wire w2100;
	wire w2101;
	wire w2102;
	wire w2103;
	wire w2104;
	wire w2105;
	wire w2106;
	wire w2107;
	wire w2108;
	wire w2109;
	wire w2110;
	wire w2111;
	wire w2112;
	wire w2113;
	wire w2114;
	wire w2115;
	wire w2116;
	wire w2117;
	wire w2118;
	wire w2119;
	wire w2120;
	wire w2121;
	wire w2122;
	wire w2123;
	wire PSG_CLK2;
	wire PSG_CLK1;
	wire w2126;
	wire w2127;
	wire w2128;
	wire w2129;
	wire w2130;
	wire w2131;
	wire w2132;
	wire w2133;
	wire PSG_nCLK2;
	wire PSG_nCLK1;
	wire w2136;
	wire w2137;
	wire w2138;
	wire w2139;
	wire w2140;
	wire w2141;
	wire w2142;
	wire w2143;
	wire w2144;
	wire w2145;
	wire w2146;
	wire w2147;
	wire w2148;
	wire w2149;
	wire w2150;
	wire w2151;
	wire w2152;
	wire w2153;
	wire w2154;
	wire w2155;
	wire w2156;
	wire w2157;
	wire w2158;
	wire w2159;
	wire w2160;
	wire w2161;
	wire w2162;
	wire w2163;
	wire w2164;
	wire w2165;
	wire w2166;
	wire w2167;
	wire w2168;
	wire w2169;
	wire w2170;
	wire w2171;
	wire w2172;
	wire w2173;
	wire w2174;
	wire w2175;
	wire w2176;
	wire w2177;
	wire w2178;
	wire w2179;
	wire w2180;
	wire w2181;
	wire w2182;
	wire w2183;
	wire w2184;
	wire w2185;
	wire w2186;
	wire w2187;
	wire w2188;
	wire w2189;
	wire w2190;
	wire w2191;
	wire w2192;
	wire w2193;
	wire w2194;
	wire w2195;
	wire w2196;
	wire w2197;
	wire w2198;
	wire w2199;
	wire w2200;
	wire w2201;
	wire w2202;
	wire w2203;
	wire w2204;
	wire w2205;
	wire w2206;
	wire w2207;
	wire w2208;
	wire w2209;
	wire w2210;
	wire w2211;
	wire w2212;
	wire w2213;
	wire w2214;
	wire w2215;
	wire w2216;
	wire w2217;
	wire w2218;
	wire w2219;
	wire w2220;
	wire w2221;
	wire w2222;
	wire w2223;
	wire w2224;
	wire w2225;
	wire w2226;
	wire w2227;
	wire w2228;
	wire w2229;
	wire w2230;
	wire w2231;
	wire w2232;
	wire w2233;
	wire w2234;
	wire w2235;
	wire w2236;
	wire w2237;
	wire w2238;
	wire w2239;
	wire w2240;
	wire w2241;
	wire w2242;
	wire w2243;
	wire w2244;
	wire w2245;
	wire w2246;
	wire w2247;
	wire w2248;
	wire w2249;
	wire w2250;
	wire w2251;
	wire w2252;
	wire w2253;
	wire w2254;
	wire w2255;
	wire w2256;
	wire w2257;
	wire w2258;
	wire w2259;
	wire w2260;
	wire w2261;
	wire w2262;
	wire w2263;
	wire w2264;
	wire w2265;
	wire w2266;
	wire w2267;
	wire w2268;
	wire w2269;
	wire w2270;
	wire w2271;
	wire w2272;
	wire w2273;
	wire w2274;
	wire w2275;
	wire w2276;
	wire w2277;
	wire w2278;
	wire w2279;
	wire w2280;
	wire w2281;
	wire w2282;
	wire w2283;
	wire w2284;
	wire w2285;
	wire w2286;
	wire w2287;
	wire w2288;
	wire w2289;
	wire w2290;
	wire w2291;
	wire w2292;
	wire w2293;
	wire w2294;
	wire w2295;
	wire w2296;
	wire w2297;
	wire w2298;
	wire w2299;
	wire w2300;
	wire w2301;
	wire w2302;
	wire w2303;
	wire w2304;
	wire w2305;
	wire w2306;
	wire w2307;
	wire w2308;
	wire w2309;
	wire w2310;
	wire w2311;
	wire w2312;
	wire w2313;
	wire w2314;
	wire w2315;
	wire w2316;
	wire w2317;
	wire w2318;
	wire w2319;
	wire w2320;
	wire w2321;
	wire w2322;
	wire w2323;
	wire w2324;
	wire w2325;
	wire w2326;
	wire w2327;
	wire w2328;
	wire w2329;
	wire w2330;
	wire w2331;
	wire w2332;
	wire w2333;
	wire w2334;
	wire w2335;
	wire w2336;
	wire w2337;
	wire w2338;
	wire w2339;
	wire w2340;
	wire w2341;
	wire w2342;
	wire w2343;
	wire w2344;
	wire w2345;
	wire w2346;
	wire w2347;
	wire w2348;
	wire w2349;
	wire w2350;
	wire w2351;
	wire w2352;
	wire w2353;
	wire w2354;
	wire w2355;
	wire w2356;
	wire w2357;
	wire w2358;
	wire w2359;
	wire w2360;
	wire w2361;
	wire w2362;
	wire w2363;
	wire w2364;
	wire w2365;
	wire w2366;
	wire w2367;
	wire w2368;
	wire w2369;
	wire w2370;
	wire w2371;
	wire w2372;
	wire w2373;
	wire w2374;
	wire w2375;
	wire w2376;
	wire w2377;
	wire w2378;
	wire w2379;
	wire w2380;
	wire w2381;
	wire w2382;
	wire w2383;
	wire w2384;
	wire w2385;
	wire w2386;
	wire w2387;
	wire w2388;
	wire w2389;
	wire w2390;
	wire w2391;
	wire w2392;
	wire w2393;
	wire w2394;
	wire w2395;
	wire w2396;
	wire w2397;
	wire w2398;
	wire w2399;
	wire w2400;
	wire w2401;
	wire w2402;
	wire w2403;
	wire w2404;
	wire w2405;
	wire w2406;
	wire w2407;
	wire w2408;
	wire w2409;
	wire w2410;
	wire w2411;
	wire w2412;
	wire w2413;
	wire w2414;
	wire w2415;
	wire w2416;
	wire w2417;
	wire w2418;
	wire w2419;
	wire w2420;
	wire w2421;
	wire w2422;
	wire w2423;
	wire w2424;
	wire w2425;
	wire w2426;
	wire w2427;
	wire w2428;
	wire w2429;
	wire w2430;
	wire w2431;
	wire w2432;
	wire w2433;
	wire w2434;
	wire w2435;
	wire w2436;
	wire w2437;
	wire w2438;
	wire w2439;
	wire w2440;
	wire w2441;
	wire w2442;
	wire w2443;
	wire w2444;
	wire w2445;
	wire w2446;
	wire w2447;
	wire w2448;
	wire w2449;
	wire w2450;
	wire w2451;
	wire w2452;
	wire w2453;
	wire w2454;
	wire w2455;
	wire w2456;
	wire w2457;
	wire w2458;
	wire w2459;
	wire w2460;
	wire w2461;
	wire w2462;
	wire w2463;
	wire w2464;
	wire w2465;
	wire w2466;
	wire w2467;
	wire w2468;
	wire w2469;
	wire w2470;
	wire w2471;
	wire w2472;
	wire w2473;
	wire w2474;
	wire w2475;
	wire w2476;
	wire w2477;
	wire w2478;
	wire w2479;
	wire w2480;
	wire w2481;
	wire w2482;
	wire w2483;
	wire w2484;
	wire w2485;
	wire w2486;
	wire w2487;
	wire w2488;
	wire w2489;
	wire w2490;
	wire w2491;
	wire w2492;
	wire w2493;
	wire w2494;
	wire w2495;
	wire w2496;
	wire w2497;
	wire w2498;
	wire w2499;
	wire w2500;
	wire w2501;
	wire w2502;
	wire w2503;
	wire w2504;
	wire w2505;
	wire w2506;
	wire w2507;
	wire w2508;
	wire w2509;
	wire w2510;
	wire w2511;
	wire w2512;
	wire w2513;
	wire w2514;
	wire w2515;
	wire w2516;
	wire w2517;
	wire w2518;
	wire w2519;
	wire w2520;
	wire w2521;
	wire w2522;
	wire w2523;
	wire w2524;
	wire w2525;
	wire w2526;
	wire w2527;
	wire w2528;
	wire w2529;
	wire w2530;
	wire w2531;
	wire w2532;
	wire w2533;
	wire w2534;
	wire w2535;
	wire w2536;
	wire w2537;
	wire w2538;
	wire w2539;
	wire w2540;
	wire w2541;
	wire w2542;
	wire RES;
	wire w2544;
	wire w2545;
	wire w2546;
	wire w2547;
	wire EDCLK_O;
	wire nYS;
	wire w2550;
	wire w2551;
	wire w2552;
	wire w2553;
	wire w2554;
	wire w2555;
	wire w2556;
	wire w2557;
	wire w2558;
	wire w2559;
	wire w2560;
	wire w2561;
	wire w2562;
	wire w2563;
	wire w2564;
	wire w2565;
	wire w2566;
	wire w2567;
	wire w2568;
	wire w2569;
	wire w2570;
	wire w2571;
	wire w2572;
	wire w2573;
	wire w2574;
	wire w2575;
	wire w2576;
	wire w2577;
	wire w2578;
	wire w2579;
	wire w2580;
	wire w2581;
	wire w2582;
	wire w2583;
	wire w2584;
	wire w2585;
	wire w2586;
	wire w2587;
	wire w2588;
	wire w2589;
	wire w2590;
	wire w2591;
	wire w2592;
	wire w2593;
	wire w2594;
	wire w2595;
	wire w2596;
	wire w2597;
	wire w2598;
	wire w2599;
	wire w2600;
	wire w2601;
	wire w2602;
	wire w2603;
	wire w2604;
	wire w2605;
	wire w2606;
	wire w2607;
	wire SPR_PRIO;
	wire w2609;
	wire w2610;
	wire w2611;
	wire w2612;
	wire w2613;
	wire w2614;
	wire w2615;
	wire w2616;
	wire w2617;
	wire w2618;
	wire w2619;
	wire w2620;
	wire w2621;
	wire w2622;
	wire w2623;
	wire w2624;
	wire w2625;
	wire w2626;
	wire w2627;
	wire w2628;
	wire w2629;
	wire w2630;
	wire w2631;
	wire w2632;
	wire w2633;
	wire w2634;
	wire w2635;
	wire w2636;
	wire w2637;
	wire w2638;
	wire w2639;
	wire w2640;
	wire w2641;
	wire w2642;
	wire w2643;
	wire w2644;
	wire w2645;
	wire w2646;
	wire w2647;
	wire w2648;
	wire w2649;
	wire w2650;
	wire w2651;
	wire w2652;
	wire w2653;
	wire w2654;
	wire w2655;
	wire w2656;
	wire w2657;
	wire w2658;
	wire w2659;
	wire w2660;
	wire w2661;
	wire w2662;
	wire w2663;
	wire w2664;
	wire w2665;
	wire w2666;
	wire w2667;
	wire w2668;
	wire w2669;
	wire w2670;
	wire w2671;
	wire w2672;
	wire w2673;
	wire w2674;
	wire w2675;
	wire w2676;
	wire PLANE_A_PRIO;
	wire PLANE_B_PRIO;
	wire w2679;
	wire w2680;
	wire w2681;
	wire w2682;
	wire w2683;
	wire w2684;
	wire w2685;
	wire w2686;
	wire w2687;
	wire w2688;
	wire w2689;
	wire w2690;
	wire w2691;
	wire w2692;
	wire w2693;
	wire w2694;
	wire w2695;
	wire w2696;
	wire w2697;
	wire w2698;
	wire w2699;
	wire w2700;
	wire w2701;
	wire w2702;
	wire w2703;
	wire w2704;
	wire w2705;
	wire w2706;
	wire w2707;
	wire w2708;
	wire w2709;
	wire w2710;
	wire w2711;
	wire w2712;
	wire w2713;
	wire w2714;
	wire w2715;
	wire w2716;
	wire w2717;
	wire w2718;
	wire w2719;
	wire w2720;
	wire w2721;
	wire w2722;
	wire w2723;
	wire w2724;
	wire w2725;
	wire w2726;
	wire w2727;
	wire w2728;
	wire w2729;
	wire w2730;
	wire w2731;
	wire w2732;
	wire w2733;
	wire w2734;
	wire w2735;
	wire w2736;
	wire w2737;
	wire w2738;
	wire w2739;
	wire w2740;
	wire w2741;
	wire w2742;
	wire w2743;
	wire w2744;
	wire w2745;
	wire w2746;
	wire w2747;
	wire w2748;
	wire w2749;
	wire w2750;
	wire w2751;
	wire w2752;
	wire w2753;
	wire w2754;
	wire w2755;
	wire w2756;
	wire w2757;
	wire w2758;
	wire w2759;
	wire w2760;
	wire w2761;
	wire HIGHLIGHT;
	wire w2763;
	wire w2764;
	wire w2765;
	wire w2766;
	wire w2767;
	wire w2768;
	wire w2769;
	wire w2770;
	wire w2771;
	wire w2772;
	wire w2773;
	wire w2774;
	wire w2775;
	wire w2776;
	wire w2777;
	wire w2778;
	wire w2779;
	wire w2780;
	wire w2781;
	wire w2782;
	wire w2783;
	wire w2784;
	wire SHADOW;
	wire w2786;
	wire w2787;
	wire w2788;
	wire w2789;
	wire w2790;
	wire w2791;
	wire w2792;
	wire w2793;
	wire w2794;
	wire w2795;
	wire w2796;
	wire w2797;
	wire w2798;
	wire w2799;
	wire w2800;
	wire w2801;
	wire w2802;
	wire w2803;
	wire w2804;
	wire w2805;
	wire w2806;
	wire w2807;
	wire w2808;
	wire w2809;
	wire w2810;
	wire w2811;
	wire w2812;
	wire w2813;
	wire w2814;
	wire w2815;
	wire w2816;
	wire w2817;
	wire w2818;
	wire w2819;
	wire w2820;
	wire w2821;
	wire w2822;
	wire w2823;
	wire w2824;
	wire w2825;
	wire w2826;
	wire w2827;
	wire w2828;
	wire w2829;
	wire w2830;
	wire w2831;
	wire w2832;
	wire w2833;
	wire w2834;
	wire w2835;
	wire w2836;
	wire w2837;
	wire w2838;
	wire w2839;
	wire w2840;
	wire w2841;
	wire w2842;
	wire w2843;
	wire w2844;
	wire w2845;
	wire w2846;
	wire w2847;
	wire w2848;
	wire w2849;
	wire w2850;
	wire w2851;
	wire w2852;
	wire w2853;
	wire w2854;
	wire w2855;
	wire w2856;
	wire w2857;
	wire w2858;
	wire w2859;
	wire w2860;
	wire w2861;
	wire w2862;
	wire w2863;
	wire w2864;
	wire w2865;
	wire w2866;
	wire w2867;
	wire w2868;
	wire w2869;
	wire w2870;
	wire w2871;
	wire w2872;
	wire w2873;
	wire w2874;
	wire w2875;
	wire w2876;
	wire w2877;
	wire w2878;
	wire w2879;
	wire w2880;
	wire w2881;
	wire w2882;
	wire w2883;
	wire w2884;
	wire w2885;
	wire w2886;
	wire w2887;
	wire w2888;
	wire w2889;
	wire w2890;
	wire w2891;
	wire w2892;
	wire w2893;
	wire w2894;
	wire w2895;
	wire w2896;
	wire w2897;
	wire w2898;
	wire w2899;
	wire w2900;
	wire w2901;
	wire w2902;
	wire w2903;
	wire w2904;
	wire w2905;
	wire w2906;
	wire w2907;
	wire w2908;
	wire w2909;
	wire w2910;
	wire w2911;
	wire w2912;
	wire w2913;
	wire w2914;
	wire w2915;
	wire w2916;
	wire w2917;
	wire w2918;
	wire w2919;
	wire w2920;
	wire w2921;
	wire w2922;
	wire w2923;
	wire w2924;
	wire w2925;
	wire w2926;
	wire w2927;
	wire w2928;
	wire w2929;
	wire w2930;
	wire w2931;
	wire w2932;
	wire w2933;
	wire w2934;
	wire w2935;
	wire w2936;
	wire w2937;
	wire w2938;
	wire w2939;
	wire w2940;
	wire w2941;
	wire w2942;
	wire w2943;
	wire w2944;
	wire w2945;
	wire w2946;
	wire w2947;
	wire w2948;
	wire w2949;
	wire S[3];
	wire w2951;
	wire w2952;
	wire S[7];
	wire S[2];
	wire w2955;
	wire w2956;
	wire w2957;
	wire w2958;
	wire w2959;
	wire w2960;
	wire S[6];
	wire S[1];
	wire S[5];
	wire S[0];
	wire S[4];
	wire w2966;
	wire w2967;
	wire w2968;
	wire w2969;
	wire w2970;
	wire w2971;
	wire w2972;
	wire w2973;
	wire w2974;
	wire w2975;
	wire w2976;
	wire w2977;
	wire w2978;
	wire w2979;
	wire w2980;
	wire w2981;
	wire w2982;
	wire w2983;
	wire w2984;
	wire w2985;
	wire w2986;
	wire w2987;
	wire w2988;
	wire w2989;
	wire w2990;
	wire w2991;
	wire w2992;
	wire w2993;
	wire w2994;
	wire w2995;
	wire w2996;
	wire w2997;
	wire w2998;
	wire w2999;
	wire w3000;
	wire w3001;
	wire w3002;
	wire w3003;
	wire w3004;
	wire w3005;
	wire w3006;
	wire w3007;
	wire w3008;
	wire w3009;
	wire w3010;
	wire w3011;
	wire w3012;
	wire w3013;
	wire w3014;
	wire w3015;
	wire w3016;
	wire w3017;
	wire w3018;
	wire w3019;
	wire w3020;
	wire w3021;
	wire w3022;
	wire w3023;
	wire w3024;
	wire w3025;
	wire w3026;
	wire w3027;
	wire w3028;
	wire w3029;
	wire w3030;
	wire w3031;
	wire w3032;
	wire w3033;
	wire w3034;
	wire w3035;
	wire w3036;
	wire w3037;
	wire w3038;
	wire w3039;
	wire w3040;
	wire w3041;
	wire w3042;
	wire w3043;
	wire w3044;
	wire w3045;
	wire w3046;
	wire w3047;
	wire w3048;
	wire w3049;
	wire w3050;
	wire w3051;
	wire w3052;
	wire w3053;
	wire w3054;
	wire w3055;
	wire w3056;
	wire w3057;
	wire w3058;
	wire w3059;
	wire w3060;
	wire w3061;
	wire w3062;
	wire w3063;
	wire w3064;
	wire w3065;
	wire w3066;
	wire w3067;
	wire w3068;
	wire w3069;
	wire w3070;
	wire w3071;
	wire w3072;
	wire w3073;
	wire w3074;
	wire w3075;
	wire w3076;
	wire w3077;
	wire w3078;
	wire w3079;
	wire w3080;
	wire w3081;
	wire w3082;
	wire w3083;
	wire w3084;
	wire w3085;
	wire w3086;
	wire w3087;
	wire w3088;
	wire w3089;
	wire w3090;
	wire w3091;
	wire w3092;
	wire w3093;
	wire w3094;
	wire w3095;
	wire w3096;
	wire w3097;
	wire w3098;
	wire w3099;
	wire w3100;
	wire w3101;
	wire w3102;
	wire w3103;
	wire w3104;
	wire w3105;
	wire w3106;
	wire w3107;
	wire w3108;
	wire w3109;
	wire w3110;
	wire w3111;
	wire w3112;
	wire w3113;
	wire w3114;
	wire w3115;
	wire w3116;
	wire w3117;
	wire w3118;
	wire w3119;
	wire w3120;
	wire w3121;
	wire w3122;
	wire w3123;
	wire w3124;
	wire w3125;
	wire w3126;
	wire w3127;
	wire w3128;
	wire w3129;
	wire w3130;
	wire w3131;
	wire w3132;
	wire w3133;
	wire w3134;
	wire w3135;
	wire w3136;
	wire w3137;
	wire w3138;
	wire w3139;
	wire w3140;
	wire w3141;
	wire w3142;
	wire w3143;
	wire w3144;
	wire w3145;
	wire w3146;
	wire w3147;
	wire w3148;
	wire w3149;
	wire w3150;
	wire w3151;
	wire w3152;
	wire w3153;
	wire w3154;
	wire w3155;
	wire w3156;
	wire w3157;
	wire w3158;
	wire w3159;
	wire w3160;
	wire w3161;
	wire w3162;
	wire w3163;
	wire w3164;
	wire w3165;
	wire w3166;
	wire w3167;
	wire w3168;
	wire w3169;
	wire w3170;
	wire w3171;
	wire w3172;
	wire w3173;
	wire w3174;
	wire w3175;
	wire w3176;
	wire w3177;
	wire w3178;
	wire w3179;
	wire w3180;
	wire w3181;
	wire w3182;
	wire w3183;
	wire w3184;
	wire w3185;
	wire w3186;
	wire w3187;
	wire w3188;
	wire w3189;
	wire w3190;
	wire w3191;
	wire w3192;
	wire w3193;
	wire w3194;
	wire w3195;
	wire w3196;
	wire w3197;
	wire w3198;
	wire w3199;
	wire w3200;
	wire w3201;
	wire w3202;
	wire w3203;
	wire w3204;
	wire w3205;
	wire w3206;
	wire w3207;
	wire w3208;
	wire w3209;
	wire w3210;
	wire w3211;
	wire w3212;
	wire w3213;
	wire w3214;
	wire w3215;
	wire w3216;
	wire w3217;
	wire w3218;
	wire w3219;
	wire w3220;
	wire w3221;
	wire w3222;
	wire w3223;
	wire w3224;
	wire w3225;
	wire w3226;
	wire w3227;
	wire w3228;
	wire w3229;
	wire w3230;
	wire w3231;
	wire w3232;
	wire w3233;
	wire w3234;
	wire w3235;
	wire w3236;
	wire w3237;
	wire w3238;
	wire w3239;
	wire w3240;
	wire w3241;
	wire w3242;
	wire w3243;
	wire w3244;
	wire w3245;
	wire w3246;
	wire w3247;
	wire w3248;
	wire w3249;
	wire w3250;
	wire w3251;
	wire w3252;
	wire w3253;
	wire w3254;
	wire w3255;
	wire w3256;
	wire w3257;
	wire w3258;
	wire w3259;
	wire w3260;
	wire w3261;
	wire w3262;
	wire w3263;
	wire w3264;
	wire w3265;
	wire w3266;
	wire w3267;
	wire w3268;
	wire w3269;
	wire w3270;
	wire w3271;
	wire w3272;
	wire w3273;
	wire w3274;
	wire w3275;
	wire w3276;
	wire w3277;
	wire w3278;
	wire w3279;
	wire w3280;
	wire w3281;
	wire w3282;
	wire w3283;
	wire w3284;
	wire w3285;
	wire w3286;
	wire w3287;
	wire w3288;
	wire w3289;
	wire w3290;
	wire w3291;
	wire w3292;
	wire w3293;
	wire w3294;
	wire w3295;
	wire w3296;
	wire w3297;
	wire w3298;
	wire w3299;
	wire w3300;
	wire w3301;
	wire w3302;
	wire w3303;
	wire w3304;
	wire w3305;
	wire w3306;
	wire w3307;
	wire w3308;
	wire w3309;
	wire w3310;
	wire w3311;
	wire w3312;
	wire w3313;
	wire w3314;
	wire w3315;
	wire w3316;
	wire w3317;
	wire w3318;
	wire w3319;
	wire w3320;
	wire w3321;
	wire w3322;
	wire w3323;
	wire w3324;
	wire w3325;
	wire w3326;
	wire w3327;
	wire w3328;
	wire w3329;
	wire w3330;
	wire w3331;
	wire w3332;
	wire w3333;
	wire w3334;
	wire w3335;
	wire w3336;
	wire w3337;
	wire w3338;
	wire w3339;
	wire w3340;
	wire w3341;
	wire w3342;
	wire w3343;
	wire w3344;
	wire w3345;
	wire w3346;
	wire w3347;
	wire w3348;
	wire w3349;
	wire w3350;
	wire w3351;
	wire w3352;
	wire w3353;
	wire w3354;
	wire w3355;
	wire w3356;
	wire w3357;
	wire w3358;
	wire w3359;
	wire w3360;
	wire w3361;
	wire w3362;
	wire w3363;
	wire w3364;
	wire w3365;
	wire w3366;
	wire w3367;
	wire w3368;
	wire w3369;
	wire w3370;
	wire w3371;
	wire w3372;
	wire w3373;
	wire w3374;
	wire w3375;
	wire w3376;
	wire w3377;
	wire w3378;
	wire w3379;
	wire w3380;
	wire w3381;
	wire w3382;
	wire w3383;
	wire w3384;
	wire w3385;
	wire w3386;
	wire w3387;
	wire w3388;
	wire w3389;
	wire w3390;
	wire w3391;
	wire w3392;
	wire w3393;
	wire w3394;
	wire w3395;
	wire w3396;
	wire w3397;
	wire w3398;
	wire w3399;
	wire w3400;
	wire w3401;
	wire w3402;
	wire w3403;
	wire w3404;
	wire w3405;
	wire w3406;
	wire w3407;
	wire w3408;
	wire w3409;
	wire w3410;
	wire w3411;
	wire w3412;
	wire w3413;
	wire w3414;
	wire w3415;
	wire w3416;
	wire w3417;
	wire w3418;
	wire w3419;
	wire w3420;
	wire w3421;
	wire w3422;
	wire w3423;
	wire w3424;
	wire w3425;
	wire w3426;
	wire w3427;
	wire w3428;
	wire w3429;
	wire w3430;
	wire w3431;
	wire w3432;
	wire w3433;
	wire w3434;
	wire w3435;
	wire w3436;
	wire w3437;
	wire w3438;
	wire w3439;
	wire w3440;
	wire w3441;
	wire w3442;
	wire w3443;
	wire w3444;
	wire w3445;
	wire w3446;
	wire w3447;
	wire w3448;
	wire w3449;
	wire w3450;
	wire w3451;
	wire w3452;
	wire w3453;
	wire w3454;
	wire w3455;
	wire w3456;
	wire w3457;
	wire w3458;
	wire w3459;
	wire w3460;
	wire w3461;
	wire w3462;
	wire w3463;
	wire w3464;
	wire w3465;
	wire w3466;
	wire w3467;
	wire w3468;
	wire w3469;
	wire w3470;
	wire w3471;
	wire w3472;
	wire w3473;
	wire w3474;
	wire w3475;
	wire w3476;
	wire w3477;
	wire w3478;
	wire w3479;
	wire w3480;
	wire w3481;
	wire w3482;
	wire w3483;
	wire w3484;
	wire w3485;
	wire w3486;
	wire w3487;
	wire w3488;
	wire w3489;
	wire w3490;
	wire w3491;
	wire w3492;
	wire w3493;
	wire w3494;
	wire w3495;
	wire w3496;
	wire w3497;
	wire w3498;
	wire w3499;
	wire w3500;
	wire w3501;
	wire w3502;
	wire w3503;
	wire w3504;
	wire w3505;
	wire w3506;
	wire w3507;
	wire w3508;
	wire w3509;
	wire w3510;
	wire w3511;
	wire w3512;
	wire w3513;
	wire w3514;
	wire w3515;
	wire w3516;
	wire w3517;
	wire w3518;
	wire w3519;
	wire w3520;
	wire w3521;
	wire w3522;
	wire w3523;
	wire w3524;
	wire w3525;
	wire w3526;
	wire w3527;
	wire w3528;
	wire w3529;
	wire w3530;
	wire w3531;
	wire w3532;
	wire w3533;
	wire w3534;
	wire w3535;
	wire w3536;
	wire w3537;
	wire w3538;
	wire w3539;
	wire w3540;
	wire w3541;
	wire w3542;
	wire w3543;
	wire w3544;
	wire w3545;
	wire w3546;
	wire w3547;
	wire w3548;
	wire w3549;
	wire w3550;
	wire w3551;
	wire w3552;
	wire w3553;
	wire w3554;
	wire w3555;
	wire w3556;
	wire w3557;
	wire w3558;
	wire w3559;
	wire w3560;
	wire w3561;
	wire w3562;
	wire w3563;
	wire w3564;
	wire w3565;
	wire w3566;
	wire w3567;
	wire w3568;
	wire w3569;
	wire w3570;
	wire w3571;
	wire w3572;
	wire w3573;
	wire w3574;
	wire w3575;
	wire w3576;
	wire w3577;
	wire w3578;
	wire w3579;
	wire w3580;
	wire w3581;
	wire w3582;
	wire w3583;
	wire w3584;
	wire w3585;
	wire w3586;
	wire w3587;
	wire w3588;
	wire w3589;
	wire w3590;
	wire w3591;
	wire w3592;
	wire w3593;
	wire w3594;
	wire w3595;
	wire w3596;
	wire w3597;
	wire w3598;
	wire w3599;
	wire w3600;
	wire w3601;
	wire w3602;
	wire w3603;
	wire w3604;
	wire w3605;
	wire w3606;
	wire w3607;
	wire w3608;
	wire w3609;
	wire w3610;
	wire w3611;
	wire w3612;
	wire w3613;
	wire w3614;
	wire w3615;
	wire w3616;
	wire w3617;
	wire w3618;
	wire w3619;
	wire w3620;
	wire w3621;
	wire w3622;
	wire w3623;
	wire w3624;
	wire w3625;
	wire w3626;
	wire w3627;
	wire w3628;
	wire w3629;
	wire w3630;
	wire w3631;
	wire w3632;
	wire w3633;
	wire w3634;
	wire w3635;
	wire w3636;
	wire w3637;
	wire w3638;
	wire w3639;
	wire w3640;
	wire w3641;
	wire w3642;
	wire w3643;
	wire w3644;
	wire w3645;
	wire w3646;
	wire w3647;
	wire w3648;
	wire w3649;
	wire w3650;
	wire w3651;
	wire w3652;
	wire w3653;
	wire w3654;
	wire w3655;
	wire w3656;
	wire w3657;
	wire w3658;
	wire w3659;
	wire w3660;
	wire w3661;
	wire w3662;
	wire w3663;
	wire w3664;
	wire w3665;
	wire w3666;
	wire w3667;
	wire w3668;
	wire w3669;
	wire w3670;
	wire w3671;
	wire w3672;
	wire w3673;
	wire w3674;
	wire w3675;
	wire w3676;
	wire w3677;
	wire w3678;
	wire w3679;
	wire w3680;
	wire w3681;
	wire w3682;
	wire w3683;
	wire w3684;
	wire w3685;
	wire w3686;
	wire w3687;
	wire w3688;
	wire w3689;
	wire w3690;
	wire w3691;
	wire w3692;
	wire w3693;
	wire w3694;
	wire w3695;
	wire w3696;
	wire w3697;
	wire w3698;
	wire w3699;
	wire w3700;
	wire w3701;
	wire w3702;
	wire w3703;
	wire w3704;
	wire w3705;
	wire w3706;
	wire w3707;
	wire w3708;
	wire w3709;
	wire w3710;
	wire w3711;
	wire w3712;
	wire w3713;
	wire w3714;
	wire w3715;
	wire w3716;
	wire w3717;
	wire w3718;
	wire w3719;
	wire w3720;
	wire w3721;
	wire w3722;
	wire w3723;
	wire w3724;
	wire w3725;
	wire w3726;
	wire w3727;
	wire w3728;
	wire w3729;
	wire w3730;
	wire w3731;
	wire w3732;
	wire w3733;
	wire w3734;
	wire w3735;
	wire w3736;
	wire w3737;
	wire w3738;
	wire w3739;
	wire w3740;
	wire w3741;
	wire w3742;
	wire w3743;
	wire w3744;
	wire w3745;
	wire w3746;
	wire w3747;
	wire w3748;
	wire w3749;
	wire w3750;
	wire w3751;
	wire w3752;
	wire w3753;
	wire w3754;
	wire w3755;
	wire w3756;
	wire w3757;
	wire w3758;
	wire w3759;
	wire w3760;
	wire w3761;
	wire w3762;
	wire w3763;
	wire w3764;
	wire w3765;
	wire w3766;
	wire w3767;
	wire w3768;
	wire w3769;
	wire w3770;
	wire w3771;
	wire w3772;
	wire w3773;
	wire w3774;
	wire w3775;
	wire w3776;
	wire w3777;
	wire w3778;
	wire w3779;
	wire w3780;
	wire w3781;
	wire w3782;
	wire w3783;
	wire w3784;
	wire w3785;
	wire w3786;
	wire w3787;
	wire w3788;
	wire w3789;
	wire w3790;
	wire w3791;
	wire w3792;
	wire w3793;
	wire w3794;
	wire w3795;
	wire w3796;
	wire w3797;
	wire w3798;
	wire w3799;
	wire w3800;
	wire w3801;
	wire w3802;
	wire w3803;
	wire w3804;
	wire w3805;
	wire w3806;
	wire w3807;
	wire w3808;
	wire w3809;
	wire w3810;
	wire w3811;
	wire w3812;
	wire w3813;
	wire w3814;
	wire w3815;
	wire w3816;
	wire w3817;
	wire w3818;
	wire w3819;
	wire w3820;
	wire w3821;
	wire w3822;
	wire w3823;
	wire w3824;
	wire w3825;
	wire w3826;
	wire w3827;
	wire w3828;
	wire w3829;
	wire w3830;
	wire w3831;
	wire w3832;
	wire w3833;
	wire w3834;
	wire w3835;
	wire w3836;
	wire w3837;
	wire w3838;
	wire w3839;
	wire w3840;
	wire w3841;
	wire w3842;
	wire w3843;
	wire w3844;
	wire w3845;
	wire w3846;
	wire w3847;
	wire w3848;
	wire w3849;
	wire w3850;
	wire w3851;
	wire w3852;
	wire w3853;
	wire w3854;
	wire w3855;
	wire w3856;
	wire w3857;
	wire w3858;
	wire w3859;
	wire w3860;
	wire w3861;
	wire w3862;
	wire w3863;
	wire w3864;
	wire w3865;
	wire w3866;
	wire w3867;
	wire w3868;
	wire w3869;
	wire w3870;
	wire w3871;
	wire w3872;
	wire w3873;
	wire w3874;
	wire w3875;
	wire w3876;
	wire w3877;
	wire w3878;
	wire w3879;
	wire w3880;
	wire w3881;
	wire w3882;
	wire w3883;
	wire w3884;
	wire w3885;
	wire w3886;
	wire w3887;
	wire w3888;
	wire w3889;
	wire w3890;
	wire w3891;
	wire w3892;
	wire w3893;
	wire w3894;
	wire w3895;
	wire w3896;
	wire w3897;
	wire w3898;
	wire w3899;
	wire w3900;
	wire w3901;
	wire w3902;
	wire w3903;
	wire w3904;
	wire w3905;
	wire w3906;
	wire w3907;
	wire w3908;
	wire w3909;
	wire w3910;
	wire w3911;
	wire w3912;
	wire w3913;
	wire w3914;
	wire w3915;
	wire w3916;
	wire w3917;
	wire w3918;
	wire w3919;
	wire w3920;
	wire w3921;
	wire w3922;
	wire w3923;
	wire w3924;
	wire w3925;
	wire w3926;
	wire w3927;
	wire w3928;
	wire w3929;
	wire w3930;
	wire w3931;
	wire w3932;
	wire w3933;
	wire w3934;
	wire w3935;
	wire w3936;
	wire w3937;
	wire w3938;
	wire w3939;
	wire w3940;
	wire w3941;
	wire w3942;
	wire w3943;
	wire w3944;
	wire w3945;
	wire w3946;
	wire w3947;
	wire w3948;
	wire w3949;
	wire w3950;
	wire w3951;
	wire w3952;
	wire w3953;
	wire w3954;
	wire w3955;
	wire w3956;
	wire w3957;
	wire w3958;
	wire w3959;
	wire w3960;
	wire w3961;
	wire w3962;
	wire w3963;
	wire w3964;
	wire w3965;
	wire w3966;
	wire w3967;
	wire w3968;
	wire w3969;
	wire w3970;
	wire w3971;
	wire w3972;
	wire w3973;
	wire w3974;
	wire w3975;
	wire w3976;
	wire w3977;
	wire w3978;
	wire w3979;
	wire w3980;
	wire w3981;
	wire w3982;
	wire w3983;
	wire w3984;
	wire w3985;
	wire w3986;
	wire w3987;
	wire w3988;
	wire w3989;
	wire w3990;
	wire w3991;
	wire w3992;
	wire w3993;
	wire w3994;
	wire w3995;
	wire w3996;
	wire w3997;
	wire w3998;
	wire w3999;
	wire w4000;
	wire w4001;
	wire w4002;
	wire w4003;
	wire w4004;
	wire w4005;
	wire w4006;
	wire w4007;
	wire w4008;
	wire w4009;
	wire w4010;
	wire w4011;
	wire w4012;
	wire w4013;
	wire w4014;
	wire w4015;
	wire w4016;
	wire w4017;
	wire w4018;
	wire w4019;
	wire w4020;
	wire w4021;
	wire w4022;
	wire w4023;
	wire w4024;
	wire w4025;
	wire w4026;
	wire w4027;
	wire w4028;
	wire w4029;
	wire w4030;
	wire w4031;
	wire w4032;
	wire w4033;
	wire w4034;
	wire w4035;
	wire w4036;
	wire w4037;
	wire w4038;
	wire w4039;
	wire w4040;
	wire w4041;
	wire w4042;
	wire w4043;
	wire w4044;
	wire w4045;
	wire w4046;
	wire w4047;
	wire w4048;
	wire w4049;
	wire w4050;
	wire w4051;
	wire w4052;
	wire w4053;
	wire w4054;
	wire w4055;
	wire w4056;
	wire w4057;
	wire w4058;
	wire w4059;
	wire w4060;
	wire w4061;
	wire w4062;
	wire w4063;
	wire w4064;
	wire w4065;
	wire w4066;
	wire w4067;
	wire w4068;
	wire w4069;
	wire w4070;
	wire w4071;
	wire w4072;
	wire w4073;
	wire w4074;
	wire w4075;
	wire w4076;
	wire w4077;
	wire w4078;
	wire w4079;
	wire w4080;
	wire w4081;
	wire w4082;
	wire w4083;
	wire w4084;
	wire w4085;
	wire w4086;
	wire w4087;
	wire w4088;
	wire w4089;
	wire w4090;
	wire w4091;
	wire w4092;
	wire w4093;
	wire w4094;
	wire w4095;
	wire w4096;
	wire w4097;
	wire w4098;
	wire w4099;
	wire w4100;
	wire w4101;
	wire w4102;
	wire w4103;
	wire w4104;
	wire w4105;
	wire w4106;
	wire w4107;
	wire w4108;
	wire w4109;
	wire w4110;
	wire w4111;
	wire w4112;
	wire w4113;
	wire w4114;
	wire w4115;
	wire w4116;
	wire w4117;
	wire w4118;
	wire w4119;
	wire w4120;
	wire w4121;
	wire w4122;
	wire w4123;
	wire w4124;
	wire w4125;
	wire w4126;
	wire w4127;
	wire w4128;
	wire w4129;
	wire w4130;
	wire w4131;
	wire w4132;
	wire w4133;
	wire w4134;
	wire w4135;
	wire w4136;
	wire w4137;
	wire w4138;
	wire w4139;
	wire w4140;
	wire w4141;
	wire w4142;
	wire w4143;
	wire w4144;
	wire w4145;
	wire w4146;
	wire w4147;
	wire w4148;
	wire w4149;
	wire w4150;
	wire w4151;
	wire w4152;
	wire w4153;
	wire w4154;
	wire w4155;
	wire w4156;
	wire w4157;
	wire w4158;
	wire w4159;
	wire w4160;
	wire w4161;
	wire w4162;
	wire w4163;
	wire w4164;
	wire w4165;
	wire w4166;
	wire w4167;
	wire w4168;
	wire w4169;
	wire w4170;
	wire w4171;
	wire w4172;
	wire w4173;
	wire w4174;
	wire w4175;
	wire w4176;
	wire w4177;
	wire w4178;
	wire w4179;
	wire w4180;
	wire w4181;
	wire w4182;
	wire w4183;
	wire w4184;
	wire w4185;
	wire w4186;
	wire w4187;
	wire w4188;
	wire w4189;
	wire w4190;
	wire w4191;
	wire w4192;
	wire w4193;
	wire w4194;
	wire w4195;
	wire w4196;
	wire w4197;
	wire w4198;
	wire w4199;
	wire w4200;
	wire w4201;
	wire w4202;
	wire w4203;
	wire w4204;
	wire w4205;
	wire w4206;
	wire w4207;
	wire w4208;
	wire w4209;
	wire w4210;
	wire w4211;
	wire w4212;
	wire w4213;
	wire w4214;
	wire w4215;
	wire w4216;
	wire w4217;
	wire w4218;
	wire w4219;
	wire w4220;
	wire w4221;
	wire w4222;
	wire w4223;
	wire w4224;
	wire w4225;
	wire w4226;
	wire w4227;
	wire w4228;
	wire w4229;
	wire w4230;
	wire w4231;
	wire w4232;
	wire w4233;
	wire w4234;
	wire w4235;
	wire w4236;
	wire w4237;
	wire w4238;
	wire w4239;
	wire w4240;
	wire w4241;
	wire w4242;
	wire w4243;
	wire w4244;
	wire w4245;
	wire w4246;
	wire w4247;
	wire w4248;
	wire w4249;
	wire w4250;
	wire w4251;
	wire w4252;
	wire w4253;
	wire w4254;
	wire w4255;
	wire w4256;
	wire w4257;
	wire w4258;
	wire w4259;
	wire w4260;
	wire w4261;
	wire w4262;
	wire w4263;
	wire w4264;
	wire w4265;
	wire w4266;
	wire w4267;
	wire w4268;
	wire w4269;
	wire w4270;
	wire w4271;
	wire w4272;
	wire w4273;
	wire w4274;
	wire w4275;
	wire w4276;
	wire w4277;
	wire w4278;
	wire w4279;
	wire w4280;
	wire w4281;
	wire w4282;
	wire w4283;
	wire w4284;
	wire w4285;
	wire w4286;
	wire w4287;
	wire w4288;
	wire w4289;
	wire w4290;
	wire w4291;
	wire w4292;
	wire w4293;
	wire w4294;
	wire w4295;
	wire w4296;
	wire w4297;
	wire w4298;
	wire w4299;
	wire w4300;
	wire w4301;
	wire w4302;
	wire w4303;
	wire w4304;
	wire w4305;
	wire w4306;
	wire w4307;
	wire w4308;
	wire w4309;
	wire M68K_CPU_CLOCK;
	wire w4311;
	wire w4312;
	wire w4313;
	wire w4314;
	wire w4315;
	wire w4316;
	wire w4317;
	wire w4318;
	wire w4319;
	wire w4320;
	wire w4321;
	wire w4322;
	wire w4323;
	wire w4324;
	wire w4325;
	wire w4326;
	wire w4327;
	wire w4328;
	wire w4329;
	wire w4330;
	wire w4331;
	wire w4332;
	wire w4333;
	wire w4334;
	wire w4335;
	wire w4336;
	wire w4337;
	wire w4338;
	wire w4339;
	wire w4340;
	wire w4341;
	wire w4342;
	wire w4343;
	wire w4344;
	wire w4345;
	wire w4346;
	wire w4347;
	wire w4348;
	wire w4349;
	wire w4350;
	wire w4351;
	wire w4352;
	wire nRAS1;
	wire nCAS1;
	wire nWE1;
	wire nWE0;
	wire nOE1;
	wire AD_RD_DIR;
	wire w4359;
	wire w4360;
	wire w4361;
	wire w4362;
	wire w4363;
	wire w4364;
	wire w4365;
	wire w4366;
	wire w4367;
	wire w4368;
	wire w4369;
	wire w4370;
	wire w4371;
	wire w4372;
	wire w4373;
	wire w4374;
	wire w4375;
	wire w4376;
	wire w4377;
	wire w4378;
	wire w4379;
	wire w4380;
	wire w4381;
	wire w4382;
	wire w4383;
	wire w4384;
	wire w4385;
	wire w4386;
	wire w4387;
	wire w4388;
	wire w4389;
	wire w4390;
	wire w4391;
	wire w4392;
	wire w4393;
	wire w4394;
	wire w4395;
	wire w4396;
	wire w4397;
	wire w4398;
	wire w4399;
	wire w4400;
	wire w4401;
	wire w4402;
	wire w4403;
	wire w4404;
	wire w4405;
	wire w4406;
	wire w4407;
	wire w4408;
	wire w4409;
	wire w4410;
	wire w4411;
	wire w4412;
	wire w4413;
	wire w4414;
	wire w4415;
	wire w4416;
	wire w4417;
	wire w4418;
	wire w4419;
	wire w4420;
	wire w4421;
	wire w4422;
	wire w4423;
	wire w4424;
	wire w4425;
	wire w4426;
	wire w4427;
	wire w4428;
	wire w4429;
	wire w4430;
	wire w4431;
	wire w4432;
	wire w4433;
	wire w4434;
	wire w4435;
	wire w4436;
	wire w4437;
	wire w4438;
	wire w4439;
	wire w4440;
	wire w4441;
	wire w4442;
	wire w4443;
	wire w4444;
	wire w4445;
	wire w4446;
	wire w4447;
	wire w4448;
	wire w4449;
	wire w4450;
	wire w4451;
	wire w4452;
	wire w4453;
	wire w4454;
	wire w4455;
	wire w4456;
	wire w4457;
	wire w4458;
	wire w4459;
	wire w4460;
	wire w4461;
	wire w4462;
	wire w4463;
	wire w4464;
	wire w4465;
	wire w4466;
	wire w4467;
	wire w4468;
	wire w4469;
	wire w4470;
	wire w4471;
	wire w4472;
	wire w4473;
	wire w4474;
	wire w4475;
	wire w4476;
	wire w4477;
	wire w4478;
	wire w4479;
	wire w4480;
	wire w4481;
	wire w4482;
	wire w4483;
	wire w4484;
	wire w4485;
	wire w4486;
	wire w4487;
	wire w4488;
	wire w4489;
	wire w4490;
	wire w4491;
	wire w4492;
	wire w4493;
	wire w4494;
	wire w4495;
	wire w4496;
	wire w4497;
	wire w4498;
	wire w4499;
	wire w4500;
	wire w4501;
	wire w4502;
	wire w4503;
	wire w4504;
	wire w4505;
	wire w4506;
	wire w4507;
	wire w4508;
	wire w4509;
	wire w4510;
	wire w4511;
	wire w4512;
	wire w4513;
	wire w4514;
	wire w4515;
	wire w4516;
	wire w4517;
	wire w4518;
	wire w4519;
	wire w4520;
	wire w4521;
	wire w4522;
	wire w4523;
	wire w4524;
	wire w4525;
	wire w4526;
	wire w4527;
	wire w4528;
	wire w4529;
	wire w4530;
	wire w4531;
	wire w4532;
	wire w4533;
	wire w4534;
	wire w4535;
	wire w4536;
	wire w4537;
	wire w4538;
	wire w4539;
	wire w4540;
	wire w4541;
	wire w4542;
	wire w4543;
	wire w4544;
	wire w4545;
	wire w4546;
	wire w4547;
	wire w4548;
	wire w4549;
	wire w4550;
	wire w4551;
	wire w4552;
	wire w4553;
	wire w4554;
	wire w4555;
	wire w4556;
	wire w4557;
	wire w4558;
	wire w4559;
	wire w4560;
	wire w4561;
	wire w4562;
	wire w4563;
	wire w4564;
	wire w4565;
	wire w4566;
	wire w4567;
	wire w4568;
	wire w4569;
	wire w4570;
	wire w4571;
	wire w4572;
	wire w4573;
	wire w4574;
	wire w4575;
	wire w4576;
	wire w4577;
	wire w4578;
	wire w4579;
	wire w4580;
	wire w4581;
	wire w4582;
	wire w4583;
	wire w4584;
	wire w4585;
	wire w4586;
	wire w4587;
	wire w4588;
	wire w4589;
	wire w4590;
	wire w4591;
	wire w4592;
	wire w4593;
	wire w4594;
	wire w4595;
	wire w4596;
	wire w4597;
	wire w4598;
	wire w4599;
	wire w4600;
	wire w4601;
	wire w4602;
	wire w4603;
	wire w4604;
	wire w4605;
	wire w4606;
	wire w4607;
	wire w4608;
	wire w4609;
	wire w4610;
	wire w4611;
	wire w4612;
	wire w4613;
	wire w4614;
	wire w4615;
	wire w4616;
	wire w4617;
	wire w4618;
	wire w4619;
	wire w4620;
	wire w4621;
	wire w4622;
	wire w4623;
	wire w4624;
	wire w4625;
	wire w4626;
	wire w4627;
	wire w4628;
	wire w4629;
	wire w4630;
	wire w4631;
	wire w4632;
	wire w4633;
	wire w4634;
	wire w4635;
	wire w4636;
	wire w4637;
	wire w4638;
	wire w4639;
	wire w4640;
	wire w4641;
	wire w4642;
	wire w4643;
	wire w4644;
	wire w4645;
	wire w4646;
	wire w4647;
	wire w4648;
	wire w4649;
	wire w4650;
	wire w4651;
	wire w4652;
	wire w4653;
	wire w4654;
	wire w4655;
	wire w4656;
	wire w4657;
	wire w4658;
	wire w4659;
	wire w4660;
	wire w4661;
	wire w4662;
	wire w4663;
	wire w4664;
	wire w4665;
	wire w4666;
	wire w4667;
	wire w4668;
	wire w4669;
	wire w4670;
	wire w4671;
	wire w4672;
	wire w4673;
	wire w4674;
	wire w4675;
	wire w4676;
	wire w4677;
	wire w4678;
	wire w4679;
	wire w4680;
	wire w4681;
	wire w4682;
	wire w4683;
	wire w4684;
	wire w4685;
	wire w4686;
	wire w4687;
	wire w4688;
	wire w4689;
	wire w4690;
	wire w4691;
	wire w4692;
	wire w4693;
	wire w4694;
	wire w4695;
	wire w4696;
	wire w4697;
	wire w4698;
	wire w4699;
	wire w4700;
	wire w4701;
	wire w4702;
	wire w4703;
	wire w4704;
	wire w4705;
	wire w4706;
	wire w4707;
	wire w4708;
	wire w4709;
	wire w4710;
	wire w4711;
	wire w4712;
	wire w4713;
	wire w4714;
	wire w4715;
	wire w4716;
	wire w4717;
	wire w4718;
	wire w4719;
	wire w4720;
	wire w4721;
	wire w4722;
	wire w4723;
	wire w4724;
	wire w4725;
	wire w4726;
	wire w4727;
	wire w4728;
	wire w4729;
	wire w4730;
	wire w4731;
	wire w4732;
	wire w4733;
	wire w4734;
	wire w4735;
	wire w4736;
	wire w4737;
	wire w4738;
	wire w4739;
	wire w4740;
	wire w4741;
	wire w4742;
	wire w4743;
	wire w4744;
	wire w4745;
	wire w4746;
	wire w4747;
	wire w4748;
	wire w4749;
	wire w4750;
	wire w4751;
	wire w4752;
	wire w4753;
	wire w4754;
	wire w4755;
	wire w4756;
	wire w4757;
	wire w4758;
	wire w4759;
	wire w4760;
	wire w4761;
	wire w4762;
	wire w4763;
	wire w4764;
	wire w4765;
	wire w4766;
	wire w4767;
	wire w4768;
	wire w4769;
	wire w4770;
	wire w4771;
	wire w4772;
	wire w4773;
	wire w4774;
	wire w4775;
	wire w4776;
	wire w4777;
	wire w4778;
	wire w4779;
	wire w4780;
	wire w4781;
	wire w4782;
	wire w4783;
	wire w4784;
	wire w4785;
	wire w4786;
	wire w4787;
	wire w4788;
	wire w4789;
	wire w4790;
	wire w4791;
	wire w4792;
	wire w4793;
	wire w4794;
	wire w4795;
	wire w4796;
	wire w4797;
	wire w4798;
	wire w4799;
	wire w4800;
	wire w4801;
	wire w4802;
	wire w4803;
	wire w4804;
	wire w4805;
	wire w4806;
	wire w4807;
	wire w4808;
	wire w4809;
	wire w4810;
	wire w4811;
	wire w4812;
	wire w4813;
	wire w4814;
	wire w4815;
	wire w4816;
	wire w4817;
	wire w4818;
	wire w4819;
	wire w4820;
	wire w4821;
	wire w4822;
	wire w4823;
	wire w4824;
	wire w4825;
	wire w4826;
	wire w4827;
	wire w4828;
	wire w4829;
	wire w4830;
	wire w4831;
	wire w4832;
	wire w4833;
	wire w4834;
	wire w4835;
	wire w4836;
	wire w4837;
	wire w4838;
	wire w4839;
	wire w4840;
	wire w4841;
	wire w4842;
	wire w4843;
	wire w4844;
	wire w4845;
	wire w4846;
	wire w4847;
	wire w4848;
	wire w4849;
	wire w4850;
	wire w4851;
	wire w4852;
	wire w4853;
	wire w4854;
	wire w4855;
	wire w4856;
	wire w4857;
	wire w4858;
	wire w4859;
	wire w4860;
	wire w4861;
	wire w4862;
	wire w4863;
	wire w4864;
	wire w4865;
	wire w4866;
	wire w4867;
	wire w4868;
	wire w4869;
	wire w4870;
	wire w4871;
	wire w4872;
	wire w4873;
	wire w4874;
	wire w4875;
	wire w4876;
	wire w4877;
	wire w4878;
	wire w4879;
	wire w4880;
	wire w4881;
	wire w4882;
	wire w4883;
	wire w4884;
	wire w4885;
	wire w4886;
	wire w4887;
	wire w4888;
	wire w4889;
	wire w4890;
	wire w4891;
	wire w4892;
	wire w4893;
	wire w4894;
	wire w4895;
	wire w4896;
	wire w4897;
	wire w4898;
	wire w4899;
	wire w4900;
	wire w4901;
	wire w4902;
	wire w4903;
	wire w4904;
	wire w4905;
	wire w4906;
	wire w4907;
	wire w4908;
	wire w4909;
	wire w4910;
	wire w4911;
	wire w4912;
	wire w4913;
	wire w4914;
	wire w4915;
	wire w4916;
	wire w4917;
	wire w4918;
	wire w4919;
	wire w4920;
	wire w4921;
	wire w4922;
	wire w4923;
	wire w4924;
	wire w4925;
	wire w4926;
	wire w4927;
	wire w4928;
	wire w4929;
	wire w4930;
	wire w4931;
	wire w4932;
	wire w4933;
	wire w4934;
	wire w4935;
	wire w4936;
	wire w4937;
	wire w4938;
	wire w4939;
	wire w4940;
	wire w4941;
	wire w4942;
	wire w4943;
	wire w4944;
	wire w4945;
	wire w4946;
	wire w4947;
	wire w4948;
	wire w4949;
	wire w4950;
	wire w4951;
	wire w4952;
	wire w4953;
	wire w4954;
	wire w4955;
	wire w4956;
	wire w4957;
	wire w4958;
	wire w4959;
	wire w4960;
	wire w4961;
	wire w4962;
	wire w4963;
	wire w4964;
	wire w4965;
	wire w4966;
	wire w4967;
	wire w4968;
	wire w4969;
	wire w4970;
	wire w4971;
	wire w4972;
	wire w4973;
	wire w4974;
	wire w4975;
	wire w4976;
	wire w4977;
	wire w4978;
	wire w4979;
	wire w4980;
	wire w4981;
	wire w4982;
	wire w4983;
	wire w4984;
	wire w4985;
	wire w4986;
	wire w4987;
	wire w4988;
	wire w4989;
	wire w4990;
	wire w4991;
	wire w4992;
	wire w4993;
	wire w4994;
	wire w4995;
	wire w4996;
	wire w4997;
	wire w4998;
	wire w4999;
	wire w5000;
	wire w5001;
	wire w5002;
	wire w5003;
	wire w5004;
	wire w5005;
	wire w5006;
	wire w5007;
	wire w5008;
	wire w5009;
	wire w5010;
	wire w5011;
	wire w5012;
	wire w5013;
	wire w5014;
	wire w5015;
	wire w5016;
	wire w5017;
	wire w5018;
	wire w5019;
	wire w5020;
	wire w5021;
	wire w5022;
	wire w5023;
	wire w5024;
	wire w5025;
	wire w5026;
	wire w5027;
	wire w5028;
	wire w5029;
	wire w5030;
	wire w5031;
	wire w5032;
	wire w5033;
	wire w5034;
	wire w5035;
	wire w5036;
	wire w5037;
	wire w5038;
	wire w5039;
	wire w5040;
	wire w5041;
	wire w5042;
	wire w5043;
	wire w5044;
	wire w5045;
	wire w5046;
	wire w5047;
	wire w5048;
	wire w5049;
	wire w5050;
	wire w5051;
	wire w5052;
	wire w5053;
	wire w5054;
	wire w5055;
	wire w5056;
	wire w5057;
	wire w5058;
	wire w5059;
	wire w5060;
	wire w5061;
	wire w5062;
	wire w5063;
	wire w5064;
	wire w5065;
	wire w5066;
	wire w5067;
	wire w5068;
	wire w5069;
	wire w5070;
	wire w5071;
	wire w5072;
	wire w5073;
	wire w5074;
	wire w5075;
	wire w5076;
	wire w5077;
	wire w5078;
	wire w5079;
	wire w5080;
	wire w5081;
	wire w5082;
	wire w5083;
	wire w5084;
	wire w5085;
	wire w5086;
	wire w5087;
	wire w5088;
	wire w5089;
	wire w5090;
	wire w5091;
	wire w5092;
	wire w5093;
	wire w5094;
	wire w5095;
	wire w5096;
	wire w5097;
	wire w5098;
	wire w5099;
	wire w5100;
	wire w5101;
	wire w5102;
	wire w5103;
	wire w5104;
	wire w5105;
	wire w5106;
	wire w5107;
	wire w5108;
	wire w5109;
	wire w5110;
	wire w5111;
	wire w5112;
	wire w5113;
	wire w5114;
	wire w5115;
	wire w5116;
	wire w5117;
	wire w5118;
	wire w5119;
	wire w5120;
	wire w5121;
	wire w5122;
	wire w5123;
	wire w5124;
	wire w5125;
	wire w5126;
	wire w5127;
	wire w5128;
	wire w5129;
	wire w5130;
	wire w5131;
	wire w5132;
	wire w5133;
	wire w5134;
	wire w5135;
	wire w5136;
	wire w5137;
	wire w5138;
	wire w5139;
	wire w5140;
	wire w5141;
	wire w5142;
	wire w5143;
	wire w5144;
	wire w5145;
	wire w5146;
	wire w5147;
	wire w5148;
	wire w5149;
	wire w5150;
	wire w5151;
	wire w5152;
	wire w5153;
	wire w5154;
	wire w5155;
	wire w5156;
	wire w5157;
	wire w5158;
	wire w5159;
	wire w5160;
	wire w5161;
	wire w5162;
	wire w5163;
	wire nSRLOAD;
	wire w5165;
	wire w5166;
	wire w5167;
	wire w5168;
	wire w5169;
	wire w5170;
	wire w5171;
	wire w5172;
	wire w5173;
	wire w5174;
	wire w5175;
	wire w5176;
	wire w5177;
	wire w5178;
	wire w5179;
	wire w5180;
	wire w5181;
	wire w5182;
	wire w5183;
	wire w5184;
	wire w5185;
	wire w5186;
	wire w5187;
	wire w5188;
	wire w5189;
	wire w5190;
	wire w5191;
	wire w5192;
	wire w5193;
	wire w5194;
	wire w5195;
	wire w5196;
	wire w5197;
	wire w5198;
	wire w5199;
	wire w5200;
	wire w5201;
	wire w5202;
	wire w5203;
	wire w5204;
	wire w5205;
	wire w5206;
	wire w5207;
	wire w5208;
	wire w5209;
	wire w5210;
	wire w5211;
	wire w5212;
	wire w5213;
	wire w5214;
	wire w5215;
	wire w5216;
	wire w5217;
	wire w5218;
	wire w5219;
	wire w5220;
	wire w5221;
	wire w5222;
	wire w5223;
	wire w5224;
	wire w5225;
	wire w5226;
	wire w5227;
	wire w5228;
	wire w5229;
	wire w5230;
	wire w5231;
	wire w5232;
	wire w5233;
	wire w5234;
	wire w5235;
	wire w5236;
	wire w5237;
	wire w5238;
	wire w5239;
	wire w5240;
	wire w5241;
	wire w5242;
	wire w5243;
	wire w5244;
	wire w5245;
	wire w5246;
	wire w5247;
	wire w5248;
	wire w5249;
	wire w5250;
	wire w5251;
	wire w5252;
	wire w5253;
	wire w5254;
	wire w5255;
	wire w5256;
	wire w5257;
	wire w5258;
	wire w5259;
	wire w5260;
	wire w5261;
	wire w5262;
	wire w5263;
	wire w5264;
	wire w5265;
	wire w5266;
	wire w5267;
	wire w5268;
	wire w5269;
	wire w5270;
	wire w5271;
	wire w5272;
	wire w5273;
	wire w5274;
	wire w5275;
	wire w5276;
	wire w5277;
	wire w5278;
	wire w5279;
	wire w5280;
	wire w5281;
	wire w5282;
	wire w5283;
	wire w5284;
	wire w5285;
	wire w5286;
	wire w5287;
	wire w5288;
	wire w5289;
	wire w5290;
	wire w5291;
	wire w5292;
	wire w5293;
	wire w5294;
	wire w5295;
	wire w5296;
	wire w5297;
	wire w5298;
	wire w5299;
	wire w5300;
	wire w5301;
	wire w5302;
	wire w5303;
	wire w5304;
	wire w5305;
	wire w5306;
	wire w5307;
	wire w5308;
	wire w5309;
	wire w5310;
	wire w5311;
	wire w5312;
	wire w5313;
	wire w5314;
	wire w5315;
	wire w5316;
	wire w5317;
	wire w5318;
	wire w5319;
	wire w5320;
	wire w5321;
	wire w5322;
	wire w5323;
	wire w5324;
	wire w5325;
	wire w5326;
	wire w5327;
	wire w5328;
	wire w5329;
	wire w5330;
	wire w5331;
	wire w5332;
	wire w5333;
	wire w5334;
	wire w5335;
	wire w5336;
	wire w5337;
	wire w5338;
	wire w5339;
	wire w5340;
	wire w5341;
	wire w5342;
	wire w5343;
	wire w5344;
	wire w5345;
	wire w5346;
	wire w5347;
	wire w5348;
	wire w5349;
	wire w5350;
	wire w5351;
	wire w5352;
	wire w5353;
	wire w5354;
	wire w5355;
	wire w5356;
	wire w5357;
	wire w5358;
	wire w5359;
	wire w5360;
	wire w5361;
	wire w5362;
	wire w5363;
	wire w5364;
	wire w5365;
	wire w5366;
	wire w5367;
	wire w5368;
	wire w5369;
	wire w5370;
	wire w5371;
	wire w5372;
	wire w5373;
	wire w5374;
	wire w5375;
	wire w5376;
	wire w5377;
	wire w5378;
	wire w5379;
	wire w5380;
	wire w5381;
	wire w5382;
	wire w5383;
	wire w5384;
	wire w5385;
	wire w5386;
	wire w5387;
	wire w5388;
	wire w5389;
	wire w5390;
	wire w5391;
	wire w5392;
	wire w5393;
	wire w5394;
	wire w5395;
	wire w5396;
	wire w5397;
	wire w5398;
	wire w5399;
	wire w5400;
	wire w5401;
	wire w5402;
	wire w5403;
	wire w5404;
	wire w5405;
	wire w5406;
	wire w5407;
	wire w5408;
	wire w5409;
	wire w5410;
	wire w5411;
	wire w5412;
	wire w5413;
	wire w5414;
	wire w5415;
	wire w5416;
	wire w5417;
	wire w5418;
	wire w5419;
	wire w5420;
	wire w5421;
	wire w5422;
	wire w5423;
	wire w5424;
	wire w5425;
	wire w5426;
	wire w5427;
	wire w5428;
	wire w5429;
	wire w5430;
	wire w5431;
	wire w5432;
	wire w5433;
	wire w5434;
	wire w5435;
	wire w5436;
	wire w5437;
	wire w5438;
	wire w5439;
	wire w5440;
	wire w5441;
	wire w5442;
	wire w5443;
	wire w5444;
	wire w5445;
	wire w5446;
	wire w5447;
	wire w5448;
	wire w5449;
	wire w5450;
	wire w5451;
	wire w5452;
	wire w5453;
	wire w5454;
	wire w5455;
	wire w5456;
	wire w5457;
	wire w5458;
	wire w5459;
	wire w5460;
	wire w5461;
	wire w5462;
	wire w5463;
	wire w5464;
	wire w5465;
	wire w5466;
	wire w5467;
	wire w5468;
	wire w5469;
	wire w5470;
	wire w5471;
	wire w5472;
	wire w5473;
	wire w5474;
	wire w5475;
	wire w5476;
	wire w5477;
	wire w5478;
	wire w5479;
	wire w5480;
	wire w5481;
	wire w5482;
	wire w5483;
	wire w5484;
	wire w5485;
	wire w5486;
	wire w5487;
	wire w5488;
	wire w5489;
	wire w5490;
	wire w5491;
	wire w5492;
	wire w5493;
	wire w5494;
	wire w5495;
	wire w5496;
	wire w5497;
	wire w5498;
	wire w5499;
	wire w5500;
	wire w5501;
	wire w5502;
	wire w5503;
	wire w5504;
	wire w5505;
	wire w5506;
	wire w5507;
	wire w5508;
	wire w5509;
	wire w5510;
	wire w5511;
	wire w5512;
	wire w5513;
	wire w5514;
	wire w5515;
	wire w5516;
	wire w5517;
	wire w5518;
	wire w5519;
	wire w5520;
	wire w5521;
	wire w5522;
	wire w5523;
	wire w5524;
	wire w5525;
	wire w5526;
	wire w5527;
	wire w5528;
	wire w5529;
	wire w5530;
	wire w5531;
	wire w5532;
	wire w5533;
	wire w5534;
	wire w5535;
	wire w5536;
	wire w5537;
	wire w5538;
	wire w5539;
	wire w5540;
	wire w5541;
	wire w5542;
	wire w5543;
	wire w5544;
	wire w5545;
	wire w5546;
	wire w5547;
	wire w5548;
	wire w5549;
	wire w5550;
	wire w5551;
	wire w5552;
	wire w5553;
	wire w5554;
	wire w5555;
	wire w5556;
	wire w5557;
	wire w5558;
	wire w5559;
	wire w5560;
	wire w5561;
	wire w5562;
	wire w5563;
	wire w5564;
	wire w5565;
	wire w5566;
	wire w5567;
	wire w5568;
	wire w5569;
	wire w5570;
	wire w5571;
	wire w5572;
	wire w5573;
	wire w5574;
	wire w5575;
	wire w5576;
	wire w5577;
	wire w5578;
	wire w5579;
	wire w5580;
	wire w5581;
	wire w5582;
	wire w5583;
	wire w5584;
	wire w5585;
	wire w5586;
	wire w5587;
	wire w5588;
	wire w5589;
	wire w5590;
	wire w5591;
	wire w5592;
	wire w5593;
	wire w5594;
	wire w5595;
	wire w5596;
	wire w5597;
	wire w5598;
	wire w5599;
	wire w5600;
	wire w5601;
	wire w5602;
	wire w5603;
	wire w5604;
	wire w5605;
	wire w5606;
	wire w5607;
	wire w5608;
	wire w5609;
	wire w5610;
	wire w5611;
	wire w5612;
	wire w5613;
	wire w5614;
	wire w5615;
	wire w5616;
	wire w5617;
	wire w5618;
	wire w5619;
	wire w5620;
	wire w5621;
	wire w5622;
	wire w5623;
	wire w5624;
	wire w5625;
	wire w5626;
	wire w5627;
	wire w5628;
	wire w5629;
	wire w5630;
	wire w5631;
	wire w5632;
	wire w5633;
	wire w5634;
	wire w5635;
	wire w5636;
	wire w5637;
	wire w5638;
	wire w5639;
	wire w5640;
	wire w5641;
	wire w5642;
	wire w5643;
	wire w5644;
	wire w5645;
	wire w5646;
	wire w5647;
	wire w5648;
	wire w5649;
	wire w5650;
	wire w5651;
	wire w5652;
	wire w5653;
	wire w5654;
	wire w5655;
	wire w5656;
	wire w5657;
	wire w5658;
	wire w5659;
	wire w5660;
	wire w5661;
	wire w5662;
	wire w5663;
	wire w5664;
	wire w5665;
	wire w5666;
	wire w5667;
	wire w5668;
	wire w5669;
	wire w5670;
	wire w5671;
	wire w5672;
	wire w5673;
	wire w5674;
	wire w5675;
	wire w5676;
	wire w5677;
	wire w5678;
	wire w5679;
	wire w5680;
	wire w5681;
	wire w5682;
	wire w5683;
	wire w5684;
	wire w5685;
	wire w5686;
	wire w5687;
	wire w5688;
	wire w5689;
	wire w5690;
	wire w5691;
	wire w5692;
	wire w5693;
	wire w5694;
	wire w5695;
	wire w5696;
	wire w5697;
	wire w5698;
	wire w5699;
	wire w5700;
	wire w5701;
	wire w5702;
	wire w5703;
	wire w5704;
	wire w5705;
	wire w5706;
	wire w5707;
	wire w5708;
	wire w5709;
	wire w5710;
	wire w5711;
	wire w5712;
	wire w5713;
	wire w5714;
	wire w5715;
	wire w5716;
	wire w5717;
	wire w5718;
	wire w5719;
	wire w5720;
	wire w5721;
	wire w5722;
	wire w5723;
	wire w5724;
	wire w5725;
	wire w5726;
	wire w5727;
	wire w5728;
	wire w5729;
	wire w5730;
	wire w5731;
	wire w5732;
	wire w5733;
	wire w5734;
	wire w5735;
	wire w5736;
	wire w5737;
	wire w5738;
	wire w5739;
	wire w5740;
	wire w5741;
	wire w5742;
	wire w5743;
	wire w5744;
	wire w5745;
	wire w5746;
	wire w5747;
	wire w5748;
	wire w5749;
	wire w5750;
	wire w5751;
	wire w5752;
	wire w5753;
	wire w5754;
	wire w5755;
	wire w5756;
	wire w5757;
	wire w5758;
	wire w5759;
	wire w5760;
	wire w5761;
	wire w5762;
	wire w5763;
	wire w5764;
	wire w5765;
	wire w5766;
	wire w5767;
	wire w5768;
	wire w5769;
	wire w5770;
	wire w5771;
	wire w5772;
	wire w5773;
	wire w5774;
	wire w5775;
	wire w5776;
	wire w5777;
	wire w5778;
	wire w5779;
	wire w5780;
	wire w5781;
	wire w5782;
	wire w5783;
	wire w5784;
	wire w5785;
	wire w5786;
	wire w5787;
	wire w5788;
	wire w5789;
	wire w5790;
	wire w5791;
	wire w5792;
	wire w5793;
	wire w5794;
	wire w5795;
	wire w5796;
	wire w5797;
	wire w5798;
	wire w5799;
	wire w5800;
	wire w5801;
	wire w5802;
	wire w5803;
	wire w5804;
	wire w5805;
	wire w5806;
	wire w5807;
	wire w5808;
	wire w5809;
	wire w5810;
	wire w5811;
	wire w5812;
	wire w5813;
	wire w5814;
	wire w5815;
	wire w5816;
	wire w5817;
	wire w5818;
	wire w5819;
	wire w5820;
	wire w5821;
	wire w5822;
	wire w5823;
	wire w5824;
	wire w5825;
	wire w5826;
	wire w5827;
	wire w5828;
	wire w5829;
	wire w5830;
	wire w5831;
	wire w5832;
	wire w5833;
	wire w5834;
	wire w5835;
	wire w5836;
	wire w5837;
	wire w5838;
	wire w5839;
	wire w5840;
	wire w5841;
	wire w5842;
	wire w5843;
	wire w5844;
	wire w5845;
	wire w5846;
	wire w5847;
	wire w5848;
	wire w5849;
	wire w5850;
	wire w5851;
	wire w5852;
	wire w5853;
	wire w5854;
	wire w5855;
	wire w5856;
	wire w5857;
	wire w5858;
	wire w5859;
	wire w5860;
	wire w5861;
	wire w5862;
	wire w5863;
	wire w5864;
	wire w5865;
	wire w5866;
	wire w5867;
	wire w5868;
	wire w5869;
	wire w5870;
	wire w5871;
	wire w5872;
	wire w5873;
	wire w5874;
	wire w5875;
	wire w5876;
	wire w5877;
	wire w5878;
	wire w5879;
	wire w5880;
	wire w5881;
	wire w5882;
	wire w5883;
	wire w5884;
	wire w5885;
	wire w5886;
	wire w5887;
	wire w5888;
	wire w5889;
	wire w5890;
	wire w5891;
	wire w5892;
	wire w5893;
	wire w5894;
	wire w5895;
	wire w5896;
	wire w5897;
	wire w5898;
	wire w5899;
	wire w5900;
	wire w5901;
	wire w5902;
	wire w5903;
	wire w5904;
	wire w5905;
	wire w5906;
	wire w5907;
	wire w5908;
	wire w5909;
	wire w5910;
	wire w5911;
	wire w5912;
	wire w5913;
	wire w5914;
	wire w5915;
	wire w5916;
	wire w5917;
	wire w5918;
	wire w5919;
	wire w5920;
	wire w5921;
	wire w5922;
	wire w5923;
	wire w5924;
	wire w5925;
	wire w5926;
	wire w5927;
	wire w5928;
	wire w5929;
	wire w5930;
	wire w5931;
	wire w5932;
	wire w5933;
	wire w5934;
	wire w5935;
	wire w5936;
	wire w5937;
	wire w5938;
	wire w5939;
	wire w5940;
	wire w5941;
	wire w5942;
	wire w5943;
	wire w5944;
	wire w5945;
	wire w5946;
	wire w5947;
	wire w5948;
	wire w5949;
	wire w5950;
	wire w5951;
	wire w5952;
	wire w5953;
	wire w5954;
	wire w5955;
	wire w5956;
	wire w5957;
	wire w5958;
	wire w5959;
	wire w5960;
	wire w5961;
	wire w5962;
	wire w5963;
	wire w5964;
	wire w5965;
	wire w5966;
	wire w5967;
	wire w5968;
	wire w5969;
	wire w5970;
	wire w5971;
	wire w5972;
	wire w5973;
	wire w5974;
	wire w5975;
	wire w5976;
	wire w5977;
	wire w5978;
	wire w5979;
	wire w5980;
	wire w5981;
	wire w5982;
	wire w5983;
	wire w5984;
	wire w5985;
	wire w5986;
	wire w5987;
	wire w5988;
	wire w5989;
	wire w5990;
	wire w5991;
	wire w5992;
	wire w5993;
	wire w5994;
	wire w5995;
	wire w5996;
	wire w5997;
	wire w5998;
	wire w5999;
	wire w6000;
	wire w6001;
	wire w6002;
	wire w6003;
	wire w6004;
	wire w6005;
	wire w6006;
	wire w6007;
	wire w6008;
	wire w6009;
	wire w6010;
	wire w6011;
	wire w6012;
	wire w6013;
	wire w6014;
	wire w6015;
	wire w6016;
	wire w6017;
	wire w6018;
	wire w6019;
	wire w6020;
	wire w6021;
	wire w6022;
	wire w6023;
	wire w6024;
	wire w6025;
	wire w6026;
	wire w6027;
	wire w6028;
	wire w6029;
	wire w6030;
	wire w6031;
	wire w6032;
	wire w6033;
	wire w6034;
	wire w6035;
	wire w6036;
	wire w6037;
	wire w6038;
	wire w6039;
	wire w6040;
	wire w6041;
	wire w6042;
	wire w6043;
	wire w6044;
	wire w6045;
	wire w6046;
	wire w6047;
	wire w6048;
	wire w6049;
	wire w6050;
	wire w6051;
	wire w6052;
	wire w6053;
	wire w6054;
	wire w6055;
	wire w6056;
	wire w6057;
	wire w6058;
	wire w6059;
	wire w6060;
	wire w6061;
	wire w6062;
	wire w6063;
	wire w6064;
	wire w6065;
	wire w6066;
	wire w6067;
	wire w6068;
	wire w6069;
	wire w6070;
	wire w6071;
	wire w6072;
	wire w6073;
	wire w6074;
	wire w6075;
	wire w6076;
	wire w6077;
	wire w6078;
	wire w6079;
	wire w6080;
	wire w6081;
	wire w6082;
	wire w6083;
	wire w6084;
	wire w6085;
	wire w6086;
	wire w6087;
	wire w6088;
	wire w6089;
	wire w6090;
	wire w6091;
	wire w6092;
	wire w6093;
	wire w6094;
	wire w6095;
	wire w6096;
	wire w6097;
	wire w6098;
	wire w6099;
	wire w6100;
	wire w6101;
	wire w6102;
	wire w6103;
	wire w6104;
	wire w6105;
	wire w6106;
	wire w6107;
	wire w6108;
	wire w6109;
	wire w6110;
	wire w6111;
	wire w6112;
	wire w6113;
	wire w6114;
	wire w6115;
	wire w6116;
	wire w6117;
	wire w6118;
	wire w6119;
	wire w6120;
	wire w6121;
	wire w6122;
	wire w6123;
	wire w6124;
	wire w6125;
	wire w6126;
	wire w6127;
	wire w6128;
	wire w6129;
	wire w6130;
	wire w6131;
	wire w6132;
	wire w6133;
	wire w6134;
	wire w6135;
	wire w6136;
	wire w6137;
	wire w6138;
	wire w6139;
	wire w6140;
	wire w6141;
	wire w6142;
	wire w6143;
	wire w6144;
	wire w6145;
	wire w6146;
	wire w6147;
	wire w6148;
	wire w6149;
	wire w6150;
	wire w6151;
	wire w6152;
	wire w6153;
	wire w6154;
	wire w6155;
	wire w6156;
	wire w6157;
	wire w6158;
	wire w6159;
	wire w6160;
	wire w6161;
	wire w6162;
	wire w6163;
	wire w6164;
	wire w6165;
	wire w6166;
	wire w6167;
	wire w6168;
	wire w6169;
	wire w6170;
	wire w6171;
	wire w6172;
	wire w6173;
	wire w6174;
	wire w6175;
	wire w6176;
	wire w6177;
	wire w6178;
	wire w6179;
	wire w6180;
	wire w6181;
	wire w6182;
	wire w6183;
	wire w6184;
	wire w6185;
	wire w6186;
	wire w6187;
	wire w6188;
	wire w6189;
	wire w6190;
	wire w6191;
	wire w6192;
	wire w6193;
	wire w6194;
	wire w6195;
	wire w6196;
	wire w6197;
	wire w6198;
	wire w6199;
	wire w6200;
	wire w6201;
	wire w6202;
	wire w6203;
	wire w6204;
	wire w6205;
	wire w6206;
	wire w6207;
	wire w6208;
	wire w6209;
	wire w6210;
	wire w6211;
	wire w6212;
	wire w6213;
	wire w6214;
	wire w6215;
	wire w6216;
	wire w6217;
	wire w6218;
	wire w6219;
	wire w6220;
	wire w6221;
	wire w6222;
	wire w6223;
	wire w6224;
	wire w6225;
	wire w6226;
	wire w6227;
	wire w6228;
	wire w6229;
	wire w6230;
	wire w6231;
	wire w6232;
	wire w6233;
	wire w6234;
	wire w6235;
	wire w6236;
	wire w6237;
	wire w6238;
	wire w6239;
	wire w6240;
	wire w6241;
	wire w6242;
	wire w6243;
	wire w6244;
	wire w6245;
	wire w6246;
	wire w6247;
	wire w6248;
	wire w6249;
	wire w6250;
	wire w6251;
	wire w6252;
	wire w6253;
	wire w6254;
	wire w6255;
	wire w6256;
	wire w6257;
	wire w6258;
	wire w6259;
	wire w6260;
	wire w6261;
	wire w6262;
	wire w6263;
	wire w6264;
	wire w6265;
	wire w6266;
	wire w6267;
	wire w6268;
	wire w6269;
	wire w6270;
	wire w6271;
	wire w6272;
	wire w6273;
	wire w6274;
	wire w6275;
	wire w6276;
	wire w6277;
	wire w6278;
	wire w6279;
	wire w6280;
	wire w6281;
	wire w6282;
	wire w6283;
	wire w6284;
	wire w6285;
	wire w6286;
	wire w6287;
	wire w6288;
	wire w6289;
	wire w6290;
	wire w6291;
	wire w6292;
	wire w6293;
	wire w6294;
	wire w6295;
	wire w6296;
	wire w6297;
	wire w6298;
	wire w6299;
	wire w6300;
	wire w6301;
	wire w6302;
	wire w6303;
	wire w6304;
	wire w6305;
	wire w6306;
	wire w6307;
	wire w6308;
	wire w6309;
	wire w6310;
	wire w6311;
	wire w6312;
	wire w6313;
	wire w6314;
	wire w6315;
	wire w6316;
	wire w6317;
	wire w6318;
	wire w6319;
	wire w6320;
	wire w6321;
	wire w6322;
	wire w6323;
	wire w6324;
	wire w6325;
	wire w6326;
	wire w6327;
	wire w6328;
	wire w6329;
	wire w6330;
	wire w6331;
	wire w6332;
	wire w6333;
	wire w6334;
	wire w6335;
	wire w6336;
	wire w6337;
	wire w6338;
	wire w6339;
	wire w6340;
	wire w6341;
	wire w6342;
	wire w6343;
	wire w6344;
	wire w6345;
	wire w6346;
	wire w6347;
	wire w6348;
	wire w6349;
	wire w6350;
	wire w6351;
	wire w6352;
	wire w6353;
	wire w6354;
	wire w6355;
	wire w6356;
	wire w6357;
	wire w6358;
	wire w6359;
	wire w6360;
	wire w6361;
	wire w6362;
	wire w6363;
	wire w6364;
	wire w6365;
	wire w6366;
	wire w6367;
	wire w6368;
	wire w6369;
	wire w6370;
	wire w6371;
	wire w6372;
	wire w6373;
	wire w6374;
	wire w6375;
	wire w6376;
	wire w6377;
	wire w6378;
	wire w6379;
	wire w6380;
	wire w6381;
	wire w6382;
	wire w6383;
	wire w6384;
	wire w6385;
	wire w6386;
	wire w6387;
	wire w6388;
	wire w6389;
	wire w6390;
	wire w6391;
	wire w6392;
	wire w6393;
	wire w6394;
	wire w6395;
	wire w6396;
	wire w6397;
	wire w6398;
	wire w6399;
	wire w6400;
	wire w6401;
	wire w6402;
	wire w6403;
	wire w6404;
	wire w6405;
	wire w6406;
	wire w6407;
	wire w6408;
	wire w6409;
	wire w6410;
	wire w6411;
	wire w6412;
	wire w6413;
	wire w6414;
	wire w6415;
	wire w6416;
	wire w6417;
	wire w6418;
	wire w6419;
	wire w6420;
	wire w6421;
	wire w6422;
	wire w6423;
	wire w6424;
	wire w6425;
	wire w6426;
	wire w6427;
	wire w6428;
	wire w6429;
	wire w6430;
	wire w6431;
	wire w6432;
	wire w6433;
	wire w6434;
	wire w6435;
	wire w6436;
	wire w6437;
	wire w6438;
	wire w6439;
	wire w6440;
	wire w6441;
	wire w6442;
	wire w6443;
	wire w6444;
	wire w6445;
	wire w6446;
	wire w6447;
	wire w6448;
	wire w6449;
	wire w6450;
	wire w6451;
	wire w6452;
	wire w6453;
	wire w6454;
	wire w6455;
	wire w6456;
	wire w6457;
	wire w6458;
	wire w6459;
	wire w6460;
	wire w6461;
	wire w6462;
	wire w6463;
	wire w6464;
	wire w6465;
	wire w6466;
	wire w6467;
	wire w6468;
	wire w6469;
	wire w6470;
	wire w6471;
	wire w6472;
	wire w6473;
	wire w6474;
	wire w6475;
	wire w6476;
	wire w6477;
	wire w6478;
	wire w6479;
	wire w6480;
	wire w6481;
	wire w6482;
	wire w6483;
	wire w6484;
	wire w6485;
	wire w6486;
	wire w6487;
	wire w6488;
	wire w6489;
	wire w6490;
	wire w6491;
	wire w6492;
	wire w6493;
	wire w6494;
	wire w6495;
	wire w6496;
	wire w6497;
	wire w6498;
	wire w6499;
	wire w6500;
	wire w6501;
	wire w6502;
	wire w6503;
	wire w6504;
	wire w6505;
	wire w6506;
	wire w6507;
	wire w6508;
	wire w6509;
	wire w6510;
	wire w6511;
	wire w6512;
	wire w6513;
	wire w6514;
	wire w6515;
	wire w6516;
	wire w6517;
	wire w6518;
	wire w6519;
	wire w6520;
	wire w6521;
	wire w6522;
	wire w6523;
	wire w6524;
	wire w6525;
	wire w6526;
	wire w6527;
	wire w6528;
	wire w6529;
	wire w6530;
	wire w6531;
	wire w6532;
	wire w6533;
	wire w6534;
	wire w6535;
	wire w6536;
	wire w6537;
	wire w6538;
	wire w6539;
	wire w6540;
	wire w6541;
	wire w6542;
	wire w6543;
	wire w6544;
	wire w6545;
	wire w6546;
	wire w6547;
	wire w6548;
	wire w6549;
	wire w6550;
	wire w6551;
	wire w6552;
	wire w6553;
	wire w6554;
	wire w6555;
	wire w6556;
	wire w6557;
	wire w6558;
	wire w6559;
	wire w6560;
	wire w6561;
	wire w6562;
	wire w6563;
	wire w6564;
	wire w6565;
	wire w6566;
	wire w6567;
	wire w6568;
	wire w6569;
	wire w6570;
	wire w6571;
	wire w6572;
	wire w6573;
	wire w6574;
	wire w6575;
	wire w6576;
	wire w6577;
	wire w6578;
	wire w6579;
	wire w6580;
	wire w6581;
	wire w6582;
	wire w6583;
	wire w6584;
	wire w6585;
	wire w6586;
	wire w6587;
	wire w6588;
	wire w6589;
	wire w6590;
	wire w6591;
	wire w6592;
	wire w6593;
	wire w6594;
	wire w6595;
	wire w6596;
	wire w6597;
	wire w6598;
	wire w6599;
	wire w6600;
	wire w6601;
	wire w6602;
	wire w6603;
	wire w6604;
	wire w6605;
	wire w6606;
	wire w6607;
	wire w6608;
	wire w6609;
	wire w6610;
	wire w6611;
	wire w6612;
	wire w6613;
	wire w6614;
	wire w6615;
	wire w6616;

	assign CH0_EN = w1941;
	assign CH0VOL[0] = w1944;
	assign CH0VOL[1] = w1945;
	assign CH1_EN = w1942;
	assign CH1VOL[0] = w2004;
	assign CH1VOL[1] = w2005;
	assign CH2_EN = w1939;
	assign CH2VOL[0] = w2024;
	assign CH2VOL[1] = w2023;
	assign CH3_EN = w1940;
	assign CH3VOL[0] = w2046;
	assign CH3VOL[1] = w2045;
	assign PSGDAC0[0] = w1946;
	assign PSGDAC0[1] = w1947;
	assign PSGDAC0[2] = w1948;
	assign PSGDAC0[3] = w1949;
	assign PSGDAC0[4] = w1950;
	assign PSGDAC0[5] = w1951;
	assign PSGDAC0[6] = w1952;
	assign PSGDAC0[7] = w1953;
	assign PSGDAC1[0] = w2006;
	assign PSGDAC1[1] = w2007;
	assign PSGDAC1[2] = w2008;
	assign PSGDAC1[3] = w2009;
	assign PSGDAC1[4] = w2010;
	assign PSGDAC1[5] = w2011;
	assign PSGDAC1[6] = w2012;
	assign PSGDAC1[7] = w2013;
	assign PSGDAC2[0] = w2035;
	assign PSGDAC2[1] = w2036;
	assign PSGDAC2[2] = w2037;
	assign PSGDAC2[3] = w2038;
	assign PSGDAC2[4] = w2039;
	assign PSGDAC2[5] = w2040;
	assign PSGDAC2[6] = w2041;
	assign PSGDAC2[7] = w2042;
	assign PSGDAC3[0] = w2044;
	assign PSGDAC3[1] = w2043;
	assign PSGDAC3[2] = w2051;
	assign PSGDAC3[3] = w2050;
	assign PSGDAC3[4] = w2049;
	assign PSGDAC3[5] = w2048;
	assign PSGDAC3[6] = w2047;
	assign PSGDAC3[7] = w2052;
	assign w1156 = CAi[22];
	assign CAo[22] = w1304;
	assign CA[19] = CA[19];
	assign DTACK_OUT = w1013;
	assign Z80_INT = w1014;
	assign RA[7] = w1063;
	assign RA[6] = w1075;
	assign RA[5] = w1064;
	assign RA[4] = w1065;
	assign RA[2] = w1067;
	assign RA[1] = w1074;
	assign RA[0] = w1068;
	assign nRAS0 = w1371;
	assign RA[3] = w1066;
	assign nCAS0 = w1370;
	assign nOE0 = w1340;
	assign nLWR = w1341;
	assign nUWR = w1259;
	assign w1328 = DTACK_IN;
	assign w958 = RnW;
	assign w1323 = nLDS;
	assign w1315 = nUDS;
	assign w1204 = nAS;
	assign w1313 = nM1;
	assign w1314 = nWR;
	assign w1311 = nRD;
	assign w1312 = nIORQ;
	assign nILP2 = w1317;
	assign nILP1 = w1316;
	assign w1186 = nINTAK;
	assign w1310 = nMREQ;
	assign w1187 = nBG;
	assign BGACK_OUT = w1202;
	assign w1327 = BGACK_IN;
	assign nBR = w1372;
	assign VSYNC = w1913;
	assign nCSYNC = w1927;
	assign w1632 = nCSYNC_IN;
	assign nHSYNC = w1694;
	assign w1896 = nHSYNC_IN;
	assign DB[15] = DB[15];
	assign DB[14] = DB[14];
	assign DB[13] = DB[13];
	assign DB[12] = DB[12];
	assign DB[11] = DB[11];
	assign DB[10] = DB[10];
	assign DB[9] = DB[9];
	assign DB[8] = DB[8];
	assign DB[7] = DB[7];
	assign DB[6] = DB[6];
	assign DB[5] = DB[5];
	assign DB[4] = DB[4];
	assign DB[3] = DB[3];
	assign DB[2] = DB[2];
	assign DB[1] = DB[1];
	assign DB[0] = DB[0];
	assign CA[0] = CA[0];
	assign CA[1] = CA[1];
	assign CA[2] = CA[2];
	assign CA[3] = CA[3];
	assign CA[4] = CA[4];
	assign CA[5] = CA[5];
	assign CA[6] = CA[6];
	assign CA[7] = CA[7];
	assign CA[8] = CA[8];
	assign CA[9] = CA[9];
	assign CA[10] = CA[10];
	assign CA[11] = CA[11];
	assign CA[12] = CA[12];
	assign CA[13] = CA[13];
	assign CA[14] = CA[14];
	assign CA[15] = CA[15];
	assign CA[17] = CA[17];
	assign CA[18] = CA[18];
	assign CA[20] = CA[20];
	assign CA[21] = CA[21];
	assign R_DAC[0] = w2848;
	assign R_DAC[1] = w2813;
	assign R_DAC[2] = w2847;
	assign R_DAC[3] = w2812;
	assign R_DAC[4] = w2846;
	assign R_DAC[5] = w2845;
	assign R_DAC[6] = w2844;
	assign R_DAC[7] = w2843;
	assign R_DAC[8] = w2809;
	assign G_DAC[0] = w2841;
	assign G_DAC[1] = w2840;
	assign G_DAC[2] = w2803;
	assign G_DAC[3] = w2802;
	assign G_DAC[4] = w2801;
	assign G_DAC[5] = w2800;
	assign G_DAC[6] = w2799;
	assign G_DAC[7] = w2798;
	assign G_DAC[8] = w2797;
	assign R_DAC[9] = w2810;
	assign R_DAC[10] = w2807;
	assign R_DAC[11] = w2811;
	assign R_DAC[12] = w2806;
	assign R_DAC[13] = w2808;
	assign R_DAC[14] = w2805;
	assign R_DAC[15] = w2804;
	assign R_DAC[16] = w2842;
	assign B_DAC[0] = w2789;
	assign B_DAC[1] = w2839;
	assign B_DAC[2] = w2835;
	assign B_DAC[3] = w2836;
	assign B_DAC[4] = w2837;
	assign B_DAC[5] = w2834;
	assign B_DAC[6] = w2838;
	assign B_DAC[7] = w2894;
	assign B_DAC[8] = w2790;
	assign G_DAC[9] = w2791;
	assign G_DAC[10] = w2796;
	assign G_DAC[11] = w2795;
	assign G_DAC[12] = w2892;
	assign G_DAC[13] = w2794;
	assign G_DAC[14] = w2793;
	assign G_DAC[15] = w2792;
	assign G_DAC[16] = w2893;
	assign B_DAC[9] = w2787;
	assign B_DAC[10] = w2788;
	assign B_DAC[11] = w2833;
	assign B_DAC[12] = w2832;
	assign B_DAC[13] = w2831;
	assign B_DAC[14] = w2830;
	assign B_DAC[15] = w2828;
	assign B_DAC[16] = w2829;
	assign nOE1 = nOE1;
	assign nWE0 = nWE0;
	assign nWE1 = nWE1;
	assign nCAS1 = nCAS1;
	assign nRAS1 = nRAS1;
	assign AD_RD_DIR = AD_RD_DIR;
	assign nYS = nYS;
	assign nSC = w2512;
	assign nSE0_1 = w2407;
	assign ADo[7] = w2490;
	assign ADo[6] = w2600;
	assign ADo[5] = w2589;
	assign ADo[4] = w2602;
	assign ADo[3] = w2594;
	assign ADo[2] = w2592;
	assign ADo[1] = w2601;
	assign ADo[0] = w2590;
	assign RDo[6] = w2550;
	assign RDo[5] = w2568;
	assign RDo[4] = w2554;
	assign RDo[3] = w2553;
	assign RDo[2] = w2569;
	assign RDo[1] = w2591;
	assign RDo[0] = w2414;
	assign w2453 = RDi[6];
	assign w2370 = RDi[7];
	assign w2382 = RDi[4];
	assign w2579 = RDi[5];
	assign w2447 = RDi[2];
	assign w2455 = RDi[3];
	assign w2612 = RDi[0];
	assign w2489 = RDi[1];
	assign w2454 = ADi[6];
	assign w2607 = ADi[7];
	assign w2400 = ADi[4];
	assign w2606 = ADi[5];
	assign w2442 = ADi[2];
	assign w2446 = ADi[3];
	assign w2415 = ADi[0];
	assign w2434 = ADi[1];
	assign RDo[7] = w2552;
	assign w5096 = SD[7];
	assign w5097 = SD[6];
	assign w6418 = SD[5];
	assign w6420 = SD[4];
	assign w5098 = SD[3];
	assign w5095 = SD[2];
	assign w6419 = SD[1];
	assign w5094 = SD[0];
	assign CLK1 = M68K_CPU_CLOCK;
	assign CLK0 = w1343;
	assign w4331 = EDCLKi;
	assign EDCLKo = EDCLK_O;
	assign w4309 = MCLK;
	assign SUB_CLK = w4298;
	assign w4349 = nRES_PAD;
	assign w1373 = M68kCLKi;
	assign EDCLKd = w1431;
	assign CA_PAD_DIR = w2367;
	assign DB_PAD_DIR = w2368;
	assign nSEL0_M3 = nSEL0_M3;
	assign w6424 = nPAL;
	assign w406 = nHL;
	assign SPA_Bo = w2722;
	assign w2699 = SPA_Bi;

	// Instances

	vdp_slatch g1 (.nQ(w330), .D(VPOS[7]), .C(w1507), .nC(w1508) );
	vdp_slatch g2 (.nQ(w1470), .D(HPOS[8]), .C(w351), .nC(w352) );
	vdp_slatch g3 (.nQ(w335), .D(w277), .C(w1403), .nC(w353) );
	vdp_slatch g4 (.D(w278), .C(w1505), .nC(w1506), .nQ(w6526) );
	vdp_slatch g5 (.nQ(w336), .D(w337), .C(w1503), .nC(w1504) );
	vdp_slatch g6 (.nQ(w280), .D(w281), .C(w1501), .nC(w1502) );
	vdp_slatch g7 (.nQ(w338), .D(w337), .C(w354), .nC(w355) );
	vdp_slatch g8 (.nQ(w341), .D(w281), .C(w356), .nC(w357) );
	vdp_slatch g9 (.nQ(w339), .D(w337), .C(w395), .nC(w1400) );
	vdp_slatch g10 (.nQ(w342), .D(w281), .C(w1399), .nC(w362) );
	vdp_slatch g11 (.nQ(w340), .D(w337), .C(w360), .nC(w359) );
	vdp_slatch g12 (.nQ(w283), .D(w281), .C(w358), .nC(w1398) );
	vdp_slatch g13 (.Q(w281), .D(DB[7]), .C(w344), .nC(w343) );
	vdp_slatch g14 (.Q(w337), .D(w890), .C(w347), .nC(w346) );
	vdp_sr_bit g15 (.D(w284), .C2(HCLK2), .C1(HCLK1), .Q(FIFOo[7]), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g16 (.A(1'b1), .nZ(DB[7]), .nE(w1397) );
	vdp_notif0 g17 (.A(w283), .nZ(w284), .nE(w1943) );
	vdp_notif0 g18 (.A(w340), .nZ(w334), .nE(w361) );
	vdp_notif0 g19 (.A(w282), .nZ(AD_DATA[7]), .nE(w1551) );
	vdp_notif0 g20 (.A(w342), .nZ(w284), .nE(w1500) );
	vdp_notif0 g21 (.A(w339), .nZ(w334), .nE(w1550) );
	vdp_notif0 g22 (.A(w1476), .nZ(AD_DATA[7]), .nE(w371) );
	vdp_notif0 g23 (.A(w341), .nZ(w284), .nE(w370) );
	vdp_notif0 g24 (.A(w338), .nZ(w334), .nE(w1401) );
	vdp_notif0 g25 (.A(w1475), .nZ(AD_DATA[7]), .nE(w384) );
	vdp_notif0 g26 (.A(w280), .nZ(w284), .nE(w363) );
	vdp_notif0 g27 (.A(w279), .nZ(AD_DATA[7]), .nE(w383) );
	vdp_notif0 g28 (.A(w335), .nZ(DB[7]), .nE(w1547) );
	vdp_notif0 g29 (.nZ(DB[15]), .nE(w364), .A(w6526) );
	vdp_notif0 g30 (.A(w336), .nZ(w334), .nE(w1548) );
	vdp_notif0 g31 (.A(w330), .nZ(DB[15]), .nE(w1546) );
	vdp_notif0 g32 (.A(w398), .nZ(DB[7]), .nE(w365) );
	vdp_aon22 g33 (.Z(w398), .A1(w1470), .A2(w1509), .B1(w369), .B2(w330) );
	vdp_aon22 g34 (.A2(w367), .B1(w368), .B2(AD_DATA[7]), .A1(w334), .Z(w277) );
	vdp_aon22 g35 (.A2(w6432), .B1(w6433), .B2(w334), .A1(AD_DATA[7]), .Z(w278) );
	vdp_aon22 g36 (.Z(w279), .A2(w366), .B1(w1510), .B2(w280), .A1(w336) );
	vdp_aon22 g37 (.Z(w1475), .A2(w389), .B1(w388), .B2(w338), .A1(w341) );
	vdp_aon22 g38 (.Z(w1476), .A2(w396), .B1(w397), .B2(w339), .A1(w342) );
	vdp_aon22 g39 (.Z(w282), .A2(w6428), .B1(w6429), .B2(w283), .A1(w340) );
	vdp_aon22 g40 (.Z(w890), .A1(DB[15]), .A2(w345), .B1(w349), .B2(DB[7]) );
	vdp_slatch g41 (.nQ(w204), .D(VPOS[6]), .C(w1507), .nC(w1508) );
	vdp_slatch g42 (.nQ(w207), .D(HPOS[7]), .C(w351), .nC(w352) );
	vdp_slatch g43 (.nQ(w209), .D(w243), .C(w1403), .nC(w353) );
	vdp_slatch g44 (.nQ(w244), .D(w1366), .C(w1505), .nC(w1506) );
	vdp_slatch g45 (.nQ(w210), .D(w211), .C(w1503), .nC(w1504) );
	vdp_slatch g46 (.nQ(w246), .D(w247), .C(w1501), .nC(w1502) );
	vdp_slatch g47 (.nQ(w212), .D(w211), .C(w354), .nC(w355) );
	vdp_slatch g48 (.nQ(w214), .D(w247), .C(w356), .nC(w357) );
	vdp_slatch g49 (.nQ(w215), .D(w211), .C(w395), .nC(w1400) );
	vdp_slatch g50 (.nQ(w217), .D(w247), .C(w1399), .nC(w362) );
	vdp_slatch g51 (.nQ(w218), .D(w211), .C(w360), .nC(w359) );
	vdp_slatch g52 (.nQ(w249), .D(w247), .C(w358), .nC(w1398) );
	vdp_slatch g53 (.Q(w247), .D(DB[6]), .C(w344), .nC(w343) );
	vdp_slatch g54 (.Q(w211), .D(w250), .C(w347), .nC(w346) );
	vdp_sr_bit g55 (.D(w1466), .Q(FIFOo[6]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g56 (.A(1'b1), .nZ(DB[6]), .nE(w1397) );
	vdp_notif0 g57 (.A(w249), .nZ(w1466), .nE(w1943) );
	vdp_notif0 g58 (.A(w218), .nZ(RD_DATA[6]), .nE(w361) );
	vdp_notif0 g59 (.A(w248), .nZ(AD_DATA[6]), .nE(w1551) );
	vdp_notif0 g60 (.A(w217), .nZ(w1466), .nE(w1500) );
	vdp_notif0 g61 (.A(w215), .nZ(RD_DATA[6]), .nE(w1550) );
	vdp_notif0 g62 (.A(w216), .nZ(AD_DATA[6]), .nE(w371) );
	vdp_notif0 g63 (.A(w214), .nZ(w1466), .nE(w370) );
	vdp_notif0 g64 (.A(w212), .nZ(RD_DATA[6]), .nE(w1401) );
	vdp_notif0 g65 (.A(w213), .nZ(AD_DATA[6]), .nE(w384) );
	vdp_notif0 g66 (.A(w246), .nZ(w1466), .nE(w363) );
	vdp_notif0 g67 (.A(w245), .nZ(AD_DATA[6]), .nE(w383) );
	vdp_notif0 g68 (.A(w209), .nZ(DB[6]), .nE(w1547) );
	vdp_notif0 g69 (.A(w244), .nZ(DB[14]), .nE(w364) );
	vdp_notif0 g70 (.A(w210), .nZ(RD_DATA[6]), .nE(w1548) );
	vdp_notif0 g71 (.A(w204), .nZ(DB[14]), .nE(w1546) );
	vdp_notif0 g72 (.A(w208), .nZ(DB[6]), .nE(w365) );
	vdp_aon22 g73 (.A2(w1509), .B1(w369), .B2(w204), .A1(w207), .Z(w208) );
	vdp_aon22 g74 (.Z(w243), .A2(w367), .B1(w368), .B2(AD_DATA[6]), .A1(RD_DATA[6]) );
	vdp_aon22 g75 (.Z(w1366), .A2(w6432), .B1(w6433), .B2(RD_DATA[6]), .A1(AD_DATA[6]) );
	vdp_aon22 g76 (.Z(w245), .A2(w366), .B1(w1510), .B2(w246), .A1(w210) );
	vdp_aon22 g77 (.Z(w213), .A2(w389), .B1(w388), .B2(w214), .A1(w212) );
	vdp_aon22 g78 (.Z(w216), .A2(w396), .B1(w397), .B2(w217), .A1(w215) );
	vdp_aon22 g79 (.Z(w248), .A2(w6428), .B1(w6429), .B2(w249), .A1(w218) );
	vdp_aon22 g80 (.Z(w250), .A1(DB[14]), .A2(w345), .B1(w349), .B2(DB[6]) );
	vdp_slatch g81 (.nQ(w314), .D(VPOS[5]), .C(w1507), .nC(w1508) );
	vdp_slatch g82 (.nQ(w1471), .D(HPOS[6]), .C(w351), .nC(w352) );
	vdp_slatch g83 (.nQ(w319), .D(w268), .C(w1403), .nC(w353) );
	vdp_slatch g84 (.D(w269), .C(w1505), .nC(w1506), .nQ(w6527) );
	vdp_slatch g85 (.nQ(w320), .D(w326), .C(w1503), .nC(w1504) );
	vdp_slatch g86 (.nQ(w271), .D(w272), .C(w1501), .nC(w1502) );
	vdp_slatch g87 (.nQ(w322), .D(w326), .C(w354), .nC(w355) );
	vdp_slatch g88 (.nQ(w321), .D(w272), .C(w356), .nC(w357) );
	vdp_slatch g89 (.nQ(w324), .D(w326), .C(w395), .nC(w1400) );
	vdp_slatch g90 (.nQ(w327), .D(w272), .C(w1399), .nC(w362) );
	vdp_slatch g91 (.nQ(w328), .D(w326), .C(w360), .nC(w359) );
	vdp_slatch g92 (.nQ(w274), .D(w272), .C(w358), .nC(w1398) );
	vdp_slatch g93 (.Q(w272), .D(DB[5]), .C(w344), .nC(w343) );
	vdp_slatch g94 (.Q(w326), .D(w275), .C(w347), .nC(w346) );
	vdp_sr_bit g95 (.D(w276), .Q(FIFOo[5]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g96 (.A(1'b1), .nZ(DB[5]), .nE(w1397) );
	vdp_notif0 g97 (.A(w274), .nZ(w276), .nE(w1943) );
	vdp_notif0 g98 (.A(w328), .nZ(RD_DATA[5]), .nE(w361) );
	vdp_notif0 g99 (.A(w273), .nZ(AD_DATA[5]), .nE(w1551) );
	vdp_notif0 g100 (.A(w327), .nZ(w276), .nE(w1500) );
	vdp_notif0 g101 (.A(w324), .nZ(RD_DATA[5]), .nE(w1550) );
	vdp_notif0 g102 (.A(w325), .nZ(AD_DATA[5]), .nE(w371) );
	vdp_notif0 g103 (.A(w321), .nZ(w276), .nE(w370) );
	vdp_notif0 g104 (.A(w322), .nZ(RD_DATA[5]), .nE(w1401) );
	vdp_notif0 g105 (.A(w323), .nZ(AD_DATA[5]), .nE(w384) );
	vdp_notif0 g106 (.A(w271), .nZ(w276), .nE(w363) );
	vdp_notif0 g107 (.A(w270), .nZ(AD_DATA[5]), .nE(w383) );
	vdp_notif0 g108 (.A(w319), .nZ(DB[5]), .nE(w1547) );
	vdp_notif0 g109 (.nZ(DB[13]), .nE(w364), .A(w6527) );
	vdp_notif0 g110 (.A(w320), .nZ(RD_DATA[5]), .nE(w1548) );
	vdp_notif0 g111 (.A(w314), .nZ(DB[13]), .nE(w1546) );
	vdp_notif0 g112 (.A(w318), .nZ(DB[5]), .nE(w365) );
	vdp_aon22 g113 (.Z(w318), .A1(w1471), .A2(w1509), .B1(w369), .B2(w314) );
	vdp_aon22 g114 (.A2(w367), .B1(w368), .B2(AD_DATA[5]), .A1(RD_DATA[5]), .Z(w268) );
	vdp_aon22 g115 (.A2(w6432), .B1(w6433), .B2(RD_DATA[5]), .A1(AD_DATA[5]), .Z(w269) );
	vdp_aon22 g116 (.Z(w270), .A2(w366), .B1(w1510), .B2(w271), .A1(w320) );
	vdp_aon22 g117 (.Z(w323), .A2(w389), .B1(w388), .B2(w322), .A1(w321) );
	vdp_aon22 g118 (.Z(w325), .A2(w396), .B1(w397), .B2(w324), .A1(w327) );
	vdp_aon22 g119 (.Z(w273), .A2(w6428), .B1(w6429), .B2(w274), .A1(w328) );
	vdp_aon22 g120 (.Z(w275), .A1(DB[13]), .A2(w345), .B1(w349), .B2(DB[5]) );
	vdp_slatch g121 (.nQ(w189), .D(VPOS[4]), .C(w1507), .nC(w1508) );
	vdp_slatch g122 (.nQ(w192), .D(HPOS[5]), .C(w351), .nC(w352) );
	vdp_slatch g123 (.nQ(w1511), .D(w236), .C(w1403), .nC(w353) );
	vdp_slatch g124 (.D(w1474), .C(w1505), .nC(w1506), .nQ(w6528) );
	vdp_slatch g125 (.nQ(w194), .D(w195), .C(w1503), .nC(w1504) );
	vdp_slatch g126 (.nQ(w238), .D(w239), .C(w1501), .nC(w1502) );
	vdp_slatch g127 (.nQ(w196), .D(w195), .C(w354), .nC(w355) );
	vdp_slatch g128 (.nQ(w198), .D(w239), .C(w356), .nC(w357) );
	vdp_slatch g129 (.nQ(w199), .D(w195), .C(w395), .nC(w1400) );
	vdp_slatch g130 (.nQ(w201), .D(w239), .C(w1399), .nC(w362) );
	vdp_slatch g131 (.nQ(w202), .D(w195), .C(w360), .nC(w359) );
	vdp_slatch g132 (.nQ(w241), .D(w239), .C(w358), .nC(w1398) );
	vdp_slatch g133 (.Q(w239), .D(DB[4]), .C(w344), .nC(w343) );
	vdp_slatch g134 (.Q(w195), .D(w888), .C(w347), .nC(w346) );
	vdp_sr_bit g135 (.D(w242), .Q(FIFOo[4]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g136 (.A(1'b1), .nZ(DB[4]), .nE(w1397) );
	vdp_notif0 g137 (.A(w241), .nZ(w242), .nE(w1943) );
	vdp_notif0 g138 (.A(w202), .nZ(RD_DATA[4]), .nE(w361) );
	vdp_notif0 g139 (.A(w240), .nZ(AD_DATA[4]), .nE(w1551) );
	vdp_notif0 g140 (.A(w201), .nZ(w242), .nE(w1500) );
	vdp_notif0 g141 (.A(w199), .nZ(RD_DATA[4]), .nE(w1550) );
	vdp_notif0 g142 (.A(w200), .nZ(AD_DATA[4]), .nE(w371) );
	vdp_notif0 g143 (.A(w198), .nZ(w242), .nE(w370) );
	vdp_notif0 g144 (.A(w196), .nZ(RD_DATA[4]), .nE(w1401) );
	vdp_notif0 g145 (.A(w197), .nZ(AD_DATA[4]), .nE(w384) );
	vdp_notif0 g146 (.A(w238), .nZ(w242), .nE(w363) );
	vdp_notif0 g147 (.A(w237), .nZ(AD_DATA[4]), .nE(w383) );
	vdp_notif0 g148 (.A(w1511), .nZ(DB[4]), .nE(w1547) );
	vdp_notif0 g149 (.nZ(DB[12]), .nE(w364), .A(w6528) );
	vdp_notif0 g150 (.A(w194), .nZ(RD_DATA[4]), .nE(w1548) );
	vdp_notif0 g151 (.A(w189), .nZ(DB[12]), .nE(w1546) );
	vdp_notif0 g152 (.A(w193), .nZ(DB[4]), .nE(w365) );
	vdp_aon22 g153 (.A2(w1509), .B1(w369), .B2(w189), .A1(w192), .Z(w193) );
	vdp_aon22 g154 (.Z(w236), .A2(w367), .B1(w368), .B2(AD_DATA[4]), .A1(RD_DATA[4]) );
	vdp_aon22 g155 (.Z(w1474), .A2(w6432), .B1(w6433), .B2(RD_DATA[4]), .A1(AD_DATA[4]) );
	vdp_aon22 g156 (.Z(w237), .A2(w366), .B1(w1510), .B2(w238), .A1(w194) );
	vdp_aon22 g157 (.Z(w197), .A2(w389), .B1(w388), .B2(w198), .A1(w196) );
	vdp_aon22 g158 (.Z(w200), .A2(w396), .B1(w397), .B2(w201), .A1(w199) );
	vdp_aon22 g159 (.Z(w240), .A2(w6428), .B1(w6429), .B2(w241), .A1(w202) );
	vdp_aon22 g160 (.Z(w888), .A1(DB[12]), .A2(w345), .B1(w349), .B2(DB[4]) );
	vdp_slatch g161 (.nQ(w298), .D(VPOS[3]), .C(w1507), .nC(w1508) );
	vdp_slatch g162 (.nQ(w1472), .D(HPOS[4]), .C(w351), .nC(w352) );
	vdp_slatch g163 (.nQ(w303), .D(w260), .C(w1403), .nC(w353) );
	vdp_slatch g164 (.D(w261), .C(w1505), .nC(w1506), .nQ(w6529) );
	vdp_slatch g165 (.nQ(w304), .D(w307), .C(w1503), .nC(w1504) );
	vdp_slatch g166 (.nQ(w263), .D(w264), .C(w1501), .nC(w1502) );
	vdp_slatch g167 (.nQ(w305), .D(w307), .C(w354), .nC(w355) );
	vdp_slatch g168 (.nQ(w306), .D(w264), .C(w356), .nC(w357) );
	vdp_slatch g169 (.nQ(w309), .D(w307), .C(w395), .nC(w1400) );
	vdp_slatch g170 (.nQ(w311), .D(w264), .C(w1399), .nC(w362) );
	vdp_slatch g171 (.nQ(w312), .D(w307), .C(w360), .nC(w359) );
	vdp_slatch g172 (.nQ(w266), .D(w264), .C(w358), .nC(w1398) );
	vdp_slatch g173 (.Q(w264), .D(DB[3]), .C(w344), .nC(w343) );
	vdp_slatch g174 (.Q(w307), .D(w267), .C(w347), .nC(w346) );
	vdp_sr_bit g175 (.D(w1465), .Q(FIFOo[3]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g176 (.A(1'b1), .nZ(DB[3]), .nE(w1397) );
	vdp_notif0 g177 (.A(w266), .nZ(w1465), .nE(w1943) );
	vdp_notif0 g178 (.A(w312), .nZ(w300), .nE(w361) );
	vdp_notif0 g179 (.A(w265), .nZ(AD_DATA[3]), .nE(w1551) );
	vdp_notif0 g180 (.A(w311), .nZ(w1465), .nE(w1500) );
	vdp_notif0 g181 (.A(w309), .nZ(w300), .nE(w1550) );
	vdp_notif0 g182 (.A(w310), .nZ(AD_DATA[3]), .nE(w371) );
	vdp_notif0 g183 (.A(w306), .nZ(w1465), .nE(w370) );
	vdp_notif0 g184 (.A(w305), .nZ(w300), .nE(w1401) );
	vdp_notif0 g185 (.A(w308), .nZ(AD_DATA[3]), .nE(w384) );
	vdp_notif0 g186 (.A(w263), .nZ(w1465), .nE(w363) );
	vdp_notif0 g187 (.A(w262), .nZ(AD_DATA[3]), .nE(w383) );
	vdp_notif0 g188 (.A(w303), .nZ(DB[3]), .nE(w1547) );
	vdp_notif0 g189 (.nZ(DB[11]), .nE(w364), .A(w6529) );
	vdp_notif0 g190 (.A(w304), .nZ(w300), .nE(w1548) );
	vdp_notif0 g191 (.A(w298), .nZ(DB[11]), .nE(w1546) );
	vdp_notif0 g192 (.A(w302), .nZ(DB[3]), .nE(w365) );
	vdp_aon22 g193 (.Z(w302), .A1(w1472), .A2(w1509), .B1(w369), .B2(w298) );
	vdp_aon22 g194 (.A2(w367), .B1(w368), .B2(AD_DATA[3]), .A1(w300), .Z(w260) );
	vdp_aon22 g195 (.A2(w6432), .B1(w6433), .B2(w300), .A1(AD_DATA[3]), .Z(w261) );
	vdp_aon22 g196 (.Z(w262), .A2(w366), .B1(w1510), .B2(w263), .A1(w304) );
	vdp_aon22 g197 (.Z(w308), .A2(w389), .B1(w388), .B2(w305), .A1(w306) );
	vdp_aon22 g198 (.Z(w310), .A2(w396), .B1(w397), .B2(w309), .A1(w311) );
	vdp_aon22 g199 (.Z(w265), .A2(w6428), .B1(w6429), .B2(w266), .A1(w312) );
	vdp_aon22 g200 (.Z(w267), .A1(DB[11]), .A2(w345), .B1(w349), .B2(DB[3]) );
	vdp_slatch g201 (.nQ(w174), .D(VPOS[2]), .C(w1507), .nC(w1508) );
	vdp_slatch g202 (.nQ(w1512), .D(HPOS[3]), .C(w351), .nC(w352) );
	vdp_slatch g203 (.nQ(w177), .D(w227), .C(w1403), .nC(w353) );
	vdp_slatch g204 (.D(w1404), .C(w1505), .nC(w1506), .nQ(w6530) );
	vdp_slatch g205 (.nQ(w178), .D(w181), .C(w1503), .nC(w1504) );
	vdp_slatch g206 (.nQ(w229), .D(w230), .C(w1501), .nC(w1502) );
	vdp_slatch g207 (.nQ(w179), .D(w181), .C(w354), .nC(w355) );
	vdp_slatch g208 (.nQ(w182), .D(w230), .C(w356), .nC(w357) );
	vdp_slatch g209 (.nQ(w183), .D(w181), .C(w395), .nC(w1400) );
	vdp_slatch g210 (.nQ(w185), .D(w230), .C(w1399), .nC(w362) );
	vdp_slatch g211 (.nQ(w186), .D(w181), .C(w360), .nC(w359) );
	vdp_slatch g212 (.nQ(w232), .D(w230), .C(w358), .nC(w1398) );
	vdp_slatch g213 (.Q(w230), .D(DB[2]), .C(w344), .nC(w343) );
	vdp_slatch g214 (.Q(w181), .D(w233), .C(w347), .nC(w346) );
	vdp_sr_bit g215 (.D(w235), .Q(FIFOo[2]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g216 (.A(w187), .nZ(DB[2]), .nE(w1397) );
	vdp_notif0 g217 (.A(w232), .nZ(w235), .nE(w1943) );
	vdp_notif0 g218 (.A(w186), .nZ(RD_DATA[2]), .nE(w361) );
	vdp_notif0 g219 (.A(w231), .nZ(AD_DATA[2]), .nE(w1551) );
	vdp_notif0 g220 (.A(w185), .nZ(w235), .nE(w1500) );
	vdp_notif0 g221 (.A(w183), .nZ(RD_DATA[2]), .nE(w1550) );
	vdp_notif0 g222 (.A(w184), .nZ(AD_DATA[2]), .nE(w371) );
	vdp_notif0 g223 (.A(w182), .nZ(w235), .nE(w370) );
	vdp_notif0 g224 (.A(w179), .nZ(RD_DATA[2]), .nE(w1401) );
	vdp_notif0 g225 (.A(w180), .nZ(AD_DATA[2]), .nE(w384) );
	vdp_notif0 g226 (.A(w229), .nZ(w235), .nE(w363) );
	vdp_notif0 g227 (.A(w228), .nZ(AD_DATA[2]), .nE(w383) );
	vdp_notif0 g228 (.A(w177), .nZ(DB[2]), .nE(w1547) );
	vdp_notif0 g229 (.nZ(DB[10]), .nE(w364), .A(w6530) );
	vdp_notif0 g230 (.A(w178), .nZ(RD_DATA[2]), .nE(w1548) );
	vdp_notif0 g231 (.A(w174), .nZ(DB[10]), .nE(w1546) );
	vdp_notif0 g232 (.A(w176), .nZ(DB[2]), .nE(w365) );
	vdp_aon22 g233 (.A2(w1509), .B1(w369), .B2(w174), .A1(w1512), .Z(w176) );
	vdp_aon22 g234 (.Z(w227), .A2(w367), .B1(w368), .B2(AD_DATA[2]), .A1(RD_DATA[2]) );
	vdp_aon22 g235 (.Z(w1404), .A2(w6432), .B1(w6433), .B2(RD_DATA[2]), .A1(AD_DATA[2]) );
	vdp_aon22 g236 (.Z(w228), .A2(w366), .B1(w1510), .B2(w229), .A1(w178) );
	vdp_aon22 g237 (.Z(w180), .A2(w389), .B1(w388), .B2(w182), .A1(w179) );
	vdp_aon22 g238 (.Z(w184), .A2(w396), .B1(w397), .B2(w185), .A1(w183) );
	vdp_aon22 g239 (.Z(w231), .A2(w6428), .B1(w6429), .B2(w232), .A1(w186) );
	vdp_aon22 g240 (.Z(w233), .A1(DB[10]), .A2(w345), .B1(w349), .B2(DB[2]) );
	vdp_slatch g241 (.nQ(w285), .D(VPOS[1]), .C(w1507), .nC(w1508) );
	vdp_slatch g242 (.nQ(w1473), .D(HPOS[2]), .C(w351), .nC(w352) );
	vdp_slatch g243 (.nQ(w288), .D(w251), .C(w1403), .nC(w353) );
	vdp_slatch g244 (.D(w252), .C(w1505), .nC(w1506), .nQ(w6531) );
	vdp_slatch g245 (.nQ(w289), .D(w292), .C(w1503), .nC(w1504) );
	vdp_slatch g246 (.nQ(w254), .D(w255), .C(w1501), .nC(w1502) );
	vdp_slatch g247 (.nQ(w291), .D(w292), .C(w354), .nC(w355) );
	vdp_slatch g248 (.nQ(w290), .D(w255), .C(w356), .nC(w357) );
	vdp_slatch g249 (.nQ(w294), .D(w292), .C(w395), .nC(w1400) );
	vdp_slatch g250 (.nQ(w296), .D(w255), .C(w1399), .nC(w362) );
	vdp_slatch g251 (.nQ(w297), .D(w292), .C(w360), .nC(w359) );
	vdp_slatch g252 (.nQ(w257), .D(w255), .C(w358), .nC(w1398) );
	vdp_slatch g253 (.Q(w255), .D(DB[1]), .C(w344), .nC(w343) );
	vdp_slatch g254 (.Q(w292), .D(w259), .C(w347), .nC(w346) );
	vdp_sr_bit g255 (.D(w1396), .Q(FIFOo[1]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g256 (.A(w1552), .nZ(DB[1]), .nE(w1397) );
	vdp_notif0 g257 (.A(w257), .nZ(w1396), .nE(w1943) );
	vdp_notif0 g258 (.A(w297), .nZ(RD_DATA[1]), .nE(w361) );
	vdp_notif0 g259 (.A(w256), .nZ(AD_DATA[1]), .nE(w1551) );
	vdp_notif0 g260 (.A(w296), .nZ(w1396), .nE(w1500) );
	vdp_notif0 g261 (.A(w294), .nZ(RD_DATA[1]), .nE(w1550) );
	vdp_notif0 g262 (.A(w295), .nZ(AD_DATA[1]), .nE(w371) );
	vdp_notif0 g263 (.A(w290), .nZ(w1396), .nE(w370) );
	vdp_notif0 g264 (.A(w291), .nZ(RD_DATA[1]), .nE(w1401) );
	vdp_notif0 g265 (.A(w293), .nZ(AD_DATA[1]), .nE(w384) );
	vdp_notif0 g266 (.A(w254), .nZ(w1396), .nE(w363) );
	vdp_notif0 g267 (.A(w253), .nZ(AD_DATA[1]), .nE(w383) );
	vdp_notif0 g268 (.A(w288), .nZ(DB[1]), .nE(w1547) );
	vdp_notif0 g269 (.nZ(DB[9]), .nE(w364), .A(w6531) );
	vdp_notif0 g270 (.A(w289), .nZ(RD_DATA[1]), .nE(w1548) );
	vdp_notif0 g271 (.A(w285), .nZ(DB[9]), .nE(w1546) );
	vdp_notif0 g272 (.A(w1402), .nZ(DB[1]), .nE(w365) );
	vdp_aon22 g273 (.Z(w1402), .A1(w1473), .A2(w1509), .B1(w369), .B2(w285) );
	vdp_aon22 g274 (.A2(w367), .B1(w368), .B2(AD_DATA[1]), .A1(RD_DATA[1]), .Z(w251) );
	vdp_aon22 g275 (.A2(w6432), .B1(w6433), .B2(RD_DATA[1]), .A1(AD_DATA[1]), .Z(w252) );
	vdp_aon22 g276 (.Z(w253), .A2(w366), .B1(w1510), .B2(w254), .A1(w289) );
	vdp_aon22 g277 (.Z(w293), .A2(w389), .B1(w388), .B2(w291), .A1(w290) );
	vdp_aon22 g278 (.Z(w295), .A2(w396), .B1(w397), .B2(w294), .A1(w296) );
	vdp_aon22 g279 (.Z(w256), .A2(w6428), .B1(w6429), .B2(w257), .A1(w297) );
	vdp_aon22 g280 (.Z(w259), .A1(DB[9]), .A2(w345), .B1(w349), .B2(DB[1]) );
	vdp_slatch g281 (.nQ(w159), .D(VPOS_80), .C(w1507), .nC(w1508) );
	vdp_slatch g282 (.D(HPOS[1]), .nQ(w1395), .C(w351), .nC(w352) );
	vdp_slatch g283 (.nQ(w162), .D(w220), .C(w1403), .nC(w353) );
	vdp_slatch g284 (.D(w1368), .C(w1505), .nC(w1506), .nQ(w6532) );
	vdp_slatch g285 (.nQ(w163), .D(w167), .C(w1503), .nC(w1504) );
	vdp_slatch g286 (.nQ(w222), .D(w223), .C(w1501), .nC(w1502) );
	vdp_slatch g287 (.nQ(w164), .D(w167), .C(w354), .nC(w355) );
	vdp_slatch g288 (.nQ(w166), .D(w223), .C(w356), .nC(w357) );
	vdp_slatch g289 (.nQ(w168), .D(w167), .C(w395), .nC(w1400) );
	vdp_slatch g290 (.nQ(w170), .D(w223), .C(w1399), .nC(w362) );
	vdp_slatch g291 (.nQ(w171), .D(w167), .C(w360), .nC(w359) );
	vdp_slatch g292 (.nQ(w225), .D(w223), .C(w358), .nC(w1398) );
	vdp_slatch g293 (.Q(w223), .D(DB[0]), .C(w344), .nC(w343) );
	vdp_slatch g294 (.D(w226), .Q(w167), .C(w347), .nC(w346) );
	vdp_sr_bit g295 (.D(w1549), .C2(HCLK2), .C1(HCLK1), .Q(FIFOo[0]), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g296 (.A(1'b1), .nZ(DB[0]), .nE(w1397) );
	vdp_notif0 g297 (.A(w225), .nZ(w1549), .nE(w1943) );
	vdp_notif0 g298 (.A(w171), .nZ(RD_DATA[0]), .nE(w361) );
	vdp_notif0 g299 (.A(w224), .nZ(AD_DATA[0]), .nE(w1551) );
	vdp_notif0 g300 (.A(w170), .nZ(w1549), .nE(w1500) );
	vdp_notif0 g301 (.A(w168), .nZ(RD_DATA[0]), .nE(w1550) );
	vdp_notif0 g302 (.A(w169), .nZ(AD_DATA[0]), .nE(w371) );
	vdp_notif0 g303 (.A(w166), .nZ(w1549), .nE(w370) );
	vdp_notif0 g304 (.A(w164), .nZ(RD_DATA[0]), .nE(w1401) );
	vdp_notif0 g305 (.A(w165), .nZ(AD_DATA[0]), .nE(w384) );
	vdp_notif0 g306 (.A(w222), .nZ(w1549), .nE(w363) );
	vdp_notif0 g307 (.A(w221), .nZ(AD_DATA[0]), .nE(w383) );
	vdp_notif0 g308 (.A(w162), .nZ(DB[0]), .nE(w1547) );
	vdp_notif0 g309 (.nZ(DB[8]), .nE(w364), .A(w6532) );
	vdp_notif0 g310 (.A(w163), .nZ(RD_DATA[0]), .nE(w1548) );
	vdp_notif0 g311 (.A(w159), .nZ(DB[8]), .nE(w1546) );
	vdp_notif0 g312 (.A(w161), .nZ(DB[0]), .nE(w365) );
	vdp_aon22 g313 (.A2(w1509), .B1(w369), .B2(w159), .A1(w1395), .Z(w161) );
	vdp_aon22 g314 (.Z(w220), .A2(w367), .B1(w368), .B2(AD_DATA[0]), .A1(RD_DATA[0]) );
	vdp_aon22 g315 (.Z(w1368), .A2(w6432), .B1(w6433), .B2(RD_DATA[0]), .A1(AD_DATA[0]) );
	vdp_aon22 g316 (.Z(w221), .A2(w366), .B1(w1510), .B2(w222), .A1(w163) );
	vdp_aon22 g317 (.Z(w165), .A2(w389), .B1(w388), .B2(w166), .A1(w164) );
	vdp_aon22 g318 (.Z(w169), .A2(w396), .B1(w397), .B2(w170), .A1(w168) );
	vdp_aon22 g319 (.Z(w224), .A2(w6428), .B1(w6429), .B2(w225), .A1(w171) );
	vdp_aon22 g320 (.Z(w226), .A1(DB[8]), .A2(w345), .B1(w349), .B2(DB[0]) );
	vdp_not g321 (.A(w258), .nZ(w1552) );
	vdp_not g322 (.A(w234), .nZ(w187) );
	vdp_not g323 (.A(w373), .nZ(w1546) );
	vdp_not g324 (.A(w377), .nZ(w365) );
	vdp_not g325 (.A(w382), .nZ(w1547) );
	vdp_not g326 (.A(w382), .nZ(w364) );
	vdp_sr_bit g327 (.D(w381), .C2(HCLK2), .C1(HCLK1), .Q(w905), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g328 (.D(w425), .Q(w394), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g329 (.D(w394), .Q(w392), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g330 (.D(w392), .Q(w386), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g331 (.D(w390), .Q(w431), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g332 (.D(w431), .Q(w387), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g333 (.D(w432), .Q(w381), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g334 (.D(w1462), .Q(w378), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g335 (.A(w414), .nZ(w1548) );
	vdp_not g336 (.A(w414), .nZ(w383) );
	vdp_not g337 (.A(w414), .nZ(w363) );
	vdp_not g338 (.A(w416), .nZ(w1401) );
	vdp_not g339 (.A(w416), .nZ(w384) );
	vdp_not g340 (.A(w416), .nZ(w370) );
	vdp_not g341 (.A(w428), .nZ(w1550) );
	vdp_not g342 (.A(w428), .nZ(w371) );
	vdp_not g343 (.A(w428), .nZ(w1500) );
	vdp_not g344 (.A(w417), .nZ(w361) );
	vdp_not g345 (.A(w417), .nZ(w1551) );
	vdp_not g346 (.A(w417), .nZ(w1943) );
	vdp_not g347 (.A(w978), .nZ(w1397) );
	vdp_not g348 (.A(w392), .nZ(w372) );
	vdp_not g349 (.A(nSEL0_M3), .nZ(w375) );
	vdp_comp_str g350 (.A(w407), .Z(w1507), .nZ(w1508) );
	vdp_comp_str g351 (.A(w408), .Z(w351), .nZ(w352) );
	vdp_comp_str g352 (.A(w379), .Z(w1403), .nZ(w353) );
	vdp_comp_str g353 (.A(w380), .Z(w1505), .nZ(w1506) );
	vdp_comp_str g354 (.A(w433), .Z(w1503), .nZ(w1504) );
	vdp_comp_str g355 (.A(w433), .Z(w1501), .nZ(w1502) );
	vdp_comp_str g356 (.A(w430), .Z(w354), .nZ(w355) );
	vdp_comp_str g357 (.A(w430), .Z(w356), .nZ(w357) );
	vdp_comp_str g358 (.A(w473), .Z(w395), .nZ(w1400) );
	vdp_comp_str g359 (.A(w473), .Z(w1399), .nZ(w362) );
	vdp_comp_str g360 (.A(w424), .Z(w360), .nZ(w359) );
	vdp_comp_str g361 (.A(w424), .Z(w358), .nZ(w1398) );
	vdp_comp_str g362 (.A(w434), .Z(w344), .nZ(w343) );
	vdp_comp_str g363 (.A(w434), .Z(w347), .nZ(w346) );
	vdp_comp_we g364 (.A(nSEL0_M3), .Z(w345), .nZ(w349) );
	vdp_comp_we g365 (.A(w413), .Z(w6428), .nZ(w6429) );
	vdp_comp_we g366 (.A(w413), .Z(w396), .nZ(w397) );
	vdp_comp_we g367 (.A(w413), .Z(w389), .nZ(w388) );
	vdp_comp_we g368 (.A(w413), .Z(w366), .nZ(w1510) );
	vdp_comp_we g369 (.A(w418), .Z(w6432), .nZ(w6433) );
	vdp_comp_we g370 (.A(w376), .Z(w367), .nZ(w368) );
	vdp_comp_we g371 (.A(w411), .Z(w1509), .nZ(w369) );
	vdp_and g372 (.Z(w379), .B(HCLK1), .A(w378) );
	vdp_and g373 (.Z(w380), .B(HCLK1), .A(w381) );
	vdp_and g374 (.Z(w1462), .B(w387), .A(w385) );
	vdp_and g375 (.Z(w432), .B(w387), .A(w391) );
	vdp_nand g376 (.Z(w391), .B(w418), .A(w372) );
	vdp_nand g377 (.Z(w385), .B(w418), .A(w392) );
	vdp_and3 g378 (.Z(w418), .B(w404), .A(nSEL0_M3), .C(w405) );
	vdp_and3 g379 (.Z(w376), .B(w375), .A(w386), .C(VRAM128k) );
	vdp_not g380 (.A(VRAM128k), .nZ(w405) );
	vdp_sr_bit g381 (.D(w402), .C2(HCLK2), .C1(HCLK1), .Q(w401), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g382 (.D(w1379), .Q(w438), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g383 (.D(w1463), .C2(HCLK2), .C1(HCLK1), .Q(w464), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g384 (.A(w465), .nZ(w393) );
	vdp_fa g385 (.SUM(w426), .A(w464), .B(1'b0), .CI(w466) );
	vdp_not g386 (.A(w402), .nZ(w400) );
	vdp_not g387 (.A(M5), .nZ(w437) );
	vdp_not g388 (.A(w410), .nZ(w408) );
	vdp_not g389 (.A(w420), .nZ(w421) );
	vdp_not g390 (.A(w471), .nZ(w423) );
	vdp_not g391 (.A(w464), .nZ(w422) );
	vdp_slatch g392 (.Q(w458), .D(CD[1]), .C(w444), .nC(w399) );
	vdp_slatch g393 (.Q(w1450), .D(CD[1]), .C(w456), .nC(w429) );
	vdp_slatch g394 (.Q(w459), .D(CD[1]), .C(w442), .nC(w415) );
	vdp_slatch g395 (.Q(w460), .D(CD[1]), .C(w440), .nC(w412) );
	vdp_slatch g396 (.Q(w461), .D(CD[2]), .C(w444), .nC(w399) );
	vdp_slatch g397 (.Q(w463), .D(CD[2]), .C(w456), .nC(w429) );
	vdp_slatch g398 (.Q(w1449), .D(CD[2]), .E(w442), .nE(w415) );
	vdp_slatch g399 (.Q(w457), .D(CD[2]), .C(w440), .nC(w412) );
	vdp_slatch g400 (.Q(w449), .D(CD[3]), .C(w444), .nC(w399) );
	vdp_slatch g401 (.Q(w443), .D(CD[3]), .C(w456), .nC(w429) );
	vdp_slatch g402 (.Q(w447), .D(CD[3]), .C(w442), .nC(w415) );
	vdp_slatch g403 (.Q(w450), .D(CD[3]), .C(w440), .nC(w412) );
	vdp_comp_dff g404 (.D(w406), .C2(HCLK2), .C1(HCLK1), .Q(w402), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and g405 (.Z(w1379), .B(w400), .A(w401) );
	vdp_or g406 (.Z(w407), .B(w437), .A(w408) );
	vdp_or g407 (.Z(w411), .B(CA[0]), .A(nSEL0_M3) );
	vdp_and3 g408 (.Z(w414), .B(w465), .A(w422), .C(w471) );
	vdp_and3 g409 (.Z(w416), .B(w465), .A(w423), .C(w464) );
	vdp_and3 g410 (.Z(w417), .B(w422), .A(w423), .C(w465) );
	vdp_xor g411 (.Z(w419), .B(w469), .A(w468) );
	vdp_aon22 g412 (.Z(w413), .A1(w421), .A2(w469), .B1(w486), .B2(w420) );
	vdp_and3 g413 (.Z(w428), .B(w464), .A(w471), .C(w465) );
	vdp_comp_str g414 (.A(w473), .Z(w444), .nZ(w399) );
	vdp_comp_str g415 (.A(w424), .Z(w440), .nZ(w412) );
	vdp_comp_str g416 (.A(w433), .Z(w442), .nZ(w415) );
	vdp_comp_str g417 (.A(w430), .Z(w456), .nZ(w429) );
	vdp_nand g418 (.Z(w420), .B(w470), .A(w419) );
	vdp_and g419 (.Z(w1463), .B(w467), .A(w426) );
	vdp_aoi21 g420 (.Z(w410), .B(w409), .A1(HCLK1), .A2(w438) );
	vdp_nor g421 (.Z(w409), .B(M3), .A(w437) );
	vdp_nor g422 (.Z(w404), .B(CD[2]), .A(CD[3]) );
	vdp_not g423 (.A(w452), .nZ(w510) );
	vdp_not g424 (.A(w451), .nZ(w514) );
	vdp_nor g425 (.Z(w574), .A(w497), .B(w452) );
	vdp_or g426 (.A(w1378), .Z(w453), .B(w454) );
	vdp_comp_we g427 (.A(w550), .nZ(w445), .Z(w491) );
	vdp_aon22 g428 (.Z(w451), .A1(w491), .A2(CD[3]), .B1(w445), .B2(w455) );
	vdp_aon22 g429 (.Z(w513), .A1(w491), .A2(CD[0]), .B1(w445), .B2(w453) );
	vdp_aon22 g430 (.Z(w519), .A1(w491), .A2(w502), .B1(w445), .B2(w468) );
	vdp_aon22 g431 (.Z(w452), .A1(w491), .A2(CD[2]), .B1(w445), .B2(w498) );
	vdp_aon22 g432 (.Z(w516), .A1(w491), .A2(w496), .B1(w445), .B2(w469) );
	vdp_aon22 g433 (.Z(w497), .A1(w491), .A2(CD[1]), .B1(w445), .B2(w490) );
	vdp_and g434 (.Z(w509), .A(w489), .B(w488) );
	vdp_and g435 (.Z(w448), .A(w489), .B(w471) );
	vdp_and g436 (.Z(w1451), .A(w464), .B(w488) );
	vdp_and g437 (.Z(w446), .A(w464), .B(w471) );
	vdp_and g438 (.Z(w1380), .A(w467), .B(w484) );
	vdp_fa g439 (.SUM(w484), .A(w471), .B(w472), .CO(w466), .CI(w485) );
	vdp_sr_bit g440 (.D(w1380), .C2(HCLK2), .C1(HCLK1), .Q(w471), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g441 (.A(w487), .nZ(w1382) );
	vdp_not g442 (.A(w477), .nZ(w480) );
	vdp_and g443 (.Z(w472), .A(w546), .B(w1382) );
	vdp_and3 g444 (.Z(w430), .B(w478), .A(w477), .C(w481) );
	vdp_and3 g445 (.Z(w473), .B(w478), .A(w477), .C(w479) );
	vdp_xor g446 (.Z(w483), .A(w464), .B(w477) );
	vdp_not g447 (.A(w471), .nZ(w488) );
	vdp_not g448 (.A(w464), .nZ(w489) );
	vdp_not g449 (.A(w470), .nZ(w1381) );
	vdp_and5 g450 (.Z(w33), .A(w511), .B(w519), .C(w515), .D(w514), .E(w452) );
	vdp_and5 g451 (.Z(w32), .A(w511), .B(w516), .C(w515), .D(w514), .E(w452) );
	vdp_aon2222 g452 (.C2(w506), .B2(w505), .A2(w504), .C1(w1451), .B1(w448), .A1(w509), .Z(w454), .D2(w507), .D1(w446) );
	vdp_aon2222 g453 (.C2(w443), .B2(w447), .A2(w450), .C1(w1451), .B1(w448), .A1(w509), .Z(w455), .D2(w449), .D1(w446) );
	vdp_aon2222 g454 (.C2(w1393), .B2(w501), .A2(w1394), .C1(w1451), .B1(w448), .A1(w509), .Z(w468), .D2(w499), .D1(w446) );
	vdp_aon2222 g455 (.C2(w463), .B2(w1449), .A2(w457), .C1(w1451), .B1(w448), .A1(w509), .Z(w498), .D2(w461), .D1(w446) );
	vdp_aon2222 g456 (.C2(w1452), .B2(w495), .A2(w492), .C1(w1451), .B1(w448), .A1(w509), .Z(w469), .D2(w508), .D1(w446) );
	vdp_aon2222 g457 (.C2(w1450), .B2(w459), .A2(w460), .C1(w1451), .B1(w448), .A1(w509), .Z(w490), .D2(w458), .D1(w446) );
	vdp_nor g458 (.Z(w487), .A(w1381), .B(w419) );
	vdp_or g459 (.Z(w434), .B(w474), .A(w931) );
	vdp_cnt_bit g460 (.R(SYSRES), .Q(w477), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2), .CI(w475) );
	vdp_cnt_bit g461 (.R(SYSRES), .Q(w479), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2), .CI(w539), .CO(w475) );
	vdp_not g462 (.A(w479), .nZ(w481) );
	vdp_not g463 (.A(w1383), .nZ(w478) );
	vdp_and3 g464 (.Z(w424), .B(w478), .A(w480), .C(w481) );
	vdp_and3 g465 (.Z(w433), .B(w478), .A(w480), .C(w479) );
	vdp_xor g466 (.Z(w482), .A(w471), .B(w479) );
	vdp_fa g467 (.SUM(w1514), .A(w547), .B(w486), .CO(w485), .CI(1'b0) );
	vdp_and g468 (.Z(w547), .A(w487), .B(w546) );
	vdp_and g469 (.Z(w1392), .A(w467), .B(w1514) );
	vdp_sr_bit g470 (.D(w1392), .C2(HCLK2), .C1(HCLK1), .Q(w486), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g471 (.A(w1390), .nZ(w532) );
	vdp_comp_str g472 (.A(w424), .Z(w526), .nZ(w503) );
	vdp_comp_str g473 (.A(w433), .Z(w534), .nZ(w493) );
	vdp_comp_str g474 (.A(w430), .Z(w533), .nZ(w500) );
	vdp_comp_str g475 (.A(w473), .Z(w535), .nZ(w494) );
	vdp_slatch g476 (.Q(w508), .D(w496), .C(w535), .nC(w494) );
	vdp_slatch g477 (.Q(w1452), .D(w496), .C(w533), .nC(w500) );
	vdp_slatch g478 (.Q(w495), .D(w496), .C(w534), .nC(w493) );
	vdp_slatch g479 (.Q(w492), .D(w496), .C(w526), .nC(w503) );
	vdp_slatch g480 (.Q(w499), .D(w502), .C(w535), .nC(w494) );
	vdp_slatch g481 (.Q(w1393), .D(w502), .C(w533), .nC(w500) );
	vdp_slatch g482 (.Q(w501), .D(w502), .C(w534), .nC(w493) );
	vdp_slatch g483 (.Q(w1394), .D(w502), .C(w526), .nC(w503) );
	vdp_slatch g484 (.Q(w507), .D(CD[0]), .C(w535), .nC(w494) );
	vdp_slatch g485 (.Q(w506), .D(CD[0]), .C(w533), .nC(w500) );
	vdp_slatch g486 (.Q(w505), .D(CD[0]), .C(w534), .nC(w493) );
	vdp_slatch g487 (.Q(w504), .D(CD[0]), .C(w526), .nC(w503) );
	vdp_and5 g488 (.Z(w1434), .A(w511), .B(w519), .C(w514), .D(w497), .E(w510) );
	vdp_and5 g489 (.Z(w1435), .A(w511), .B(w516), .C(w514), .D(w497), .E(w510) );
	vdp_not g490 (.A(M5), .nZ(w1378) );
	vdp_not g491 (.A(w497), .nZ(w515) );
	vdp_not g492 (.A(w512), .nZ(w511) );
	vdp_oai21 g493 (.A1(w550), .Z(w512), .A2(w546), .B(w513) );
	vdp_and3 g494 (.Z(w537), .B(w546), .A(w470), .C(w486) );
	vdp_nor g495 (.Z(w1391), .A(w536), .B(w486) );
	vdp_nor g496 (.Z(w544), .A(w483), .B(w482) );
	vdp_aoi21 g497 (.A1(DCLK1), .Z(w1383), .A2(w474), .B(w538) );
	vdp_comb1 g498 (.Z(w1390), .C1(w546), .B(w548), .C2(w1391), .A(HCLK1) );
	vdp_not g499 (.A(w524), .nZ(w517) );
	vdp_not g500 (.A(w1454), .nZ(w518) );
	vdp_not g501 (.A(VRAM128k), .nZ(w522) );
	vdp_not g502 (.A(w521), .nZ(w118) );
	vdp_not g503 (.A(w1455), .nZ(w119) );
	vdp_not g504 (.A(w1456), .nZ(w520) );
	vdp_not g505 (.A(VRAMA[0]), .nZ(w1457) );
	vdp_not g506 (.A(w528), .nZ(w527) );
	vdp_not g507 (.A(w464), .nZ(w571) );
	vdp_not g508 (.A(w471), .nZ(w573) );
	vdp_not g509 (.A(w549), .nZ(w570) );
	vdp_not g510 (.A(nSEL0_M3), .nZ(w569) );
	vdp_not g511 (.A(VRAM128k), .nZ(w1461) );
	vdp_not g512 (.A(w486), .nZ(w565) );
	vdp_not g513 (.A(SYSRES), .nZ(w467) );
	vdp_not g514 (.A(FIFO_EMPTY), .nZ(w1385) );
	vdp_not g515 (.A(w561), .nZ(w1384) );
	vdp_not g516 (.A(w545), .nZ(w560) );
	vdp_not g517 (.A(w538), .nZ(w542) );
	vdp_not g518 (.A(w542), .nZ(w543) );
	vdp_sr_bit g519 (.D(w1386), .C2(HCLK2), .C1(HCLK1), .Q(w546), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g520 (.D(w1389), .Q(w550), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_slatch g521 (.Q(w425), .D(VRAMA[0]), .C(w560), .nC(w545) );
	vdp_and g522 (.A(w30), .Z(w1386), .B(w1385) );
	vdp_and g523 (.A(w1384), .Z(w465), .B(w3) );
	vdp_and g524 (.A(w3), .Z(w545), .B(HCLK1) );
	vdp_and g525 (.A(FIFO_EMPTY), .Z(w561), .B(w552) );
	vdp_and g526 (.A(w553), .Z(w31), .B(FIFO_EMPTY) );
	vdp_and g527 (.A(w553), .B(w537) );
	vdp_or g528 (.A(w541), .Z(w539), .B(w474) );
	vdp_or g529 (.A(w543), .Z(w904), .B(1'b0) );
	vdp_or g530 (.A(SYSRES), .Z(w563), .B(w1007) );
	vdp_and g531 (.A(w546), .Z(w1387), .B(DMA_BUSY) );
	vdp_and g532 (.A(w574), .Z(w470), .B(w1460) );
	vdp_and g533 (.A(w1461), .Z(w1460), .B(nSEL0_M3) );
	vdp_or g534 (.A(w537), .Z(w568), .B(w536) );
	vdp_or g535 (.A(DMA_BUSY), .Z(w1458), .B(w531) );
	vdp_or g536 (.A(DMA_BUSY), .Z(w1459), .B(w530) );
	vdp_and g537 (.A(M5), .Z(w549), .B(REG_BUS[0]) );
	vdp_or g538 (.A(w519), .Z(w523), .B(w522) );
	vdp_and g539 (.A(w516), .Z(w1453), .B(VRAM128k) );
	vdp_aon22 g540 (.Z(w496), .A2(w1458), .B1(w569), .B2(w549), .A1(nSEL0_M3) );
	vdp_aon22 g541 (.Z(w502), .A2(w1459), .B1(w570), .B2(w569), .A1(nSEL0_M3) );
	vdp_and3 g542 (.A(w30), .Z(w1389), .B(w31), .C(w1388) );
	vdp_rs_ff g543 (.Q(w1388), .R(w563), .S(w1387) );
	vdp_oai21 g544 (.A1(VRAMA[0]), .Z(w528), .A2(VRAM128k), .B(w555) );
	vdp_oai21 g545 (.A1(VRAM128k), .Z(w1456), .A2(w1457), .B(w555) );
	vdp_aoi21 g546 (.A1(w516), .Z(w1455), .A2(w525), .B(w527) );
	vdp_aoi21 g547 (.A1(w519), .Z(w521), .A2(w525), .B(w520) );
	vdp_aoi21 g548 (.A1(w525), .Z(w1454), .A2(w523), .B(w555) );
	vdp_aoi21 g549 (.A1(w525), .Z(w524), .A2(w1453), .B(w555) );
	vdp_and4 g550 (.A(w511), .Z(w525), .B(w515), .C(w510), .D(w514) );
	vdp_not g551 (.A(w599), .nZ(w1377) );
	vdp_not g552 (.A(w611), .nZ(w610) );
	vdp_and3 g553 (.A(w565), .Z(w566), .B(w601), .C(w610) );
	vdp_and3 g554 (.A(w573), .Z(w587), .B(w575), .C(w571) );
	vdp_and3 g555 (.A(w471), .Z(w591), .B(w575), .C(w571) );
	vdp_and3 g556 (.A(w573), .Z(w579), .B(w575), .C(w464) );
	vdp_and3 g557 (.A(w471), .Z(w583), .B(w575), .C(w464) );
	vdp_or g558 (.A(w567), .Z(w598), .B(w600) );
	vdp_or g559 (.A(w567), .Z(w604), .B(w608) );
	vdp_or g560 (.A(w632), .Z(w757), .B(w607) );
	vdp_and3 g561 (.Z(w553), .B(DMA_BUSY), .A(w631), .C(w606) );
	vdp_or3 g562 (.Z(w556), .B(w550), .A(w555), .C(w605) );
	vdp_and g563 (.A(w558), .Z(w474), .B(w557) );
	vdp_and g564 (.A(w546), .Z(w575), .B(w565) );
	vdp_bufif0 g565 (.A(w559), .Z(VRAMA[8]), .nE(w612) );
	vdp_aoi221 g566 (.Z(w599), .A2(w566), .B1(FIFO_EMPTY), .B2(w544), .A1(w544), .C(SYSRES) );
	vdp_aon33 g567 (.Z(FIFO_FULL), .A2(w544), .B1(w1494), .B2(w544), .A1(w609), .A3(w1494), .B3(w562) );
	vdp_not g568 (.A(w568), .nZ(w1406) );
	vdp_comp_str g569 (.A(w532), .Z(w1407), .nZ(w594) );
	vdp_not g570 (.A(w591), .nZ(w593) );
	vdp_comp_str g571 (.A(w433), .Z(w1409), .nZ(w1408) );
	vdp_not g572 (.A(w568), .nZ(w813) );
	vdp_comp_str g573 (.A(w532), .Z(w595), .nZ(w596) );
	vdp_not g574 (.A(w548), .nZ(w612) );
	vdp_not g575 (.A(w591), .nZ(w1495) );
	vdp_comp_str g576 (.A(w433), .Z(w1410), .nZ(w592) );
	vdp_not g577 (.A(w587), .nZ(w586) );
	vdp_comp_str g578 (.A(w424), .Z(w1411), .nZ(w1499) );
	vdp_not g579 (.A(w587), .nZ(w588) );
	vdp_comp_str g580 (.A(w473), .Z(w1412), .nZ(w585) );
	vdp_comp_str g581 (.A(w424), .Z(w589), .nZ(w590) );
	vdp_not g582 (.A(w579), .nZ(w576) );
	vdp_comp_str g583 (.A(w430), .Z(w577), .nZ(w578) );
	vdp_not g584 (.A(w579), .nZ(w812) );
	vdp_comp_str g585 (.A(w430), .Z(w1497), .nZ(w1498) );
	vdp_not g586 (.A(w583), .nZ(w580) );
	vdp_comp_str g587 (.A(w473), .Z(w581), .nZ(w582) );
	vdp_not g588 (.A(w583), .nZ(w1496) );
	vdp_sr_bit g589 (.D(w1377), .Q(FIFO_EMPTY), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g590 (.D(w601), .Q(w611), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g591 (.D(w546), .Q(w601), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g592 (.D(FIFO_FULL), .Q(w609), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g593 (.D(w539), .Q(w562), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_not g594 (.A(SYSRES), .nZ(w1494) );
	vdp_not g595 (.A(w1464), .nZ(w605) );
	vdp_sr_bit g596 (.D(w558), .Q(w557), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g597 (.D(w551), .C2(HCLK2), .C1(HCLK1), .Q(w1007), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_dlatch_inv g598 (.D(w558), .C(HCLK2), .Q(w1464), .nC(nHCLK2) );
	vdp_slatch g599 (.D(w622), .C(w577), .nC(w578), .nQ(w6448) );
	vdp_slatch g600 (.D(REG_BUS[7]), .C(w1497), .nC(w1498), .nQ(w6449) );
	vdp_slatch g601 (.D(w622), .C(w581), .nC(w582), .nQ(w6468) );
	vdp_slatch g602 (.D(REG_BUS[7]), .C(w1412), .nC(w585), .nQ(w6466) );
	vdp_slatch g603 (.D(w622), .C(w1411), .nC(w1499), .nQ(w6482) );
	vdp_slatch g604 (.D(REG_BUS[7]), .C(w589), .nC(w590), .nQ(w6484) );
	vdp_slatch g605 (.D(w622), .C(w1410), .nC(w592), .nQ(w6502) );
	vdp_slatch g606 (.D(REG_BUS[7]), .C(w1409), .nC(w1408), .nQ(w6500) );
	vdp_slatch g607 (.D(VRAMA[9]), .C(w1407), .nC(w594), .nQ(w6516) );
	vdp_slatch g608 (.D(VRAMA[7]), .C(w595), .nC(w596), .nQ(w6517) );
	vdp_notif0 g609 (.nZ(VRAMA[7]), .nE(w813), .A(w6517) );
	vdp_notif0 g610 (.nZ(VRAMA[9]), .nE(w1406), .A(w6516) );
	vdp_notif0 g611 (.nZ(VRAMA[7]), .nE(w593), .A(w6500) );
	vdp_notif0 g612 (.nZ(VRAMA[9]), .nE(w1495), .A(w6502) );
	vdp_notif0 g613 (.nZ(VRAMA[7]), .nE(w588), .A(w6484) );
	vdp_notif0 g614 (.nZ(VRAMA[9]), .nE(w580), .A(w6468) );
	vdp_notif0 g615 (.nZ(VRAMA[7]), .nE(w1496), .A(w6466) );
	vdp_notif0 g616 (.nZ(VRAMA[9]), .nE(w586), .A(w6482) );
	vdp_notif0 g617 (.nZ(VRAMA[9]), .nE(w576), .A(w6448) );
	vdp_notif0 g618 (.nZ(VRAMA[7]), .nE(w812), .A(w6449) );
	vdp_bufif0 g619 (.A(w622), .Z(VRAMA[9]), .nE(w612) );
	vdp_bufif0 g620 (.A(REG_BUS[7]), .Z(VRAMA[7]), .nE(w612) );
	vdp_bufif0 g621 (.A(w615), .Z(VRAMA[8]), .nE(w1445) );
	vdp_bufif0 g622 (.A(w615), .Z(CA[8]), .nE(w815) );
	vdp_bufif0 g623 (.A(w614), .Z(VRAMA[7]), .nE(w1443) );
	vdp_bufif0 g624 (.A(w614), .Z(CA[7]), .nE(w814) );
	vdp_slatch g625 (.Q(w631), .D(REG_BUS[7]), .nQ(w629), .C(w1541), .nC(w1542) );
	vdp_not g626 (.A(REG_BUS[0]), .nZ(w627) );
	vdp_not g627 (.A(REG_BUS[7]), .nZ(w633) );
	vdp_and3 g628 (.Z(w632), .B(w606), .A(w629), .C(DMA_BUSY) );
	vdp_nand g629 (.A(w625), .Z(w653), .B(w626) );
	vdp_cnt_bit_load g630 (.D(REG_BUS[0]), .nL(w1544), .L(w1554), .R(1'b0), .Q(w615), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w598), .CO(w619) );
	vdp_cnt_bit_load g631 (.D(REG_BUS[7]), .nL(w1376), .L(w762), .R(1'b0), .Q(w614), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w617), .CO(w600) );
	vdp_cnt_bit_load g632 (.D(w627), .nL(w1543), .L(w774), .R(1'b0), .Q(w625), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w604), .CO(w624) );
	vdp_cnt_bit_load g633 (.D(w633), .nL(w750), .L(w751), .R(1'b0), .Q(w628), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w630), .CO(w608) );
	vdp_slatch g634 (.D(w641), .C(w577), .nC(w578), .nQ(w6447) );
	vdp_slatch g635 (.D(REG_BUS[6]), .C(w1497), .nC(w1498), .nQ(w6450) );
	vdp_slatch g636 (.D(w641), .C(w581), .nC(w582), .nQ(w6467) );
	vdp_slatch g637 (.D(REG_BUS[6]), .C(w1412), .nC(w585), .nQ(w6465) );
	vdp_slatch g638 (.D(w641), .C(w1411), .nC(w1499), .nQ(w6481) );
	vdp_slatch g639 (.D(REG_BUS[6]), .C(w589), .nC(w590), .nQ(w6483) );
	vdp_slatch g640 (.D(w641), .C(w1410), .nC(w592), .nQ(w6501) );
	vdp_slatch g641 (.D(REG_BUS[6]), .C(w1409), .nC(w1408), .nQ(w6499) );
	vdp_slatch g642 (.D(VRAMA[10]), .C(w1407), .nC(w594), .nQ(w6515) );
	vdp_slatch g643 (.D(VRAMA[6]), .C(w595), .nC(w596), .nQ(w6518) );
	vdp_notif0 g644 (.nZ(VRAMA[6]), .nE(w813), .A(w6518) );
	vdp_notif0 g645 (.nZ(VRAMA[10]), .nE(w1406), .A(w6515) );
	vdp_notif0 g646 (.nZ(VRAMA[6]), .nE(w593), .A(w6499) );
	vdp_notif0 g647 (.nZ(VRAMA[10]), .nE(w1495), .A(w6501) );
	vdp_notif0 g648 (.nZ(VRAMA[6]), .nE(w588), .A(w6483) );
	vdp_notif0 g649 (.nZ(VRAMA[10]), .nE(w580), .A(w6467) );
	vdp_notif0 g650 (.nZ(VRAMA[6]), .nE(w1496), .A(w6465) );
	vdp_notif0 g651 (.nZ(VRAMA[10]), .nE(w586), .A(w6481) );
	vdp_notif0 g652 (.nZ(VRAMA[10]), .nE(w576), .A(w6447) );
	vdp_notif0 g653 (.nZ(VRAMA[6]), .nE(w812), .A(w6450) );
	vdp_bufif0 g654 (.A(w641), .Z(VRAMA[10]), .nE(w612) );
	vdp_bufif0 g655 (.A(REG_BUS[6]), .Z(VRAMA[6]), .nE(w1446) );
	vdp_bufif0 g656 (.A(w613), .Z(VRAMA[9]), .nE(w1445) );
	vdp_bufif0 g657 (.A(w613), .Z(CA[9]), .nE(w815) );
	vdp_bufif0 g658 (.A(w635), .Z(VRAMA[6]), .nE(w1443) );
	vdp_bufif0 g659 (.A(w635), .Z(CA[6]), .nE(w814) );
	vdp_slatch g660 (.Q(w648), .D(REG_BUS[6]), .nQ(w606), .C(w1541), .nC(w1542) );
	vdp_not g661 (.A(REG_BUS[1]), .nZ(w644) );
	vdp_not g662 (.A(REG_BUS[6]), .nZ(w646) );
	vdp_and3 g663 (.Z(w607), .B(DMA_BUSY), .A(w648), .C(w629) );
	vdp_cnt_bit_load g664 (.D(REG_BUS[1]), .nL(w1544), .L(w1554), .R(1'b0), .Q(w613), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w619), .CO(w637) );
	vdp_cnt_bit_load g665 (.D(REG_BUS[6]), .nL(w1376), .L(w762), .R(1'b0), .Q(w635), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w636), .CO(w617) );
	vdp_cnt_bit_load g666 (.D(w644), .nL(w1543), .L(w774), .R(1'b0), .Q(w626), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w624), .CO(w643) );
	vdp_cnt_bit_load g667 (.D(w646), .nL(w750), .L(w751), .R(1'b0), .Q(w645), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w649), .CO(w630) );
	vdp_nand3 g668 (.Z(w652), .B(w645), .A(w651), .C(w628) );
	vdp_slatch g669 (.D(w671), .C(w577), .nC(w578), .nQ(w6446) );
	vdp_slatch g670 (.D(REG_BUS[5]), .C(w1497), .nC(w1498), .nQ(w6451) );
	vdp_slatch g671 (.D(w671), .C(w581), .nC(w582), .nQ(w6469) );
	vdp_slatch g672 (.D(REG_BUS[5]), .C(w1412), .nC(w585), .nQ(w6464) );
	vdp_slatch g673 (.D(w671), .C(w1411), .nC(w1499), .nQ(w6480) );
	vdp_slatch g674 (.D(w671), .C(w1410), .nC(w592), .nQ(w6503) );
	vdp_slatch g675 (.D(REG_BUS[5]), .C(w1409), .nC(w1408), .nQ(w6498) );
	vdp_slatch g676 (.D(VRAMA[11]), .C(w1407), .nC(w594), .nQ(w6514) );
	vdp_slatch g677 (.D(VRAMA[5]), .C(w595), .nC(w596), .nQ(w6519) );
	vdp_notif0 g678 (.nZ(VRAMA[5]), .nE(w813), .A(w6519) );
	vdp_notif0 g679 (.nZ(VRAMA[11]), .nE(w1406), .A(w6514) );
	vdp_notif0 g680 (.nZ(VRAMA[5]), .nE(w593), .A(w6498) );
	vdp_notif0 g681 (.nZ(VRAMA[11]), .nE(w1495), .A(w6503) );
	vdp_notif0 g682 (.nZ(VRAMA[5]), .nE(w588), .A(w6485) );
	vdp_notif0 g683 (.nZ(VRAMA[11]), .nE(w580), .A(w6469) );
	vdp_notif0 g684 (.nZ(VRAMA[5]), .nE(w1496), .A(w6464) );
	vdp_notif0 g685 (.nZ(VRAMA[11]), .nE(w586), .A(w6480) );
	vdp_notif0 g686 (.nZ(VRAMA[11]), .nE(w576), .A(w6446) );
	vdp_notif0 g687 (.nZ(VRAMA[5]), .nE(w812), .A(w6451) );
	vdp_bufif0 g688 (.A(w671), .Z(VRAMA[11]), .nE(w612) );
	vdp_bufif0 g689 (.A(REG_BUS[5]), .Z(VRAMA[5]), .nE(w1446) );
	vdp_bufif0 g690 (.A(w634), .Z(VRAMA[10]), .nE(w1445) );
	vdp_bufif0 g691 (.A(w634), .Z(CA[10]), .nE(w815) );
	vdp_bufif0 g692 (.A(w665), .Z(VRAMA[5]), .nE(w1443) );
	vdp_bufif0 g693 (.A(w665), .Z(CA[5]), .nE(w814) );
	vdp_slatch g694 (.Q(CA[18]), .D(REG_BUS[2]), .C(w1541), .nC(w1542) );
	vdp_not g695 (.A(REG_BUS[2]), .nZ(w659) );
	vdp_not g696 (.A(REG_BUS[5]), .nZ(w658) );
	vdp_and3 g697 (.Z(w552), .B(DMA_BUSY), .A(w648), .C(w631) );
	vdp_cnt_bit_load g698 (.D(REG_BUS[2]), .nL(w1544), .L(w1554), .R(1'b0), .Q(w634), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w637), .CO(w668) );
	vdp_cnt_bit_load g699 (.D(REG_BUS[5]), .nL(w1376), .L(w762), .R(1'b0), .Q(w665), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w664), .CO(w636) );
	vdp_cnt_bit_load g700 (.D(w659), .nL(w1543), .L(w774), .R(1'b0), .Q(w650), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w643), .CO(w660) );
	vdp_cnt_bit_load g701 (.D(w658), .nL(w750), .L(w751), .R(1'b0), .Q(w651), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w655), .CO(w649) );
	vdp_nand3 g702 (.Z(w663), .B(w661), .A(w662), .C(w650) );
	vdp_slatch g703 (.D(w677), .C(w577), .nC(w578), .nQ(w6445) );
	vdp_slatch g704 (.D(REG_BUS[4]), .C(w1497), .nC(w1498), .nQ(w6452) );
	vdp_slatch g705 (.D(w677), .C(w581), .nC(w582), .nQ(w6470) );
	vdp_slatch g706 (.D(REG_BUS[4]), .C(w1412), .nC(w585), .nQ(w6463) );
	vdp_slatch g707 (.D(w677), .C(w1411), .nC(w1499), .nQ(w6479) );
	vdp_slatch g708 (.D(w677), .C(w1410), .nC(w592), .nQ(w6504) );
	vdp_slatch g709 (.D(REG_BUS[4]), .C(w1409), .nC(w1408), .nQ(w6497) );
	vdp_slatch g710 (.D(VRAMA[12]), .C(w1407), .nC(w594), .nQ(w6513) );
	vdp_slatch g711 (.D(VRAMA[4]), .C(w595), .nC(w596), .nQ(w6520) );
	vdp_notif0 g712 (.nZ(VRAMA[4]), .nE(w813), .A(w6520) );
	vdp_notif0 g713 (.nZ(VRAMA[12]), .nE(w1406), .A(w6513) );
	vdp_notif0 g714 (.nZ(VRAMA[4]), .nE(w593), .A(w6497) );
	vdp_notif0 g715 (.nZ(VRAMA[12]), .nE(w1495), .A(w6504) );
	vdp_notif0 g716 (.nZ(VRAMA[4]), .nE(w588), .A(w6486) );
	vdp_notif0 g717 (.nZ(VRAMA[12]), .nE(w580), .A(w6470) );
	vdp_notif0 g718 (.nZ(VRAMA[4]), .nE(w1496), .A(w6463) );
	vdp_notif0 g719 (.nZ(VRAMA[12]), .nE(w586), .A(w6479) );
	vdp_notif0 g720 (.nZ(VRAMA[12]), .nE(w576), .A(w6445) );
	vdp_notif0 g721 (.nZ(VRAMA[4]), .nE(w812), .A(w6452) );
	vdp_bufif0 g722 (.A(w677), .Z(VRAMA[12]), .nE(w612) );
	vdp_bufif0 g723 (.A(REG_BUS[4]), .Z(VRAMA[4]), .nE(w1446) );
	vdp_bufif0 g724 (.A(w667), .Z(VRAMA[11]), .nE(w1445) );
	vdp_bufif0 g725 (.A(w667), .Z(CA[11]), .nE(w815) );
	vdp_bufif0 g726 (.A(w678), .Z(VRAMA[4]), .nE(w1443) );
	vdp_bufif0 g727 (.A(w678), .Z(CA[4]), .nE(w814) );
	vdp_slatch g728 (.Q(CA[19]), .D(REG_BUS[3]), .C(w1541), .nC(w1542) );
	vdp_not g729 (.A(REG_BUS[3]), .nZ(w679) );
	vdp_not g730 (.A(REG_BUS[4]), .nZ(w681) );
	vdp_and g731 (.Z(w551), .B(w657), .A(w689) );
	vdp_cnt_bit_load g732 (.D(REG_BUS[3]), .nL(w1544), .L(w1554), .R(1'b0), .Q(w667), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w668), .CO(w673) );
	vdp_cnt_bit_load g733 (.D(REG_BUS[4]), .nL(w1376), .L(w762), .R(1'b0), .Q(w678), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w683), .CO(w664) );
	vdp_cnt_bit_load g734 (.D(w679), .nL(w1543), .L(w774), .R(1'b0), .Q(w661), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w660), .CO(w684) );
	vdp_cnt_bit_load g735 (.D(w681), .nL(w750), .L(w751), .R(1'b0), .Q(w687), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w688), .CO(w655) );
	vdp_nor3 g736 (.Z(w657), .B(w663), .A(w686), .C(w653) );
	vdp_slatch g737 (.D(w694), .C(w577), .nC(w578), .nQ(w6444) );
	vdp_slatch g738 (.D(REG_BUS[3]), .C(w1497), .nC(w1498), .nQ(w6453) );
	vdp_slatch g739 (.D(w694), .C(w581), .nC(w582), .nQ(w6471) );
	vdp_slatch g740 (.D(REG_BUS[3]), .C(w1412), .nC(w585), .nQ(w6462) );
	vdp_slatch g741 (.D(w694), .C(w1411), .nC(w1499), .nQ(w6478) );
	vdp_slatch g742 (.D(REG_BUS[3]), .C(w589), .nC(w590), .nQ(w6488) );
	vdp_slatch g743 (.D(w694), .C(w1410), .nC(w592), .nQ(w6506) );
	vdp_slatch g744 (.D(REG_BUS[3]), .C(w1409), .nC(w1408), .nQ(w6496) );
	vdp_slatch g745 (.D(VRAMA[13]), .C(w1407), .nC(w594), .nQ(w6512) );
	vdp_slatch g746 (.D(VRAMA[3]), .C(w595), .nC(w596), .nQ(w6521) );
	vdp_notif0 g747 (.nZ(VRAMA[3]), .nE(w813), .A(w6521) );
	vdp_notif0 g748 (.nZ(VRAMA[13]), .nE(w1406), .A(w6512) );
	vdp_notif0 g749 (.nZ(VRAMA[3]), .nE(w593), .A(w6496) );
	vdp_notif0 g750 (.nZ(VRAMA[13]), .nE(w1495), .A(w6506) );
	vdp_notif0 g751 (.nZ(VRAMA[3]), .nE(w588), .A(w6488) );
	vdp_notif0 g752 (.nZ(VRAMA[13]), .nE(w580), .A(w6471) );
	vdp_notif0 g753 (.nZ(VRAMA[3]), .nE(w1496), .A(w6462) );
	vdp_notif0 g754 (.nZ(VRAMA[13]), .nE(w586), .A(w6478) );
	vdp_notif0 g755 (.nZ(VRAMA[13]), .nE(w576), .A(w6444) );
	vdp_notif0 g756 (.nZ(VRAMA[3]), .nE(w812), .A(w6453) );
	vdp_bufif0 g757 (.A(w694), .Z(VRAMA[13]), .nE(w612) );
	vdp_bufif0 g758 (.A(REG_BUS[3]), .Z(VRAMA[3]), .nE(w1446) );
	vdp_bufif0 g759 (.A(w672), .Z(VRAMA[12]), .nE(w1445) );
	vdp_bufif0 g760 (.A(w672), .Z(CA[12]), .nE(w815) );
	vdp_bufif0 g761 (.A(w702), .Z(VRAMA[3]), .nE(w1443) );
	vdp_bufif0 g762 (.A(w702), .Z(CA[3]), .nE(w814) );
	vdp_slatch g763 (.Q(w708), .D(REG_BUS[4]), .C(w1541), .nC(w1542) );
	vdp_not g764 (.A(REG_BUS[4]), .nZ(w696) );
	vdp_not g765 (.A(REG_BUS[3]), .nZ(w697) );
	vdp_cnt_bit_load g766 (.D(REG_BUS[4]), .nL(w1544), .L(w1554), .R(1'b0), .Q(w672), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w673), .CO(w693) );
	vdp_cnt_bit_load g767 (.D(REG_BUS[3]), .nL(w1376), .L(w762), .R(1'b0), .Q(w702), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w691), .CO(w683) );
	vdp_cnt_bit_load g768 (.D(w696), .nL(w1543), .L(w774), .R(1'b0), .Q(w662), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w684), .CO(w701) );
	vdp_cnt_bit_load g769 (.D(w697), .nL(w750), .L(w751), .R(1'b0), .Q(w706), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w698), .CO(w688) );
	vdp_nor3 g770 (.Z(w689), .B(w707), .A(w705), .C(w652) );
	vdp_bufif0 g771 (.A(w708), .Z(CA[20]), .nE(w748) );
	vdp_slatch g772 (.D(w712), .C(w577), .nC(w578), .nQ(w6443) );
	vdp_slatch g773 (.D(REG_BUS[2]), .C(w1497), .nC(w1498), .nQ(w6454) );
	vdp_slatch g774 (.D(w712), .C(w581), .nC(w582), .nQ(w6472) );
	vdp_slatch g775 (.D(REG_BUS[2]), .C(w1412), .nC(w585), .nQ(w6461) );
	vdp_slatch g776 (.D(w712), .C(w1411), .nC(w1499), .nQ(w6477) );
	vdp_slatch g777 (.D(REG_BUS[2]), .C(w589), .nC(w590), .nQ(w6487) );
	vdp_slatch g778 (.D(w712), .C(w1410), .nC(w592), .nQ(w6505) );
	vdp_slatch g779 (.D(REG_BUS[2]), .C(w1409), .nC(w1408), .nQ(w6495) );
	vdp_slatch g780 (.D(VRAMA[14]), .C(w1407), .nC(w594), .nQ(w6511) );
	vdp_slatch g781 (.D(VRAMA[2]), .nC(w596), .C(w595), .nQ(w6522) );
	vdp_notif0 g782 (.nZ(VRAMA[2]), .nE(w813), .A(w6522) );
	vdp_notif0 g783 (.nZ(VRAMA[14]), .nE(w1406), .A(w6511) );
	vdp_notif0 g784 (.nZ(VRAMA[2]), .nE(w593), .A(w6495) );
	vdp_notif0 g785 (.nZ(VRAMA[14]), .nE(w1495), .A(w6505) );
	vdp_notif0 g786 (.nZ(VRAMA[2]), .nE(w588), .A(w6487) );
	vdp_notif0 g787 (.nZ(VRAMA[14]), .nE(w580), .A(w6472) );
	vdp_notif0 g788 (.nZ(VRAMA[2]), .nE(w1496), .A(w6461) );
	vdp_notif0 g789 (.nZ(VRAMA[14]), .nE(w586), .A(w6477) );
	vdp_notif0 g790 (.nZ(VRAMA[14]), .nE(w576), .A(w6443) );
	vdp_notif0 g791 (.nZ(VRAMA[2]), .nE(w812), .A(w6454) );
	vdp_bufif0 g792 (.A(w712), .Z(VRAMA[14]), .nE(w1444) );
	vdp_bufif0 g793 (.A(REG_BUS[2]), .Z(VRAMA[2]), .nE(w1446) );
	vdp_bufif0 g794 (.A(w692), .Z(VRAMA[13]), .nE(w1445) );
	vdp_bufif0 g795 (.A(w692), .Z(CA[13]), .nE(w815) );
	vdp_bufif0 g796 (.A(w713), .Z(VRAMA[2]), .nE(w1443) );
	vdp_bufif0 g797 (.A(w713), .Z(CA[2]), .nE(w814) );
	vdp_slatch g798 (.Q(w718), .D(REG_BUS[5]), .C(w1541), .nC(w1542) );
	vdp_not g799 (.A(REG_BUS[5]), .nZ(w714) );
	vdp_not g800 (.A(REG_BUS[2]), .nZ(w715) );
	vdp_cnt_bit_load g801 (.D(REG_BUS[5]), .nL(w1544), .L(w1554), .R(1'b0), .Q(w692), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w693), .CO(w724) );
	vdp_cnt_bit_load g802 (.D(REG_BUS[2]), .nL(w1376), .L(w762), .R(1'b0), .Q(w713), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w723), .CO(w691) );
	vdp_cnt_bit_load g803 (.D(w714), .nL(w1543), .L(w774), .R(1'b0), .Q(w722), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w701), .CO(w716) );
	vdp_cnt_bit_load g804 (.D(w715), .nL(w750), .L(w751), .R(1'b0), .Q(w720), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w726), .CO(w698) );
	vdp_nand3 g805 (.Z(w707), .B(w706), .A(w720), .C(w687) );
	vdp_bufif0 g806 (.A(w718), .Z(CA[21]), .nE(w748) );
	vdp_slatch g807 (.D(w731), .C(w577), .nC(w578), .nQ(w6442) );
	vdp_slatch g808 (.D(REG_BUS[1]), .C(w1497), .nC(w1498), .nQ(w6455) );
	vdp_slatch g809 (.D(w731), .C(w581), .nC(w582), .nQ(w6474) );
	vdp_slatch g810 (.D(REG_BUS[1]), .C(w1412), .nC(w585), .nQ(w6460) );
	vdp_slatch g811 (.D(w731), .C(w1411), .nC(w1499), .nQ(w6476) );
	vdp_slatch g812 (.D(REG_BUS[1]), .C(w589), .nC(w590), .nQ(w6490) );
	vdp_slatch g813 (.D(w731), .C(w1410), .nC(w592), .nQ(w6507) );
	vdp_slatch g814 (.D(REG_BUS[1]), .C(w1409), .nC(w1408), .nQ(w6494) );
	vdp_slatch g815 (.D(VRAMA[15]), .C(w1407), .nC(w594), .nQ(w6510) );
	vdp_slatch g816 (.D(VRAMA[1]), .C(w595), .nC(w596), .nQ(w6523) );
	vdp_notif0 g817 (.nZ(VRAMA[1]), .nE(w813), .A(w6523) );
	vdp_notif0 g818 (.nZ(VRAMA[15]), .nE(w1406), .A(w6510) );
	vdp_notif0 g819 (.nZ(VRAMA[1]), .nE(w593), .A(w6494) );
	vdp_notif0 g820 (.nZ(VRAMA[15]), .nE(w1495), .A(w6507) );
	vdp_notif0 g821 (.nZ(VRAMA[1]), .nE(w588), .A(w6490) );
	vdp_notif0 g822 (.nZ(VRAMA[15]), .nE(w580), .A(w6474) );
	vdp_notif0 g823 (.nZ(VRAMA[1]), .nE(w1496), .A(w6460) );
	vdp_notif0 g824 (.nZ(VRAMA[15]), .nE(w586), .A(w6476) );
	vdp_notif0 g825 (.nZ(VRAMA[15]), .nE(w576), .A(w6442) );
	vdp_notif0 g826 (.nZ(VRAMA[1]), .nE(w812), .A(w6455) );
	vdp_bufif0 g827 (.A(w731), .Z(VRAMA[15]), .nE(w1444) );
	vdp_bufif0 g828 (.A(REG_BUS[1]), .Z(VRAMA[1]), .nE(w1446) );
	vdp_bufif0 g829 (.A(w709), .Z(VRAMA[14]), .nE(w1445) );
	vdp_bufif0 g830 (.A(w709), .Z(CA[14]), .nE(w815) );
	vdp_bufif0 g831 (.A(w733), .Z(VRAMA[1]), .nE(w1443) );
	vdp_bufif0 g832 (.A(w733), .Z(CA[1]), .nE(w814) );
	vdp_slatch g833 (.Q(w1447), .D(REG_BUS[1]), .C(w1541), .nC(w1542) );
	vdp_not g834 (.A(REG_BUS[6]), .nZ(w736) );
	vdp_not g835 (.A(REG_BUS[1]), .nZ(w739) );
	vdp_cnt_bit_load g836 (.D(REG_BUS[6]), .nL(w1544), .L(w1554), .R(1'b0), .Q(w709), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w724), .CO(w740) );
	vdp_cnt_bit_load g837 (.D(REG_BUS[1]), .nL(w1376), .L(w762), .R(1'b0), .Q(w733), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w741), .CO(w723) );
	vdp_cnt_bit_load g838 (.D(w736), .nL(w1543), .L(w774), .R(1'b0), .Q(w721), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w716), .CO(w734) );
	vdp_cnt_bit_load g839 (.D(w739), .nL(w750), .L(w751), .R(1'b0), .Q(w738), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w737), .CO(w726) );
	vdp_nand3 g840 (.Z(w686), .B(w721), .A(w722), .C(w735) );
	vdp_bufif0 g841 (.A(w1447), .Z(CA[17]), .nE(w748) );
	vdp_slatch g842 (.nQ(w732), .D(w745), .C(w577), .nC(w578) );
	vdp_slatch g843 (.D(REG_BUS[0]), .C(w1497), .nC(w1498), .nQ(w6456) );
	vdp_slatch g844 (.D(w745), .C(w581), .nC(w582), .nQ(w6473) );
	vdp_slatch g845 (.D(REG_BUS[0]), .C(w1412), .nC(w585), .nQ(w6459) );
	vdp_slatch g846 (.D(w745), .C(w1411), .nC(w1499), .nQ(w6475) );
	vdp_slatch g847 (.D(REG_BUS[0]), .C(w589), .nC(w590), .nQ(w6489) );
	vdp_slatch g848 (.D(w745), .C(w1410), .nC(w592), .nQ(w6508) );
	vdp_slatch g849 (.D(REG_BUS[0]), .C(w1409), .nC(w1408), .nQ(w6493) );
	vdp_slatch g850 (.D(VRAMA[16]), .C(w1407), .nC(w594), .nQ(w6509) );
	vdp_slatch g851 (.Q(w6524), .D(VRAMA[0]), .C(w595), .nC(w596) );
	vdp_notif0 g852 (.nZ(VRAMA[0]), .nE(w813), .A(w6524) );
	vdp_notif0 g853 (.nZ(VRAMA[16]), .nE(w1406), .A(w6509) );
	vdp_notif0 g854 (.nZ(VRAMA[0]), .nE(w593), .A(w6493) );
	vdp_notif0 g855 (.nZ(VRAMA[16]), .nE(w1495), .A(w6508) );
	vdp_notif0 g856 (.nZ(VRAMA[0]), .nE(w588), .A(w6489) );
	vdp_notif0 g857 (.nZ(VRAMA[16]), .nE(w580), .A(w6473) );
	vdp_notif0 g858 (.nZ(VRAMA[0]), .nE(w1496), .A(w6459) );
	vdp_notif0 g859 (.nZ(VRAMA[16]), .nE(w586), .A(w6475) );
	vdp_notif0 g860 (.A(w732), .nZ(VRAMA[16]), .nE(w576) );
	vdp_notif0 g861 (.nZ(VRAMA[0]), .nE(w812), .A(w6456) );
	vdp_bufif0 g862 (.A(w745), .Z(VRAMA[16]), .nE(w1444) );
	vdp_bufif0 g863 (.A(REG_BUS[0]), .Z(VRAMA[0]), .nE(w1446) );
	vdp_bufif0 g864 (.A(w727), .Z(VRAMA[15]), .nE(w1445) );
	vdp_bufif0 g865 (.A(w727), .Z(CA[15]), .nE(w815) );
	vdp_bufif0 g866 (.A(w755), .Z(VRAMA[0]), .nE(w1443) );
	vdp_bufif0 g867 (.A(w755), .Z(CA[0]), .nE(w814) );
	vdp_slatch g868 (.Q(w746), .D(REG_BUS[0]), .C(w1541), .nC(w1542) );
	vdp_not g869 (.A(REG_BUS[7]), .nZ(w1545) );
	vdp_not g870 (.A(REG_BUS[0]), .nZ(w1414) );
	vdp_cnt_bit_load g871 (.D(REG_BUS[7]), .nL(w1544), .L(w1554), .R(1'b0), .Q(w727), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w740) );
	vdp_cnt_bit_load g872 (.D(REG_BUS[0]), .nL(w1376), .L(w762), .R(1'b0), .Q(w755), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w753), .CO(w741) );
	vdp_cnt_bit_load g873 (.D(w1545), .nL(w1543), .L(w774), .R(1'b0), .Q(w735), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w734) );
	vdp_cnt_bit_load g874 (.D(w1414), .nL(w750), .L(w751), .R(1'b0), .Q(w1413), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w753), .CO(w737) );
	vdp_nand3 g875 (.Z(w705), .B(w738), .A(w556), .C(w1369) );
	vdp_bufif0 g876 (.A(w746), .Z(CA[16]), .nE(w748) );
	vdp_slatch g877 (.D(VRAMA[8]), .C(w595), .nC(w596), .nQ(w6525) );
	vdp_slatch g878 (.D(w559), .C(w1409), .nC(w1408), .nQ(w6492) );
	vdp_slatch g879 (.D(w559), .C(w589), .nC(w590), .nQ(w6491) );
	vdp_slatch g880 (.D(w559), .C(w1412), .nC(w585), .nQ(w6458) );
	vdp_slatch g881 (.D(w559), .C(w1497), .nC(w1498), .nQ(w6457) );
	vdp_notif0 g882 (.nZ(VRAMA[8]), .nE(w812), .A(w6457) );
	vdp_notif0 g883 (.nZ(VRAMA[8]), .nE(w1496), .A(w6458) );
	vdp_notif0 g884 (.nZ(VRAMA[8]), .nE(w588), .A(w6491) );
	vdp_notif0 g885 (.nZ(VRAMA[8]), .nE(w593), .A(w6492) );
	vdp_notif0 g886 (.nZ(VRAMA[8]), .nE(w813), .A(w6525) );
	vdp_bufif0 g887 (.A(w746), .Z(VRAMA[16]), .nE(w1445) );
	vdp_not g888 (.A(w1405), .nZ(w1444) );
	vdp_not g889 (.A(w548), .nZ(w1446) );
	vdp_not g890 (.A(w760), .nZ(w1445) );
	vdp_not g891 (.A(w757), .nZ(w815) );
	vdp_not g892 (.A(w760), .nZ(w1443) );
	vdp_not g893 (.A(w757), .nZ(w814) );
	vdp_not g894 (.A(w757), .nZ(w748) );
	vdp_not g895 (.A(w1413), .nZ(w1369) );
	vdp_not g896 (.A(w749), .nZ(w1375) );
	vdp_not g897 (.A(M5), .nZ(w770) );
	vdp_and4 g898 (.Z(w766), .B(w641), .A(w775), .D(w559), .C(w776) );
	vdp_and4 g899 (.Z(w767), .B(w641), .A(w775), .D(w778), .C(w622) );
	vdp_and4 g900 (.B(w780), .A(w756), .D(w778), .C(w776), .Z(w769) );
	vdp_and4 g901 (.B(w780), .A(w756), .D(w559), .C(w776), .Z(w768) );
	vdp_and4 g902 (.Z(w759), .B(w776), .A(w559), .D(w781), .C(w641) );
	vdp_and4 g903 (.Z(w771), .B(w622), .A(w778), .D(w756), .C(w780) );
	vdp_and4 g904 (.Z(w758), .B(w622), .A(w559), .D(w781), .C(w641) );
	vdp_and4 g905 (.B(w784), .A(M5), .D(w671), .C(w785), .Z(w775) );
	vdp_comp_str g906 (.A(w787), .Z(w1541), .nZ(w1542) );
	vdp_comp_we g907 (.A(w1418), .Z(w1554), .nZ(w1544) );
	vdp_comp_we g908 (.A(w761), .Z(w762), .nZ(w1376) );
	vdp_comp_we g909 (.A(w788), .Z(w774), .nZ(w1543) );
	vdp_comp_we g910 (.A(w789), .Z(w751), .nZ(w750) );
	vdp_and g911 (.Z(w567), .B(w556), .A(w749) );
	vdp_and g912 (.Z(w753), .B(w556), .A(w1375) );
	vdp_or g913 (.Z(w787), .B(w758), .A(SYSRES) );
	vdp_or g914 (.Z(w761), .B(w759), .A(SYSRES) );
	vdp_or g915 (.Z(w1405), .B(w770), .A(w548) );
	vdp_or g916 (.B(w768), .A(SYSRES), .Z(w763) );
	vdp_or g917 (.B(w769), .A(SYSRES), .Z(w764) );
	vdp_or g918 (.Z(w765), .B(w767), .A(SYSRES) );
	vdp_or g919 (.Z(w1421), .B(w766), .A(SYSRES) );
	vdp_or g920 (.B(w1415), .A(SYSRES), .Z(w792) );
	vdp_and4 g921 (.B(w641), .A(w777), .D(w559), .C(w622), .Z(w799) );
	vdp_or g922 (.B(w799), .A(SYSRES), .Z(w811) );
	vdp_and4 g923 (.B(w780), .A(w781), .D(w778), .C(w622), .Z(w798) );
	vdp_or g924 (.B(w798), .A(SYSRES), .Z(w793) );
	vdp_and4 g925 (.B(w780), .A(w781), .D(w559), .C(w776), .Z(w797) );
	vdp_or g926 (.B(w797), .A(SYSRES), .Z(w794) );
	vdp_and4 g927 (.B(w780), .A(w781), .D(w778), .C(w776), .Z(w1416) );
	vdp_or g928 (.B(w1416), .A(SYSRES), .Z(w779) );
	vdp_and4 g929 (.B(w641), .A(w777), .D(w778), .C(w622), .Z(w796) );
	vdp_or g930 (.B(w796), .A(SYSRES), .Z(w157) );
	vdp_and4 g931 (.B(w641), .A(w777), .D(w559), .C(w776), .Z(w795) );
	vdp_or g932 (.B(w795), .A(SYSRES), .Z(w156) );
	vdp_or g933 (.B(w800), .A(SYSRES), .Z(w791) );
	vdp_and4 g934 (.B(w641), .A(w777), .D(w778), .C(w776), .Z(w1415) );
	vdp_or g935 (.B(w801), .A(SYSRES), .Z(w790) );
	vdp_and4 g936 (.B(w780), .A(w777), .D(w559), .C(w622), .Z(w800) );
	vdp_and4 g937 (.B(w780), .A(w777), .D(w778), .C(w622), .Z(w801) );
	vdp_and4 g938 (.B(w776), .A(w559), .D(w777), .C(w780), .Z(w803) );
	vdp_or g939 (.B(w803), .A(SYSRES), .Z(w1091) );
	vdp_and4 g940 (.B(w776), .A(w778), .D(w777), .C(w780), .Z(w1417) );
	vdp_or g941 (.B(w1417), .A(SYSRES), .Z(w1129) );
	vdp_and4 g942 (.B(w776), .A(w778), .D(w775), .C(w641), .Z(w802) );
	vdp_or g943 (.B(w802), .A(SYSRES), .Z(w1092) );
	vdp_and4 g944 (.B(w622), .A(w778), .D(w781), .C(w641), .Z(w804) );
	vdp_or g945 (.B(w804), .A(SYSRES), .Z(w1418) );
	vdp_and4 g946 (.B(w622), .A(w559), .D(w775), .C(w780), .Z(w1419) );
	vdp_or g947 (.B(w1419), .A(SYSRES), .Z(w1053) );
	vdp_and4 g948 (.B(w776), .A(w778), .D(w781), .C(w641), .Z(w805) );
	vdp_or g949 (.B(w805), .A(SYSRES), .Z(w788) );
	vdp_and4 g950 (.B(w622), .A(w559), .D(w781), .C(w780), .Z(w806) );
	vdp_or g951 (.B(w806), .A(SYSRES), .Z(w789) );
	vdp_and4 g952 (.B(w622), .A(w559), .D(w775), .C(w641), .Z(w807) );
	vdp_or g953 (.B(w807), .A(SYSRES), .Z(w808) );
	vdp_and4 g954 (.B(w786), .A(w784), .D(M5), .C(w677), .Z(w781) );
	vdp_and3 g955 (.B(w785), .A(w784), .C(w671), .Z(w756) );
	vdp_and3 g956 (.B(w786), .A(w784), .C(w785), .Z(w777) );
	vdp_or g957 (.Z(w809), .B(w810), .A(w6427) );
	vdp_and g958 (.B(w783), .A(HCLK1), .Z(w784) );
	vdp_dlatch_inv g959 (.D(w782), .C(DCLK2), .nQ(w810), .nC(nDCLK2) );
	vdp_dlatch_inv g960 (.D(w6426), .C(HCLK2), .nQ(w783), .nC(nHCLK2) );
	vdp_not g961 (.A(w677), .nZ(w785) );
	vdp_not g962 (.A(w671), .nZ(w786) );
	vdp_not g963 (.A(w622), .nZ(w776) );
	vdp_not g964 (.A(w641), .nZ(w780) );
	vdp_not g965 (.A(w559), .nZ(w778) );
	vdp_slatch g966 (.D(REG_BUS[5]), .C(w589), .nC(w590), .nQ(w6485) );
	vdp_slatch g967 (.D(REG_BUS[4]), .C(w589), .nC(w590), .nQ(w6486) );
	vdp_sr_bit g968 (.D(w810), .C2(DCLK2), .C1(DCLK1), .Q(w6427), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_dlatch_inv g969 (.D(w809), .C(DCLK1), .nQ(w6426), .nC(nDCLK1) );
	vdp_comp_str g970 (.A(w847), .Z(w817), .nZ(w825) );
	vdp_fa g971 (.SUM(w844), .A(REG_BUS[6]), .B(w1518), .CO(w846), .CI(w842) );
	vdp_fa g972 (.SUM(w840), .A(REG_BUS[5]), .B(w841), .CO(w842), .CI(w839) );
	vdp_fa g973 (.SUM(w837), .A(REG_BUS[4]), .B(w838), .CO(w839), .CI(w834) );
	vdp_fa g974 (.SUM(w833), .A(REG_BUS[3]), .B(w836), .CO(w834), .CI(w831) );
	vdp_fa g975 (.SUM(w829), .A(REG_BUS[2]), .B(w830), .CO(w831), .CI(w828) );
	vdp_fa g976 (.SUM(w6430), .A(REG_BUS[1]), .B(w827), .CO(w828), .CI(w824) );
	vdp_fa g977 (.SUM(w6431), .A(REG_BUS[0]), .B(w821), .CO(w824), .CI(w819) );
	vdp_fa g978 (.SUM(w1420), .A(REG_BUS[7]), .B(w1517), .CO(w848), .CI(w846) );
	vdp_slatch g979 (.Q(w845), .D(DB[7]), .C(w817), .nC(w825) );
	vdp_aon22 g980 (.Z(w1528), .A1(w845), .A2(w816), .B1(w822), .B2(w1420) );
	vdp_slatch g981 (.Q(w843), .D(DB[6]), .C(w817), .nC(w825) );
	vdp_aon22 g982 (.Z(w1529), .A1(w843), .A2(w816), .B1(w822), .B2(w844) );
	vdp_slatch g983 (.Q(w1469), .D(DB[5]), .C(w817), .nC(w825) );
	vdp_aon22 g984 (.Z(w1530), .A1(w1469), .A2(w816), .B1(w822), .B2(w840) );
	vdp_slatch g985 (.Q(w835), .D(DB[4]), .C(w817), .nC(w825) );
	vdp_aon22 g986 (.Z(w1531), .A1(w835), .A2(w816), .B1(w822), .B2(w837) );
	vdp_slatch g987 (.Q(w832), .D(DB[3]), .C(w817), .nC(w825) );
	vdp_aon22 g988 (.Z(w1532), .A1(w832), .A2(w816), .B1(w822), .B2(w833) );
	vdp_slatch g989 (.Q(w826), .D(DB[2]), .C(w817), .nC(w825) );
	vdp_aon22 g990 (.Z(w1533), .A1(w826), .A2(w816), .B1(w822), .B2(w829) );
	vdp_slatch g991 (.Q(w823), .D(DB[1]), .C(w817), .nC(w825) );
	vdp_aon22 g992 (.Z(w1534), .A1(w823), .A2(w816), .B1(w822), .B2(w6430) );
	vdp_slatch g993 (.Q(w818), .D(DB[0]), .C(w817), .nC(w825) );
	vdp_aon22 g994 (.Z(w1535), .A1(w818), .A2(w816), .B1(w822), .B2(w6431) );
	vdp_dff g995 (.Q(REG_BUS[0]), .R(SYSRES), .C(w850), .D(w1535) );
	vdp_slatch g996 (.Q(w821), .D(REG_BUS[0]), .C(w849), .nC(w820) );
	vdp_dff g997 (.Q(REG_BUS[1]), .R(SYSRES), .D(w1534), .C(w850) );
	vdp_slatch g998 (.Q(w827), .D(REG_BUS[1]), .C(w849), .nC(w820) );
	vdp_dff g999 (.Q(REG_BUS[2]), .R(SYSRES), .C(w850), .D(w1533) );
	vdp_slatch g1000 (.Q(w830), .D(REG_BUS[2]), .C(w849), .nC(w820) );
	vdp_dff g1001 (.Q(REG_BUS[3]), .R(SYSRES), .D(w1532), .C(w850) );
	vdp_slatch g1002 (.Q(w836), .D(REG_BUS[3]), .C(w849), .nC(w820) );
	vdp_dff g1003 (.Q(REG_BUS[4]), .R(SYSRES), .C(w850), .D(w1531) );
	vdp_slatch g1004 (.Q(w838), .D(REG_BUS[4]), .C(w849), .nC(w820) );
	vdp_dff g1005 (.Q(REG_BUS[5]), .R(SYSRES), .C(w850), .D(w1530) );
	vdp_slatch g1006 (.Q(w841), .D(REG_BUS[5]), .C(w849), .nC(w820) );
	vdp_dff g1007 (.Q(REG_BUS[6]), .R(SYSRES), .C(w850), .D(w1529) );
	vdp_slatch g1008 (.Q(w1518), .D(REG_BUS[6]), .C(w849), .nC(w820) );
	vdp_dff g1009 (.Q(REG_BUS[7]), .R(SYSRES), .D(w1528), .C(w850) );
	vdp_slatch g1010 (.Q(w1517), .D(REG_BUS[7]), .C(w849), .nC(w820) );
	vdp_comp_str g1011 (.A(w808), .Z(w849), .nZ(w820) );
	vdp_comp_we g1012 (.A(w851), .Z(w816), .nZ(w822) );
	vdp_dff g1013 (.Q(w745), .R(w855), .C(w850), .D(w1519) );
	vdp_dff g1014 (.Q(w731), .R(w855), .C(w850), .D(w1520) );
	vdp_dff g1015 (.Q(w712), .R(w855), .C(w850), .D(w1521) );
	vdp_dff g1016 (.Q(w694), .R(SYSRES), .C(w850), .D(w1522) );
	vdp_dff g1017 (.Q(w677), .R(SYSRES), .C(w850), .D(w1523) );
	vdp_dff g1018 (.Q(w671), .R(SYSRES), .C(w850), .D(w1524) );
	vdp_dff g1019 (.Q(w641), .R(SYSRES), .C(w850), .D(w1525) );
	vdp_dff g1020 (.Q(w622), .R(SYSRES), .C(w850), .D(w1526) );
	vdp_dff g1021 (.Q(w559), .R(SYSRES), .C(w850), .D(w1527) );
	vdp_not g1022 (.A(w877), .nZ(w850) );
	vdp_or g1023 (.Z(w855), .B(SYSRES), .A(w819) );
	vdp_not g1024 (.A(M5), .nZ(w819) );
	vdp_slatch g1025 (.Q(w874), .D(w259), .C(w887), .nC(w865) );
	vdp_aon22 g1026 (.Z(w1527), .A1(w878), .A2(w885), .B1(w852), .B2(w876) );
	vdp_slatch g1027 (.Q(w878), .D(w226), .C(w887), .nC(w865) );
	vdp_comp_str g1028 (.A(w892), .Z(w887), .nZ(w865) );
	vdp_comp_we g1029 (.A(w851), .Z(w885), .nZ(w852) );
	vdp_ha g1030 (.SUM(w876), .A(w559), .B(w848), .CO(w873) );
	vdp_slatch g1031 (.Q(w872), .D(w233), .C(w887), .nC(w865) );
	vdp_aon22 g1032 (.Z(w1526), .A1(w874), .A2(w885), .B1(w852), .B2(w875) );
	vdp_ha g1033 (.SUM(w875), .A(w622), .B(w873), .CO(w1538) );
	vdp_slatch g1034 (.Q(w870), .D(w267), .C(w887), .nC(w865) );
	vdp_aon22 g1035 (.Z(w1525), .A1(w872), .A2(w885), .B1(w852), .B2(w871) );
	vdp_ha g1036 (.SUM(w871), .A(w641), .B(w1538), .CO(w869) );
	vdp_slatch g1037 (.Q(w867), .D(w888), .C(w887), .nC(w865) );
	vdp_aon22 g1038 (.Z(w1524), .A1(w870), .A2(w885), .B1(w852), .B2(w868) );
	vdp_ha g1039 (.SUM(w868), .A(w671), .B(w869), .CO(w1537) );
	vdp_slatch g1040 (.Q(w864), .D(w275), .C(w887), .nC(w865) );
	vdp_aon22 g1041 (.Z(w1523), .A1(w867), .A2(w885), .B1(w852), .B2(w866) );
	vdp_ha g1042 (.SUM(w866), .A(w677), .B(w1537), .CO(w863) );
	vdp_aon22 g1043 (.Z(w1522), .A1(w864), .A2(w885), .B1(w852), .B2(w861) );
	vdp_ha g1044 (.SUM(w861), .A(w694), .B(w863), .CO(w862) );
	vdp_comp_str g1045 (.A(w886), .Z(w884), .nZ(w854) );
	vdp_aon22 g1046 (.Z(w1521), .A1(w860), .A2(w885), .B1(w852), .B2(w1536) );
	vdp_ha g1047 (.SUM(w1536), .A(w712), .B(w862), .CO(w857) );
	vdp_slatch_r g1048 (.Q(w860), .D(DB[0]), .R(w855), .C(w884), .nC(w854) );
	vdp_slatch_r g1049 (.Q(w859), .D(DB[1]), .R(w855), .C(w884), .nC(w854) );
	vdp_aon22 g1050 (.Z(w1520), .A1(w859), .A2(w885), .B1(w852), .B2(w858) );
	vdp_ha g1051 (.SUM(w858), .A(w731), .B(w857), .CO(w856) );
	vdp_slatch_r g1052 (.Q(w853), .D(DB[2]), .R(w855), .C(w884), .nC(w854) );
	vdp_aon22 g1053 (.Z(w1519), .A1(w853), .A2(w885), .B1(w852), .B2(w1468) );
	vdp_ha g1054 (.SUM(w1468), .A(w745), .B(w856) );
	vdp_and3 g1055 (.C(w881), .A(w879), .B(w880), .Z(w883) );
	vdp_sr_bit g1056 (.D(w1427), .C2(HCLK2), .C1(HCLK1), .nQ(w95), .nC1(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1057 (.D(w900), .Q(w1427), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK2), .nC1(nHCLK1) );
	vdp_not g1058 (.A(w942), .nZ(w902) );
	vdp_not g1059 (.A(CD[2]), .nZ(w1428) );
	vdp_not g1060 (.A(CD[3]), .nZ(w913) );
	vdp_not g1061 (.A(w879), .nZ(w914) );
	vdp_not g1062 (.A(w911), .nZ(w919) );
	vdp_not g1063 (.A(CD[0]), .nZ(w897) );
	vdp_not g1064 (.A(w552), .nZ(w908) );
	vdp_not g1065 (.A(w932), .nZ(w922) );
	vdp_not g1066 (.A(w1429), .nZ(w925) );
	vdp_not g1067 (.A(w923), .nZ(w893) );
	vdp_slatch g1068 (.Q(CD[1]), .D(w890), .C(w891), .nC(w903) );
	vdp_slatch g1069 (.Q(CD[0]), .D(w250), .C(w891), .nC(w903) );
	vdp_comp_str g1070 (.A(w892), .Z(w891), .nZ(w903) );
	vdp_dlatch_inv g1071 (.D(w558), .C(DCLK1), .nQ(w923), .nC(nDCLK1) );
	vdp_dlatch_inv g1072 (.D(w922), .C(DCLK1), .nQ(w921), .nC(nDCLK1) );
	vdp_dlatch_inv g1073 (.D(w934), .C(DCLK2), .nQ(w932), .nC(nDCLK2) );
	vdp_dlatch_inv g1074 (.D(w939), .C(DCLK1), .nQ(w934), .nC(nDCLK1) );
	vdp_slatch g1075 (.Q(w939), .D(w899), .C(DCLK2), .nC(nDCLK2) );
	vdp_slatch g1076 (.Q(w899), .D(w933), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g1077 (.D(w548), .C(HCLK1), .nQ(w898), .nC(nHCLK1) );
	vdp_rs_ff g1078 (.nQ(w895), .R(w941), .S(w940), .Q(w906) );
	vdp_rs_ff g1079 (.Q(w918), .R(w916), .S(w896) );
	vdp_and3 g1080 (.C(w390), .A(CD[3]), .B(w1428), .Z(w901) );
	vdp_and3 g1081 (.C(w913), .A(CD[2]), .B(w390), .Z(w94) );
	vdp_comp_dff g1082 (.D(w917), .C2(HCLK2), .C1(HCLK1), .Q(w910), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_comp_dff g1083 (.D(w907), .C2(HCLK2), .C1(HCLK1), .Q(w909), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g1084 (.C(w30), .A(w906), .B(FIFO_EMPTY), .Z(w907) );
	vdp_and g1085 (.A(DB[7]), .B(w886), .Z(w889) );
	vdp_and g1086 (.A(w898), .B(w939), .Z(w851) );
	vdp_and g1087 (.A(w909), .B(w908), .Z(w536) );
	vdp_and g1088 (.A(w552), .B(w909), .Z(w555) );
	vdp_and g1089 (.A(w910), .B(w908), .Z(w920) );
	vdp_and g1090 (.A(w552), .B(w910), .Z(w760) );
	vdp_or g1091 (.A(w910), .B(w930), .Z(w916) );
	vdp_or g1092 (.A(w910), .B(w536), .Z(w390) );
	vdp_or g1093 (.A(w552), .B(w418), .Z(w938) );
	vdp_aoi21 g1094 (.A1(w921), .B(SYSRES), .Z(w1429), .A2(w922) );
	vdp_or3 g1095 (.C(w894), .A(w915), .B(w883), .Z(w896) );
	vdp_or3 g1096 (.C(w555), .A(w920), .B(w550), .Z(w548) );
	vdp_or5 g1097 (.C(w904), .A(w893), .B(w548), .Z(w877), .D(w892), .E(w886) );
	vdp_nand3 g1098 (.C(w882), .A(w919), .B(w928), .Z(w782) );
	vdp_2a3oi g1099 (.A1(w881), .B(w935), .Z(w929), .A2(w928), .C(w880) );
	vdp_nand g1100 (.A(CD[1]), .B(w897), .Z(w911) );
	vdp_nor g1101 (.A(w899), .B(w934), .Z(w882) );
	vdp_and4 g1102 (.C(w895), .A(FIFO_EMPTY), .B(w30), .Z(w917), .D(w918) );
	vdp_nor5 g1103 (.C(CD[0]), .A(CD[4]), .B(w929), .Z(w894), .D(CD[1]), .E(w914) );
	vdp_and g1104 (.A(w552), .B(CD[4]), .Z(w915) );
	vdp_not g1105 (.A(w541), .nZ(w1486) );
	vdp_not g1106 (.A(w1486), .nZ(w977) );
	vdp_not g1107 (.A(w958), .nZ(w997) );
	vdp_not g1108 (.A(w934), .nZ(w1436) );
	vdp_not g1109 (.A(w939), .nZ(w979) );
	vdp_not g1110 (.A(w982), .nZ(w892) );
	vdp_not g1111 (.A(nSEL0_M3), .nZ(w912) );
	vdp_not g1112 (.A(w967), .nZ(w975) );
	vdp_not g1113 (.A(M5), .nZ(w881) );
	vdp_rs_ff g1114 (.Q(w928), .R(w926), .S(w892) );
	vdp_rs_ff g1115 (.Q(w880), .R(w926), .S(w1002) );
	vdp_rs_ff g1116 (.Q(w935), .R(w926), .S(w886) );
	vdp_rs_ff g1117 (.nQ(w937), .R(w936), .S(w905) );
	vdp_rs_ff g1118 (.Q(w999), .R(w925), .S(w931) );
	vdp_rs_ff g1119 (.Q(w531), .R(w925), .S(w992) );
	vdp_rs_ff g1120 (.Q(w530), .R(w925), .S(w949) );
	vdp_or g1121 (.A(w949), .B(w992), .Z(w1001) );
	vdp_and g1122 (.A(w999), .B(w879), .Z(w538) );
	vdp_and g1123 (.A(w998), .B(w999), .Z(w541) );
	vdp_and g1124 (.A(w979), .B(w1436), .Z(w879) );
	vdp_and g1125 (.A(w979), .B(w932), .Z(w998) );
	vdp_and g1126 (.A(w934), .B(w932), .Z(w965) );
	vdp_and g1127 (.A(w910), .B(w938), .Z(w940) );
	vdp_and g1128 (.A(w961), .B(w950), .Z(w382) );
	vdp_and g1129 (.A(w912), .B(w847), .Z(w1009) );
	vdp_and g1130 (.A(w985), .B(w984), .Z(w931) );
	vdp_or g1131 (.A(w909), .B(w930), .Z(w941) );
	vdp_or g1132 (.A(w978), .B(w981), .Z(w924) );
	vdp_or g1133 (.A(SYSRES), .B(w879), .Z(w936) );
	vdp_or g1134 (.A(SYSRES), .B(w939), .Z(w1005) );
	vdp_or g1135 (.A(w934), .B(w933), .Z(w1000) );
	vdp_or g1136 (.A(w961), .B(w985), .Z(w1006) );
	vdp_or g1137 (.A(w927), .B(SYSRES), .Z(w971) );
	vdp_or g1138 (.A(SYSRES), .B(w966), .Z(w1011) );
	vdp_or g1139 (.A(SYSRES), .B(w965), .Z(w926) );
	vdp_and g1140 (.A(w942), .B(w901), .Z(w116) );
	vdp_and g1141 (.A(w901), .B(w902), .Z(w93) );
	vdp_and g1142 (.A(w879), .B(w973), .Z(w1010) );
	vdp_nand g1143 (.A(w382), .B(w937), .Z(w990) );
	vdp_nor g1144 (.A(FIFO_FULL), .B(w977), .Z(w991) );
	vdp_or5 g1145 (.C(w892), .A(w976), .B(w989), .Z(w988), .D(w847), .E(w993) );
	vdp_or3 g1146 (.C(w980), .A(w961), .B(w377), .Z(w981) );
	vdp_nor g1147 (.A(w94), .B(w901), .Z(w900) );
	vdp_and3 g1148 (.C(w1012), .A(w1008), .B(w963), .Z(w983) );
	vdp_or4 g1149 (.C(w931), .A(w886), .B(w960), .Z(w927), .D(w382) );
	vdp_and4 g1150 (.C(w986), .A(w985), .B(w968), .Z(w847), .D(w1008) );
	vdp_aoi21 g1151 (.A1(w879), .B(SYSRES), .Z(w967), .A2(w974) );
	vdp_aoi21 g1152 (.A1(w847), .B(w983), .Z(w982), .A2(nSEL0_M3) );
	vdp_or5 g1153 (.C(w382), .A(w960), .B(w886), .Z(w966), .D(w931), .E(w892) );
	vdp_and5 g1154 (.C(w972), .A(M5), .B(w1008), .Z(w886), .D(w986), .E(w985) );
	vdp_not g1155 (.A(CA[7]), .nZ(w954) );
	vdp_not g1156 (.A(w985), .nZ(w962) );
	vdp_not g1157 (.A(w962), .nZ(w947) );
	vdp_not g1158 (.A(w961), .nZ(w946) );
	vdp_not g1159 (.A(w946), .nZ(w945) );
	vdp_slatch g1160 (.Q(w987), .D(w948), .nC(w945), .C(w946) );
	vdp_slatch g1161 (.Q(w1008), .D(w948), .nC(w947), .C(w962), .nQ(w984) );
	vdp_rs_ff g1162 (.Q(w969), .R(w965), .S(w971) );
	vdp_rs_ff g1163 (.Q(w973), .R(w1011), .S(w1009), .nQ(w974) );
	vdp_rs_ff g1164 (.Q(w1012), .R(w975), .S(w1010), .nQ(w986) );
	vdp_rs_ff g1165 (.Q(w972), .R(w970), .S(w1425), .nQ(w968) );
	vdp_slatch_r g1166 (.Q(CD[4]), .D(DB[6]), .C(w964), .nC(w944), .R(w855) );
	vdp_slatch_r g1167 (.Q(CD[3]), .D(DB[5]), .R(w855), .C(w964), .nC(w944) );
	vdp_slatch_r g1168 (.Q(CD[2]), .D(DB[4]), .R(w855), .C(w964), .nC(w944) );
	vdp_comp_str g1169 (.A(w886), .Z(w964), .nZ(w944) );
	vdp_not g1170 (.A(w1426), .nZ(w970) );
	vdp_aoi21 g1171 (.A1(w879), .B(SYSRES), .Z(w1426), .A2(w969) );
	vdp_and4 g1172 (.C(w911), .A(M5), .B(w928), .Z(w1425), .D(w879) );
	vdp_and g1173 (.A(w961), .B(w987), .Z(w1002) );
	vdp_rs_ff g1174 (.nQ(w1004), .R(w1003), .S(w1002) );
	vdp_rs_ff g1175 (.Q(w933), .R(w1005), .S(w1006) );
	vdp_not g1176 (.A(w948), .nZ(w1539) );
	vdp_not g1177 (.A(CA[2]), .nZ(w1035) );
	vdp_not g1178 (.A(CA[3]), .nZ(w1036) );
	vdp_aon22 g1179 (.Z(w948), .A1(CA[0]), .A2(w1060), .B1(nSEL0_M3), .B2(CA[1]) );
	vdp_and4 g1180 (.C(w953), .A(w954), .B(CA[6]), .Z(w996), .D(w952) );
	vdp_and4 g1181 (.C(w957), .A(w956), .B(CA[7]), .Z(w963), .D(w952) );
	vdp_and4 g1182 (.C(CA[3]), .A(w997), .B(w995), .Z(w980), .D(CA[9]) );
	vdp_and4 g1183 (.C(CA[2]), .A(w997), .B(w995), .Z(w373), .D(w1036) );
	vdp_and4 g1184 (.C(w958), .A(w1035), .B(CA[3]), .Z(w955), .D(w995) );
	vdp_or g1185 (.A(w996), .B(w373), .Z(w377) );
	vdp_and g1186 (.A(w931), .B(w991), .Z(w989) );
	vdp_and g1187 (.A(w981), .B(w990), .Z(w993) );
	vdp_and g1188 (.A(nSEL0_M3), .B(w988), .Z(w1026) );
	vdp_or g1189 (.A(SYSRES), .B(w905), .Z(w1003) );
	vdp_or g1190 (.A(w963), .B(w951), .Z(w985) );
	vdp_or g1191 (.A(SYSRES), .B(w1007), .Z(w930) );
	vdp_and3 g1192 (.C(w1034), .A(w886), .B(w1004), .Z(w976) );
	vdp_and3 g1193 (.C(w1037), .A(w1000), .B(w1160), .Z(w995) );
	vdp_and5 g1194 (.C(CA[2]), .A(w958), .B(CA[3]), .Z(w1031), .D(w1539), .E(w995) );
	vdp_and5 g1195 (.C(CA[2]), .A(w958), .B(w948), .Z(w1030), .D(CA[3]), .E(w995) );
	vdp_and5 g1196 (.C(w1035), .A(w1001), .B(w997), .Z(w959), .D(w1036), .E(w995) );
	vdp_and5 g1197 (.C(w1036), .A(w1035), .B(w1001), .Z(w951), .D(w958), .E(w995) );
	vdp_nor5 g1198 (.C(w1027), .A(w1030), .B(w1031), .Z(w1013), .D(w955), .E(w1026) );
	vdp_aon22 g1199 (.Z(w1023), .A1(w4), .A2(w1033), .B1(w34), .B2(nSEL0_M3) );
	vdp_aon22 g1200 (.Z(VPOS_80), .A1(w1016), .A2(VPOS[8]), .B1(w1021), .B2(VPOS[0]) );
	vdp_not g1201 (.A(w1016), .nZ(w1021) );
	vdp_not g1202 (.A(nSEL0_M3), .nZ(w1017) );
	vdp_not g1203 (.A(nSEL0_M3), .nZ(w1033) );
	vdp_not g1204 (.A(w1483), .nZ(w98) );
	vdp_not g1205 (.A(CA[6]), .nZ(w956) );
	vdp_not g1206 (.A(w1423), .nZ(nPSGWRITE) );
	vdp_not g1207 (.A(w948), .nZ(w950) );
	vdp_aoi21 g1208 (.A1(w949), .B(w1424), .Z(w1423), .A2(w955) );
	vdp_and4 g1209 (.C(w953), .A(w956), .B(CA[7]), .Z(w1422), .D(w952) );
	vdp_and4 g1210 (.C(w957), .A(w954), .B(CA[6]), .Z(w1424), .D(w952) );
	vdp_slatch g1211 (.Q(w100), .D(w953), .C(w1540), .nC(w1484) );
	vdp_comp_we g1212 (.A(PSG_Z80_CLK), .Z(w1540), .nZ(w1484) );
	vdp_and g1213 (.A(w44), .B(w1028), .Z(w1485) );
	vdp_and g1214 (.A(w948), .B(w961), .Z(w960) );
	vdp_or g1215 (.A(w959), .B(w1422), .Z(w961) );
	vdp_or g1216 (.A(w1027), .B(w1485), .Z(w1029) );
	vdp_or g1217 (.Z(w1022), .A(w35), .B(SYSRES) );
	vdp_and g1218 (.Z(V_INT_HAPPENED), .A(w55), .B(w1023) );
	vdp_rs_ff g1219 (.Q(w1019), .R(w1022), .S(V_INT_HAPPENED) );
	vdp_aoi221 g1220 (.Z(w1483), .A1(w97), .A2(1'b1), .B1(w1024), .B2(w1029), .C(w99) );
	vdp_aoi22 g1221 (.Z(w1014), .A1(w1020), .A2(w1017), .B1(nSEL0_M3), .B2(w1019) );
	vdp_comp_str g1222 (.Z(w1046), .A(w55), .nZ(w1047) );
	vdp_comp_str g1223 (.Z(w1072), .A(w1053), .nZ(w1073) );
	vdp_comp_str g1224 (.Z(w1084), .A(w1092), .nZ(w1085) );
	vdp_comp_str g1225 (.Z(w1081), .A(w1091), .nZ(w1080) );
	vdp_not g1226 (.A(w1090), .nZ(w1093) );
	vdp_not g1227 (.A(w1082), .nZ(w1095) );
	vdp_not g1228 (.A(w1079), .nZ(w1094) );
	vdp_not g1229 (.A(w1094), .nZ(w1059) );
	vdp_not g1230 (.A(nSEL0_M3), .nZ(w1060) );
	vdp_not g1231 (.A(w1095), .nZ(w1078) );
	vdp_not g1232 (.A(w1097), .nZ(w1077) );
	vdp_not g1233 (.A(w1096), .nZ(w1076) );
	vdp_aon222 g1234 (.C2(w1076), .B2(w1077), .A2(w1078), .C1(w1057), .B1(CA[15]), .A1(CA[7]), .Z(w1063) );
	vdp_aon222 g1235 (.C2(w1076), .B2(w1077), .A2(w1078), .C1(w1056), .B1(CA[13]), .A1(CA[6]), .Z(w1075) );
	vdp_aon222 g1236 (.C2(w1076), .B2(w1077), .A2(w1078), .C1(w1055), .B1(CA[12]), .A1(CA[5]), .Z(w1064) );
	vdp_aon222 g1237 (.C2(w1076), .B2(w1077), .A2(w1078), .C1(w1054), .B1(CA[11]), .A1(CA[4]), .Z(w1065) );
	vdp_aon222 g1238 (.C2(w1076), .B2(w1077), .A2(w1078), .C1(w1058), .B1(CA[10]), .A1(CA[3]), .Z(w1066) );
	vdp_aon222 g1239 (.C2(w1076), .B2(w1077), .A2(w1078), .C1(w1467), .B1(CA[9]), .A1(CA[2]), .Z(w1067) );
	vdp_aon222 g1240 (.C2(w1076), .B2(w1077), .A2(w1078), .C1(w1061), .B1(CA[8]), .A1(CA[1]), .Z(w1074) );
	vdp_aon222 g1241 (.C2(w1076), .B2(w1077), .A2(w1078), .C1(w1050), .B1(CA[14]), .A1(CA[0]), .Z(w1068) );
	vdp_aon222 g1242 (.C2(w1076), .B2(w1077), .A2(w1078), .C1(nHCLK1), .B1(1'b1), .A1(1'b0), .Z(w1079) );
	vdp_slatch g1243 (.Q(w1016), .D(LSM0), .C(w1046), .nC(w1047) );
	vdp_slatch g1244 (.Q(w1045), .D(LSM1), .C(w1046), .nC(w1047) );
	vdp_aon22 g1245 (.Z(w1049), .A1(COL[6]), .A2(w1086), .B1(w114), .B2(w1432) );
	vdp_not g1246 (.A(M2), .nZ(w1044) );
	vdp_not g1247 (.A(w1086), .nZ(w1432) );
	vdp_and g1248 (.Z(w1), .A(w1045), .B(w1016) );
	vdp_and g1249 (.Z(w1739), .A(M5), .B(w1044) );
	vdp_and g1250 (.Z(M2), .A(M5), .B(M2) );
	vdp_and g1251 (.Z(VRAM128k), .A(M5), .B(w1070) );
	vdp_or3 g1252 (.Z(w1090), .A(w1087), .B(w1088), .C(w1335) );
	vdp_and g1253 (.Z(w1089), .A(w1087), .B(w1059) );
	vdp_nand g1254 (.Z(w1097), .A(w1095), .B(w1090) );
	vdp_nand g1255 (.Z(w1096), .A(w1095), .B(w1093) );
	vdp_slatch g1256 (.Q(LSCR), .D(REG_BUS[0]), .C(w1072), .nC(w1073) );
	vdp_slatch g1257 (.Q(HSCR), .D(REG_BUS[1]), .C(w1072), .nC(w1073) );
	vdp_slatch g1258 (.Q(VSCR), .D(REG_BUS[2]), .C(w1072), .nC(w1073) );
	vdp_slatch g1259 (.Q(IE2), .D(REG_BUS[3]), .C(w1072), .nC(w1073) );
	vdp_slatch g1260 (.Q(w113), .D(REG_BUS[4]), .C(w1072), .nC(w1073) );
	vdp_slatch g1261 (.Q(w79), .D(REG_BUS[5]), .C(w1072), .nC(w1073) );
	vdp_slatch g1262 (.Q(w1028), .D(REG_BUS[6]), .C(w1072), .nC(w1073) );
	vdp_slatch g1263 (.Q(w1082), .D(REG_BUS[7]), .C(w1072), .nC(w1073) );
	vdp_slatch g1264 (.Q(M2), .D(REG_BUS[3]), .C(w1081), .nC(w1080) );
	vdp_slatch g1265 (.Q(w1070), .D(REG_BUS[7]), .C(w1081), .nC(w1080) );
	vdp_slatch g1266 (.Q(w18), .D(REG_BUS[4]), .C(w1084), .nC(w1085) );
	vdp_slatch g1267 (.Q(S_TE), .D(REG_BUS[3]), .C(w1084), .nC(w1085) );
	vdp_slatch g1268 (.Q(LSM1), .D(REG_BUS[2]), .C(w1084), .nC(w1085) );
	vdp_slatch g1269 (.Q(LSM0), .D(REG_BUS[1]), .C(w1084), .nC(w1085) );
	vdp_slatch g1270 (.Q(H40), .D(REG_BUS[0]), .C(w1084), .nC(w1085) );
	vdp_slatch g1271 (.Q(w42), .D(REG_BUS[0]), .C(w1081), .nC(w1080) );
	vdp_slatch g1272 (.Q(w117), .D(REG_BUS[1]), .C(w1081), .nC(w1080) );
	vdp_slatch g1273 (.Q(M5), .D(REG_BUS[2]), .C(w1081), .nC(w1080) );
	vdp_slatch g1274 (.Q(M1), .D(REG_BUS[4]), .C(w1081), .nC(w1080) );
	vdp_slatch g1275 (.Q(IE0), .D(REG_BUS[5]), .C(w1081), .nC(w1080) );
	vdp_slatch g1276 (.Q(DISP), .D(REG_BUS[6]), .C(w1081), .nC(w1080) );
	vdp_and g1277 (.Z(w106), .A(w1030), .B(w1109) );
	vdp_and g1278 (.Z(w105), .A(w980), .B(w1109) );
	vdp_and g1279 (.Z(w107), .A(w1030), .B(w1110) );
	vdp_and g1280 (.Z(w109), .A(w980), .B(w1110) );
	vdp_and g1281 (.Z(w102), .A(w1030), .B(w1104) );
	vdp_and g1282 (.Z(w112), .A(w980), .B(w1104) );
	vdp_and g1283 (.Z(w54), .A(w1030), .B(w1105) );
	vdp_and g1284 (.Z(w45), .A(w980), .B(w1105) );
	vdp_and g1285 (.Z(w75), .A(w1030), .B(w1107) );
	vdp_and g1286 (.Z(w73), .A(w980), .B(w1107) );
	vdp_and g1287 (.Z(w77), .A(w1030), .B(w1108) );
	vdp_and g1288 (.Z(PSG_TEST_OE), .A(w980), .B(w1108) );
	vdp_and g1289 (.Z(w1125), .A(w1030), .B(w1112) );
	vdp_and g1290 (.Z(w1101), .A(w1030), .B(w1113) );
	vdp_and g1291 (.Z(w53), .A(w1030), .B(w1106) );
	vdp_and g1292 (.Z(w51), .A(w980), .B(w1106) );
	vdp_dlatch g1293 (.D(COL[0]), .C(HCLK1), .Q(w1050), .nC(nHCLK1) );
	vdp_dlatch g1294 (.D(COL[1]), .Q(w1061), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch g1295 (.D(COL[2]), .Q(w1467), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch g1296 (.D(COL[3]), .Q(w1058), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch g1297 (.D(COL[4]), .Q(w1054), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch g1298 (.D(COL[5]), .Q(w1055), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch g1299 (.D(w1049), .Q(w1056), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch g1300 (.D(COL[7]), .Q(w1057), .C(HCLK1), .nC(nHCLK1) );
	vdp_slatch g1301 (.Q(w49), .D(REG_BUS[5]), .C(w1085), .nC(w1084) );
	vdp_slatch g1302 (.Q(w36), .D(REG_BUS[6]), .C(w1085), .nC(w1084) );
	vdp_slatch g1303 (.Q(RS0), .D(REG_BUS[7]), .C(w1085), .nC(w1084) );
	vdp_slatch g1304 (.Q(w22), .D(REG_BUS[3]), .nC(w1132), .C(w1130) );
	vdp_slatch g1305 (.Q(w82), .D(REG_BUS[2]), .nC(w1132), .C(w1130) );
	vdp_slatch g1306 (.Q(M3), .D(REG_BUS[1]), .nC(w1132), .C(w1130) );
	vdp_slatch g1307 (.Q(w50), .D(REG_BUS[0]), .nC(w1132), .C(w1130) );
	vdp_slatch g1308 (.Q(w80), .D(REG_BUS[7]), .nC(w1132), .C(w1130) );
	vdp_slatch g1309 (.Q(w81), .D(REG_BUS[6]), .nC(w1132), .C(w1130) );
	vdp_slatch g1310 (.Q(w56), .D(REG_BUS[5]), .nC(w1132), .C(w1130) );
	vdp_slatch g1311 (.Q(IE1), .D(REG_BUS[4]), .nC(w1132), .C(w1130) );
	vdp_slatch_r g1312 (.Q(w104), .D(DB[14]), .nC(w1124), .R(w1119), .C(w1128) );
	vdp_slatch_r g1313 (.Q(w111), .D(DB[13]), .R(w1119), .nC(w1124), .C(w1128) );
	vdp_slatch_r g1314 (.Q(w108), .D(DB[12]), .R(w1119), .nC(w1124), .C(w1128) );
	vdp_comp_str g1315 (.Z(w1130), .A(w1129), .nZ(w1132) );
	vdp_comp_str g1316 (.Z(w1127), .A(w1101), .nZ(w1126) );
	vdp_not g1317 (.A(REG_BUS[6]), .nZ(w1430) );
	vdp_not g1318 (.A(REG_BUS[7]), .nZ(w1145) );
	vdp_not g1319 (.A(REG_BUS[4]), .nZ(w1133) );
	vdp_not g1320 (.A(REG_BUS[5]), .nZ(w1131) );
	vdp_not g1321 (.A(REG_BUS[2]), .nZ(w1146) );
	vdp_not g1322 (.A(REG_BUS[3]), .nZ(w1134) );
	vdp_not g1323 (.A(REG_BUS[0]), .nZ(w1140) );
	vdp_not g1324 (.A(REG_BUS[1]), .nZ(w1141) );
	vdp_not g1325 (.A(w1117), .nZ(w1136) );
	vdp_not g1326 (.A(w1118), .nZ(w1122) );
	vdp_not g1327 (.A(w1111), .nZ(w1135) );
	vdp_not g1328 (.A(w1123), .nZ(w1137) );
	vdp_comp_str g1329 (.Z(w1121), .nZ(w1120), .A(w1031) );
	vdp_slatch_r g1330 (.Q(w1123), .R(w1119), .D(DB[11]), .nC(w1120), .C(w1121) );
	vdp_slatch_r g1331 (.Q(w1111), .D(DB[10]), .nC(w1120), .R(w1119), .C(w1121) );
	vdp_and4 g1332 (.Z(w1441), .A(w1117), .B(w1118), .C(w1123), .D(w1111) );
	vdp_and4 g1333 (.Z(w1104), .A(w1123), .B(w1135), .C(w1122), .D(w1136) );
	vdp_and4 g1334 (.Z(w1110), .A(w1137), .B(w1111), .C(w1118), .D(w1117) );
	vdp_and4 g1335 (.Z(w1109), .A(w1137), .B(w1111), .C(w1118), .D(w1136) );
	vdp_and4 g1336 (.Z(w1108), .A(w1137), .B(w1111), .C(w1122), .D(w1117) );
	vdp_and4 g1337 (.Z(w1107), .A(w1137), .B(w1111), .C(w1122), .D(w1136) );
	vdp_and4 g1338 (.Z(w1105), .A(w1137), .B(w1135), .C(w1118), .D(w1117) );
	vdp_and4 g1339 (.Z(w1106), .A(w1137), .B(w1135), .C(w1118), .D(w1136) );
	vdp_and4 g1340 (.Z(w1113), .A(w1137), .B(w1135), .C(w1122), .D(w1117) );
	vdp_and4 g1341 (.Z(w1112), .A(w1137), .B(w1135), .C(w1122), .D(w1136) );
	vdp_nand g1342 (.Z(w1374), .A(w1441), .B(w1030) );
	vdp_slatch_r g1343 (.Q(w1117), .D(DB[8]), .R(w1119), .C(w1121), .nC(w1120) );
	vdp_slatch_r g1344 (.Q(PSG_TEST11), .D(DB[11]), .R(w1119), .C(w1128), .nC(w1124) );
	vdp_slatch_r g1345 (.nC(w1120), .Q(w1118), .D(DB[9]), .R(w1119), .C(w1121) );
	vdp_slatch_r g1346 (.Q(PSG_TEST10), .D(DB[10]), .R(w1119), .C(w1128), .nC(w1124) );
	vdp_slatch_r g1347 (.Q(w84), .D(DB[8]), .R(w1119), .C(w1128), .nC(w1124) );
	vdp_slatch_r g1348 (.Q(PSG_TEST9), .D(DB[9]), .R(w1119), .C(w1128), .nC(w1124) );
	vdp_slatch_r g1349 (.Q(w83), .D(DB[7]), .R(w1119), .C(w1128), .nC(w1124) );
	vdp_slatch_r g1350 (.Q(w85), .D(DB[5]), .R(w1119), .C(w1128), .nC(w1124) );
	vdp_slatch_r g1351 (.Q(w86), .D(DB[6]), .R(w1119), .C(w1128), .nC(w1124) );
	vdp_slatch_r g1352 (.Q(w942), .D(DB[4]), .R(w1119), .C(w1128), .nC(w1124) );
	vdp_slatch_r g1353 (.Q(w1143), .D(DB[2]), .R(w1119), .C(w1128), .nC(w1124) );
	vdp_slatch_r g1354 (.Q(w1144), .D(DB[3]), .R(w1119), .C(w1128), .nC(w1124) );
	vdp_slatch_r g1355 (.Q(w1086), .D(DB[0]), .R(w1119), .C(w1128), .nC(w1124) );
	vdp_slatch_r g1356 (.Q(w749), .D(DB[1]), .R(w1119), .C(w1128), .nC(w1124) );
	vdp_slatch_r g1357 (.Q(w90), .D(DB[9]), .R(w1119), .C(w1127), .nC(w1126) );
	vdp_slatch_r g1358 (.Q(w91), .D(DB[10]), .R(w1119), .C(w1127), .nC(w1126) );
	vdp_slatch_r g1359 (.Q(w88), .D(DB[7]), .R(w1119), .C(w1127), .nC(w1126) );
	vdp_slatch_r g1360 (.Q(w89), .D(DB[8]), .R(w1119), .C(w1127), .nC(w1126) );
	vdp_slatch_r g1361 (.Q(w48), .D(DB[5]), .R(w1119), .C(w1127), .nC(w1126) );
	vdp_slatch_r g1362 (.Q(w38), .D(DB[6]), .R(w1119), .C(w1127), .nC(w1126) );
	vdp_slatch_r g1363 (.Q(w37), .D(DB[3]), .R(w1119), .C(w1127), .nC(w1126) );
	vdp_slatch_r g1364 (.Q(w39), .D(DB[4]), .R(w1119), .C(w1127), .nC(w1126) );
	vdp_slatch_r g1365 (.Q(w1431), .D(DB[1]), .R(w1119), .C(w1127), .nC(w1126) );
	vdp_slatch_r g1366 (.Q(w52), .D(DB[2]), .R(w1119), .C(w1127), .nC(w1126) );
	vdp_slatch_r g1367 (.Q(w40), .D(DB[0]), .R(w1119), .C(w1127), .nC(w1126) );
	vdp_comp_str g1368 (.Z(w1128), .nZ(w1124), .A(w1125) );
	vdp_notif0 g1369 (.A(VPOS[9]), .nZ(DB[10]), .nE(w1138) );
	vdp_notif0 g1370 (.A(VPOS[8]), .nZ(DB[9]), .nE(w1138) );
	vdp_bufif0 g1371 (.A(FIFO_EMPTY), .Z(DB[9]), .nE(w1168) );
	vdp_bufif0 g1372 (.A(FIFO_FULL), .Z(DB[8]), .nE(w1168) );
	vdp_bufif0 g1373 (.A(w1167), .Z(DB[1]), .nE(w1168) );
	vdp_bufif0 g1374 (.A(w1169), .Z(DB[0]), .nE(w1168) );
	vdp_bufif0 g1375 (.A(w1150), .Z(DB[7]), .nE(w1168) );
	vdp_bufif0 g1376 (.A(w1149), .Z(DB[6]), .nE(w1168) );
	vdp_bufif0 g1377 (.A(w1148), .Z(DB[5]), .nE(w1168) );
	vdp_bufif0 g1378 (.A(ODD_EVEN), .Z(DB[4]), .nE(w1168) );
	vdp_bufif0 g1379 (.A(w43), .Z(DB[3]), .nE(w1168) );
	vdp_bufif0 g1380 (.A(w20), .Z(DB[2]), .nE(w1168) );
	vdp_slatch_r g1381 (.Q(w69), .D(DB[4]), .R(w1119), .C(w1121), .nC(w1120) );
	vdp_slatch_r g1382 (.Q(w70), .D(DB[5]), .R(w1119), .C(w1121), .nC(w1120) );
	vdp_slatch_r g1383 (.Q(w72), .D(DB[7]), .R(w1119), .C(w1121), .nC(w1120) );
	vdp_slatch_r g1384 (.Q(w71), .D(DB[6]), .R(w1119), .C(w1121), .nC(w1120) );
	vdp_slatch_r g1385 (.Q(w65), .D(DB[0]), .R(w1119), .C(w1121), .nC(w1120) );
	vdp_slatch_r g1386 (.Q(w66), .D(DB[1]), .R(w1119), .C(w1121), .nC(w1120) );
	vdp_slatch_r g1387 (.Q(w68), .D(DB[3]), .R(w1119), .C(w1121), .nC(w1120) );
	vdp_slatch_r g1388 (.Q(w67), .D(DB[2]), .R(w1119), .C(w1121), .nC(w1120) );
	vdp_notif0 g1389 (.A(HPOS[0]), .nZ(DB[8]), .nE(w1138) );
	vdp_not g1390 (.A(nSEL0_M3), .nZ(w1442) );
	vdp_comp_str g1391 (.Z(w1139), .A(w771), .nZ(w1142) );
	vdp_slatch_r g1392 (.Q(HIT[0]), .D(w1140), .R(SYSRES), .C(w1139), .nC(w1142) );
	vdp_slatch_r g1393 (.Q(HIT[2]), .D(w1146), .R(SYSRES), .C(w1139), .nC(w1142) );
	vdp_slatch_r g1394 (.Q(HIT[1]), .D(w1141), .R(SYSRES), .C(w1139), .nC(w1142) );
	vdp_slatch_r g1395 (.Q(HIT[6]), .D(w1430), .R(SYSRES), .C(w1139), .nC(w1142) );
	vdp_slatch_r g1396 (.Q(HIT[3]), .D(w1134), .R(SYSRES), .C(w1139), .nC(w1142) );
	vdp_slatch_r g1397 (.Q(HIT[5]), .D(w1131), .R(SYSRES), .C(w1139), .nC(w1142) );
	vdp_slatch_r g1398 (.Q(HIT[4]), .D(w1133), .R(SYSRES), .C(w1139), .nC(w1142) );
	vdp_slatch_r g1399 (.Q(HIT[7]), .D(w1145), .R(SYSRES), .C(w1139), .nC(w1142) );
	vdp_aon22 g1400 (.Z(w1167), .A1(FIFO_EMPTY), .A2(w1152), .B1(w1153), .B2(DMA_BUSY) );
	vdp_aon22 g1401 (.Z(w1169), .A1(FIFO_FULL), .A2(w1152), .B1(w1153), .B2(PAL) );
	vdp_and3 g1402 (.C(w1143), .A(w377), .B(w1442), .Z(w1147) );
	vdp_not g1403 (.A(w1147), .nZ(w1138) );
	vdp_not g1404 (.A(w960), .nZ(w1168) );
	vdp_cnt_bit_load g1405 (.D(HIT[7]), .nL(w1174), .L(w1155), .R(1'b0), .Q(w1175), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1201) );
	vdp_cnt_bit_load g1406 (.D(HIT[6]), .nL(w1174), .L(w1155), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1477), .CO(w1201) );
	vdp_cnt_bit_load g1407 (.D(HIT[5]), .nL(w1174), .L(w1155), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1200), .CO(w1477) );
	vdp_cnt_bit_load g1408 (.D(HIT[4]), .nL(w1174), .L(w1155), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1199), .CO(w1200) );
	vdp_cnt_bit_load g1409 (.D(HIT[3]), .nL(w1174), .L(w1155), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1198), .CO(w1199) );
	vdp_cnt_bit_load g1410 (.D(HIT[2]), .nL(w1174), .L(w1155), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1487), .CO(w1198) );
	vdp_cnt_bit_load g1411 (.D(HIT[1]), .nL(w1174), .L(w1155), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1197), .CO(w1487) );
	vdp_cnt_bit_load g1412 (.D(HIT[0]), .nL(w1174), .L(w1155), .R(1'b0), .CI(w1172), .CO(w1197), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g1413 (.D(w1438), .C2(HCLK2), .C1(HCLK1), .Q(w1176), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_rs_ff g1414 (.Q(w1149), .R(w1191), .S(w1192) );
	vdp_rs_ff g1415 (.Q(w1150), .R(w1190), .S(V_INT_HAPPENED) );
	vdp_rs_ff g1416 (.Q(w1148), .R(w1191), .S(COLLISION) );
	vdp_not g1417 (.A(M5), .nZ(w1189) );
	vdp_not g1418 (.A(w1150), .nZ(w1171) );
	vdp_not g1419 (.A(w1156), .nZ(w1161) );
	vdp_not g1420 (.A(CA[21]), .nZ(w1439) );
	vdp_not g1421 (.A(nSEL0_M3), .nZ(w1162) );
	vdp_not g1422 (.A(w1194), .nZ(w1163) );
	vdp_comp_we g1423 (.Z(w1174), .A(w1437), .nZ(w1155) );
	vdp_or g1424 (.A(w1194), .B(w1176), .Z(w1437) );
	vdp_and g1425 (.A(w1163), .B(w1175), .Z(w1438) );
	vdp_and g1426 (.A(w1171), .B(SPRITE_OVF), .Z(w1192) );
	vdp_or g1427 (.A(w1144), .B(w4), .Z(w1172) );
	vdp_not g1428 (.A(w1152), .nZ(w1153) );
	vdp_nor3 g1429 (.A(nSEL0_M3), .B(w1189), .Z(w1152), .C(CA[1]) );
	vdp_nor3 g1430 (.A(w1144), .B(w5), .Z(w1194), .C(w29) );
	vdp_nor g1431 (.A(w1196), .B(w1177), .Z(w1160) );
	vdp_or5 g1432 (.A(w1162), .B(CA[4]), .C(CA[5]), .D(CA[15]), .Z(w1196), .E(CA[6]) );
	vdp_or5 g1433 (.A(CA[16]), .B(CA[17]), .C(CA[20]), .D(w1161), .Z(w1177), .E(w1439) );
	vdp_rs_ff g1434 (.Q(w1182), .R(w1233), .S(w1438) );
	vdp_rs_ff g1435 (.Q(w1234), .R(w1217), .S(w1440) );
	vdp_dff g1436 (.Q(w1236), .R(w1195), .C(w1185), .D(w1178) );
	vdp_dff g1437 (.Q(w1235), .R(w1195), .C(w1185), .D(w1292) );
	vdp_dff g1438 (.Q(w1237), .R(w1195), .C(w1185), .D(w1179) );
	vdp_rs_ff g1439 (.Q(w1493), .R(w1232), .S(w1492) );
	vdp_rs_ff g1440 (.Q(w1205), .R(w1206), .S(w1490) );
	vdp_dlatch_inv g1441 (.D(w1212), .Q(w1213), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g1442 (.D(w1206), .C(DCLK1), .Q(w1212), .nC(nDCLK1) );
	vdp_dlatch_inv g1443 (.D(w1215), .Q(w1191), .C(HCLK1), .nC(nHCLK1) );
	vdp_not g1444 (.A(w1228), .nZ(w1202) );
	vdp_not g1445 (.A(w631), .nZ(w1181) );
	vdp_not g1446 (.A(w1184), .nZ(w1179) );
	vdp_not g1447 (.A(w1183), .nZ(w1178) );
	vdp_not g1448 (.A(w1193), .nZ(w1195) );
	vdp_not g1449 (.A(w1209), .nZ(w1185) );
	vdp_not g1450 (.A(w1186), .nZ(w47) );
	vdp_not g1451 (.A(w1187), .nZ(w1188) );
	vdp_sr_bit g1452 (.D(w1214), .C2(HCLK2), .C1(HCLK1), .Q(w1232), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and g1453 (.A(M5), .B(w1205), .Z(w1209) );
	vdp_and g1454 (.A(nSEL0_M3), .B(w1204), .Z(w1037) );
	vdp_and g1455 (.A(w1186), .B(w1037), .Z(w1491) );
	vdp_or g1456 (.A(w978), .B(w1491), .Z(w1490) );
	vdp_or g1457 (.A(w960), .B(SYSRES), .Z(w1492) );
	vdp_and g1458 (.A(w1189), .B(w1191), .Z(w1216) );
	vdp_or g1459 (.A(w1235), .B(w1216), .Z(w1217) );
	vdp_and g1460 (.A(M5), .B(w438), .Z(w1440) );
	vdp_and g1461 (.A(M1), .B(M5), .Z(w1180) );
	vdp_or g1462 (.A(w1237), .B(w1216), .Z(w1190) );
	vdp_or g1463 (.A(w1236), .B(w1216), .Z(w1233) );
	vdp_comp_dff g1464 (.D(w1493), .C2(HCLK2), .C1(HCLK1), .Q(w1214), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_comp_dff g1465 (.D(w1209), .C2(DCLK2), .C1(DCLK1), .Q(w1206), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_nor g1466 (.A(w1214), .B(SYSRES), .Z(w1515) );
	vdp_nand g1467 (.A(w1232), .B(w1515), .Z(w1215) );
	vdp_nand g1468 (.A(w1150), .B(IE0), .Z(w1184) );
	vdp_and3 g1469 (.A(w1180), .B(w889), .Z(w1227), .C(w1181) );
	vdp_and3 g1470 (.A(w1180), .B(w889), .Z(w1226), .C(w631) );
	vdp_and4 g1471 (.A(w1183), .B(IE2), .C(w1184), .D(w1234), .Z(w1292) );
	vdp_nand3 g1472 (.C(w1182), .A(w1184), .B(IE1), .Z(w1183) );
	vdp_aoi21 g1473 (.A1(w1213), .B(SYSRES), .Z(w1193), .A2(w1212) );
	vdp_dff g1474 (.Q(w1256), .R(w1242), .C(w1239), .D(w1225) );
	vdp_dff g1475 (.Q(w1252), .R(w1242), .C(w1239), .D(w1251) );
	vdp_dff g1476 (.Q(w1222), .R(w1242), .C(w1239), .D(w1220) );
	vdp_dff g1477 (.Q(w1230), .R(w1242), .C(w1239), .D(w1229) );
	vdp_dff g1478 (.Q(w1231), .R(w1242), .C(w1239), .D(w1219) );
	vdp_dff g1479 (.Q(w1210), .R(w1242), .C(w1239), .D(w1247) );
	vdp_dff g1480 (.Q(w1207), .R(w1242), .C(w1239), .D(w1245) );
	vdp_dff g1481 (.Q(w1238), .R(1'b0), .C(w1239), .D(w1203) );
	vdp_ha g1482 (.SUM(w1245), .A(w1207), .B(w1202), .CO(w1208) );
	vdp_ha g1483 (.SUM(w1247), .A(w1210), .B(w1208), .CO(w1211) );
	vdp_ha g1484 (.SUM(w1219), .A(w1231), .B(w1211), .CO(w1218) );
	vdp_ha g1485 (.SUM(w1229), .A(w1230), .B(w1218), .CO(w1223) );
	vdp_ha g1486 (.SUM(w1220), .A(w1222), .B(w1223), .CO(w1221) );
	vdp_ha g1487 (.SUM(w1225), .A(w1256), .B(w1221), .CO(w1224) );
	vdp_ha g1488 (.SUM(w1251), .A(w1252), .B(w1224) );
	vdp_and3 g1489 (.A(w1252), .B(w1222), .Z(w1249), .C(w1256) );
	vdp_and4 g1490 (.C(w1210), .A(w1230), .B(w1249), .Z(w1255), .D(w1231) );
	vdp_nand g1491 (.A(w1238), .B(nSEL0_M3), .Z(w1372) );
	vdp_dff g1492 (.Q(w1263), .R(1'b0), .C(w1239), .D(w1244) );
	vdp_dff g1493 (.Q(w1244), .R(w1246), .C(w1239), .D(w1268) );
	vdp_dff g1494 (.Q(w1268), .R(w1246), .C(w1266), .D(w1248) );
	vdp_dff g1495 (.Q(w1248), .R(w1246), .C(w1239), .D(w1272) );
	vdp_dff g1496 (.Q(w1272), .R(w1246), .C(w1239), .D(w1273) );
	vdp_dff g1497 (.Q(w1273), .R(w1246), .C(w1239), .D(1'b1) );
	vdp_dff g1498 (.Q(w1480), .R(w1281), .C(w1257), .D(w1249) );
	vdp_dff g1499 (.Q(w1257), .R(1'b0), .C(w1239), .D(w1255) );
	vdp_dff g1500 (.Q(w1274), .R(w1254), .C(w1275), .D(w1249) );
	vdp_dff g1501 (.Q(w1253), .R(w1267), .C(w1279), .D(1'b1) );
	vdp_or g1502 (.A(SYSRES), .B(w1253), .Z(w1254) );
	vdp_or g1503 (.A(w1246), .B(w1263), .Z(w1277) );
	vdp_not g1504 (.A(w1263), .nZ(w1241) );
	vdp_not g1505 (.A(w1480), .nZ(w1246) );
	vdp_nand3 g1506 (.A(nSEL0_M3), .B(w1261), .Z(w1242), .C(w1241) );
	vdp_not g1507 (.nZ(w1266), .A(w1262) );
	vdp_not g1508 (.nZ(w1239), .A(w1240) );
	vdp_dff g1509 (.Q(w1265), .R(1'b0), .C(w1266), .D(w1284) );
	vdp_dff g1510 (.Q(w1288), .R(w1267), .C(w1266), .D(w1271) );
	vdp_dff g1511 (.Q(w1271), .R(w1267), .C(w1239), .D(w1290) );
	vdp_dff g1512 (.Q(w1290), .R(w1267), .C(w1266), .D(w1270) );
	vdp_dff g1513 (.Q(w1270), .R(w1267), .C(w1266), .D(w1280) );
	vdp_dff g1514 (.Q(w1280), .R(w1267), .C(w1239), .D(w44) );
	vdp_dff g1515 (.Q(w1296), .R(w1295), .C(w1266), .D(w1088) );
	vdp_dff g1516 (.Q(w1088), .R(w1295), .C(w1239), .D(w1276) );
	vdp_not g1517 (.A(w1282), .nZ(w97) );
	vdp_not g1518 (.A(w958), .nZ(w1260) );
	vdp_not g1519 (.A(w1271), .nZ(w1269) );
	vdp_not g1520 (.A(w1268), .nZ(w1488) );
	vdp_not g1521 (.A(w1276), .nZ(w1295) );
	vdp_not g1522 (.A(w1037), .nZ(w1279) );
	vdp_not g1523 (.A(w1186), .nZ(w1481) );
	vdp_and g1524 (.A(w1277), .B(w1037), .Z(w1276) );
	vdp_and g1525 (.A(w1278), .B(w1276), .Z(w1275) );
	vdp_and g1526 (.A(w1296), .B(w1275), .Z(w44) );
	vdp_and g1527 (.A(w1272), .B(w1488), .Z(w1285) );
	vdp_and g1528 (.A(w1273), .B(w1488), .Z(w1287) );
	vdp_and g1529 (.A(w1264), .B(w949), .Z(w1286) );
	vdp_and g1530 (.A(w1264), .B(w992), .Z(w1259) );
	vdp_and g1531 (.A(w958), .B(w1265), .Z(w1264) );
	vdp_and g1532 (.A(w97), .B(w1088), .Z(w1024) );
	vdp_nand g1533 (.A(w1270), .B(w1269), .Z(w1261) );
	vdp_nor g1534 (.A(w1267), .B(w1280), .Z(w1289) );
	vdp_or3 g1535 (.C(w1274), .A(SYSRES), .B(w1263), .Z(w1281) );
	vdp_oai21 g1536 (.A1(w992), .B(w1260), .Z(w1282), .A2(w949) );
	vdp_dff g1537 (.Q(w1351), .R(1'b0), .C(w1239), .D(w1187) );
	vdp_rs_ff g1538 (.nQ(w1034), .R(w1303), .S(w1301) );
	vdp_not g1539 (.A(w1308), .nZ(PSG_Z80_CLK) );
	vdp_not g1540 (.A(REG_BUS[7]), .nZ(w1300) );
	vdp_and3 g1541 (.C(w1300), .A(w787), .B(M5), .Z(w1301) );
	vdp_or g1542 (.A(w1187), .B(SYSRES), .Z(w1303) );
	vdp_and g1543 (.A(w1319), .B(w757), .Z(w1320) );
	vdp_not g1544 (.A(w1278), .nZ(w1322) );
	vdp_and4 g1545 (.C(CA[21]), .A(w1156), .B(CA[20]), .Z(w1278), .D(w1481) );
	vdp_dff g1546 (.Q(w1360), .R(1'b0), .C(w1308), .D(w1344) );
	vdp_dff g1547 (.Q(w1339), .R(1'b0), .C(w1308), .D(w1338) );
	vdp_dff g1548 (.Q(w1283), .R(1'b0), .C(w1325), .D(w1326) );
	vdp_dff g1549 (.Q(w1338), .R(1'b0), .C(w1325), .D(w1283) );
	vdp_dff g1550 (.Q(w1352), .R(w1353), .C(HCLK2), .D(w1355) );
	vdp_dff g1551 (.Q(DMA_BUSY), .R(w1353), .C(HCLK2), .D(w1352) );
	vdp_rs_ff g1552 (.Q(w1228), .R(w1353), .S(w1293) );
	vdp_rs_ff g1553 (.Q(w1482), .R(w1353), .S(w1226) );
	vdp_rs_ff g1554 (.Q(w1203), .R(w1294), .S(w1227) );
	vdp_sr_bit g1555 (.D(w757), .Q(w1319), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1556 (.D(w1489), .Q(w1350), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_dlatch_inv g1557 (.D(w1318), .nQ(w1299), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g1558 (.D(w1349), .nQ(w1318), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g1559 (.D(w1305), .C(HCLK1), .nQ(w1349), .nC(nHCLK1) );
	vdp_aon22 g1560 (.Z(w1346), .A2(w1298), .B1(w1349), .B2(w1356), .A1(w1299) );
	vdp_sr_bit g1561 (.D(w1357), .Q(w1362), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1562 (.D(w1321), .Q(w1357), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1563 (.D(VRAM_REFRESH), .C2(HCLK2), .C1(HCLK1), .Q(w1321), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_aon22 g1564 (.Z(w1334), .A2(w1289), .B1(w1363), .B2(w1364), .A1(w1332) );
	vdp_not g1565 (.A(w1479), .nZ(w1027) );
	vdp_not g1566 (.A(w1289), .nZ(w1364) );
	vdp_not g1567 (.A(w1350), .nZ(w1356) );
	vdp_not g1568 (.A(w1297), .nZ(w1333) );
	vdp_not g1569 (.A(w1274), .nZ(w1267) );
	vdp_or g1570 (.A(w1228), .B(w1482), .Z(w1355) );
	vdp_or g1571 (.A(SYSRES), .B(w1007), .Z(w1353) );
	vdp_or g1572 (.A(w1293), .B(w1353), .Z(w1294) );
	vdp_or g1573 (.A(w1179), .B(w1292), .Z(w258) );
	vdp_or g1574 (.A(w1179), .B(w1178), .Z(w234) );
	vdp_and g1575 (.A(w1350), .B(w607), .Z(w1298) );
	vdp_or g1576 (.A(w1299), .B(w1357) );
	vdp_and g1577 (.A(w1261), .B(w1275), .Z(w1332) );
	vdp_and g1578 (.A(w1290), .B(w1275), .Z(w1363) );
	vdp_and g1579 (.A(w1275), .B(w1267), .Z(w99) );
	vdp_and g1580 (.A(w953), .B(w100), .Z(w1345) );
	vdp_or g1581 (.A(w1286), .B(w957), .Z(w1341) );
	vdp_aon22 g1582 (.Z(w1370), .A2(w1028), .B1(w1291), .B2(w1337), .A1(w1336) );
	vdp_and g1583 (.A(w1344), .B(w1360), .Z(w1087) );
	vdp_and g1584 (.A(w1358), .B(w1365), .Z(w1347) );
	vdp_and g1585 (.A(w1365), .B(w1361), .Z(w1344) );
	vdp_not g1586 (.A(w1361), .nZ(w1358) );
	vdp_not g1587 (.A(w1359), .nZ(w1365) );
	vdp_not g1588 (.A(w1318), .nZ(w1354) );
	vdp_not g1589 (.A(w1330), .nZ(w1348) );
	vdp_and g1590 (.A(w1342), .B(w1310), .Z(w1309) );
	vdp_and g1591 (.A(w1342), .B(w1312), .Z(w952) );
	vdp_and g1592 (.A(w1342), .B(w1314), .Z(w957) );
	vdp_and g1593 (.A(w1342), .B(w1311), .Z(w953) );
	vdp_and g1594 (.A(w1342), .B(w1313), .Z(w1326) );
	vdp_and g1595 (.A(w952), .B(w1326), .Z(w978) );
	vdp_and g1596 (.A(nSEL0_M3), .B(w1323), .Z(w949) );
	vdp_and g1597 (.A(nSEL0_M3), .B(w1315), .Z(w992) );
	vdp_not g1598 (.A(nSEL0_M3), .nZ(w1342) );
	vdp_nand g1599 (.A(w1338), .B(w1339), .Z(w1361) );
	vdp_nand g1600 (.A(FIFO_FULL), .B(w1307), .Z(w1306) );
	vdp_nand g1601 (.A(nSEL0_M3), .B(w234), .Z(w1317) );
	vdp_nand g1602 (.A(w258), .B(nSEL0_M3), .Z(w1316) );
	vdp_or3 g1603 (.C(w1179), .A(w1178), .B(w1292), .Z(w1020) );
	vdp_and3 g1604 (.C(w1299), .A(w757), .B(w1350), .Z(w558) );
	vdp_aoi21 g1605 (.A2(w1298), .B(w1354), .Z(w1297), .A1(w1349) );
	vdp_nor g1606 (.A(w1321), .B(w1362), .Z(w1307) );
	vdp_nand g1607 (.A(w97), .B(w1322), .Z(w1330) );
	vdp_nand3 g1608 (.C(w1306), .A(w3), .B(w1320), .Z(w1305) );
	vdp_2a3oi g1609 (.A1(w1354), .B(w632), .Z(w1304), .A2(w1349), .C(w1350) );
	vdp_nor4 g1610 (.C(VRAM_REFRESH), .A(w1357), .B(w1321), .Z(w1489), .D(w1362) );
	vdp_comb1 g1611 (.A(w1309), .B(w1358), .Z(w1359), .C2(CA[14]), .C1(CA[15]) );
	vdp_aon22 g1612 (.Z(w1371), .A2(w1028), .B1(w1291), .B2(w1331), .A1(w1478) );
	vdp_not g1613 (.A(w1028), .nZ(w1291) );
	vdp_or4 g1614 (.C(w1333), .A(w1365), .B(w1332), .Z(w1478), .D(w1285) );
	vdp_or4 g1615 (.C(w1299), .A(w1348), .B(w1345), .Z(w1337), .D(w1299) );
	vdp_or3 g1616 (.C(w1334), .A(w1344), .B(w1335), .Z(w1331) );
	vdp_comb1 g1617 (.C1(w1088), .B(w1271), .Z(w1479), .C2(w1289), .A(w1275) );
	vdp_and6 g1618 (.C(w1328), .A(w1238), .B(w1327), .Z(w1293), .D(w1351), .E(nSEL0_M3), .F(w1279) );
	vdp_or5 g1619 (.C(w1346), .A(w1338), .B(w44), .Z(w1336), .D(w1287), .E(w1089) );
	vdp_or5 g1620 (.C(w1299), .A(w1347), .B(w98), .Z(w1340), .D(w1285), .E(w1345) );
	vdp_aoi22 g1621 (.Z(w1284), .A2(w44), .B1(w1288), .B2(w1275), .A1(w1289) );
	vdp_n_fet g1622 (.Z(w284), .A(w393) );
	vdp_n_fet g1623 (.Z(w1466), .A(w393) );
	vdp_n_fet g1624 (.A(w393), .Z(w276) );
	vdp_n_fet g1625 (.A(w393), .Z(w242) );
	vdp_n_fet g1626 (.Z(w1465), .A(w393) );
	vdp_n_fet g1627 (.Z(w235), .A(w393) );
	vdp_n_fet g1628 (.Z(w1396), .A(w393) );
	vdp_n_fet g1629 (.Z(w1549), .A(w393) );
	vdp_aon22 g1630 (.Z(w1335), .A2(w1298), .B1(w1298), .B2(w1354), .A1(w1299) );
	vdp_comp_we g1631 (.nZ(w1308), .Z(w1325), .A(w1343) );
	vdp_comp_we g1632 (.nZ(w1240), .Z(w1262), .A(w1373) );
	vdp_not g1633 (.nZ(w1572), .A(w1904) );
	vdp_not g1634 (.nZ(w1574), .A(w1575) );
	vdp_sr_bit g1635 (.Q(w5), .D(w1899), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1636 (.Q(w1580), .D(VPLA7), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1637 (.Q(w1555), .D(VPLA6), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1638 (.Q(w1603), .D(w1577), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1639 (.Q(w1557), .D(VPLA5), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1640 (.Q(w1561), .D(VPLA4), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1641 (.Q(w1740), .D(VPLA0), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1642 (.Q(w1588), .D(w1586), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1643 (.Q(w1585), .D(VPLA2), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1644 (.Q(w1562), .D(VPLA3), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1645 (.Q(w1595), .D(w1779), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1646 (.Q(w1593), .D(w1590), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1647 (.Q(w1590), .D(w1916), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1648 (.Q(w1594), .D(w1597), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1649 (.Q(w1567), .D(w1863), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_not g1650 (.nZ(w1586), .A(VPLA1) );
	vdp_not g1651 (.nZ(w55), .A(w1585) );
	vdp_not g1652 (.nZ(w1571), .A(w1585) );
	vdp_not g1653 (.nZ(w1564), .A(ODD_EVEN) );
	vdp_not g1654 (.nZ(w1573), .A(w1016) );
	vdp_not g1655 (.nZ(w1916), .A(w1900) );
	vdp_not g1656 (.nZ(w1599), .A(w1600) );
	vdp_not g1657 (.nZ(w1587), .A(w1901) );
	vdp_not g1658 (.nZ(w1592), .A(w1593) );
	vdp_not g1659 (.nZ(w1569), .A(w50) );
	vdp_and g1660 (.Z(w1591), .A(w1774), .B(w1595) );
	vdp_nor g1661 (.Z(w1589), .A(SYSRES), .B(w1561) );
	vdp_oai21 g1662 (.Z(w1900), .B(w1589), .A2(w1599), .A1(w1590) );
	vdp_oai21 g1663 (.Z(w1600), .B(w1598), .A2(w1597), .A1(w1779) );
	vdp_aoi21 g1664 (.Z(w1901), .B(SYSRES), .A2(w1594), .A1(w1774) );
	vdp_and g1665 (.Z(w1568), .A(w1571), .B(w34) );
	vdp_and3 g1666 (.Z(w1774), .A(w1592), .B(w50), .C(w1590) );
	vdp_or g1667 (.Z(w1570), .A(SYSRES), .B(w1571) );
	vdp_and g1668 (.Z(w1863), .A(w1565), .B(w1575) );
	vdp_and g1669 (.Z(w1576), .A(w1568), .B(w1569) );
	vdp_and g1670 (.Z(w1565), .A(w1568), .B(w50) );
	vdp_and g1671 (.Z(w1560), .A(w1556), .B(w1562) );
	vdp_or g1672 (.Z(w1559), .A(SYSRES), .B(w1560) );
	vdp_2a3oi g1673 (.Z(w1904), .A1(w1574), .A2(w1565), .C(SYSRES), .B(w1573) );
	vdp_or g1674 (.Z(w1556), .A(w1563), .B(w1564) );
	vdp_or g1675 (.Z(w1558), .A(SYSRES), .B(w1601) );
	vdp_and g1676 (.Z(w1601), .A(w1556), .B(w1557) );
	vdp_and g1677 (.Z(w1581), .A(w1556), .B(w1580) );
	vdp_and g1678 (.Z(w1579), .A(w1556), .B(w1555) );
	vdp_or g1679 (.Z(w1850), .A(SYSRES), .B(w1601) );
	vdp_and g1680 (.Z(w1781), .A(w1577), .B(M5) );
	vdp_not g1681 (.nZ(w43), .A(w1583) );
	vdp_not g1682 (.nZ(w1583), .A(w1582) );
	vdp_not g1683 (.nZ(w1776), .A(w1582) );
	vdp_not g1684 (.nZ(w1899), .A(w1750) );
	vdp_and g1685 (.Z(w1669), .A(M5), .B(w1578) );
	vdp_or g1686 (.Z(w1584), .A(SYSRES), .B(w1581) );
	vdp_oai21 g1687 (.Z(w1582), .B(DISP), .A2(w29), .A1(w5) );
	vdp_rs_ff g1688 (.Q(w1578), .S(w1579), .R(w1584) );
	vdp_rs_ff g1689 (.Q(w1566), .R(w1558), .S(w1560) );
	vdp_rs_ff g1690 (.Q(w29), .S(w1588), .R(w1570) );
	vdp_rs_ff g1691 (.Q(w19), .R(w1561), .S(w1559) );
	vdp_tff g1692 (.C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .CI(w1576), .R(w1572), .A(w1567), .Q(ODD_EVEN) );
	vdp_cnt_bit_load g1693 (.D(w1770), .Q(w1637), .nL(w1882), .L(w1755), .CI(w1772), .nC1(nHCLK1), .CO(w1848), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g1694 (.Q(w1563), .D(HPLA13), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1695 (.Q(w1914), .D(HPLA0), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1696 (.Q(w30), .D(w1929), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1697 (.Q(w34), .D(HPLA14), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1698 (.Q(VRAM_REFRESH), .D(HPLA23), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1699 (.Q(w1638), .D(HPLA25), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1700 (.Q(w1633), .D(HPLA24), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1701 (.Q(w1609), .D(HPLA15), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1702 (.Q(w1634), .D(w1647), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1703 (.Q(w1597), .D(HPLA1), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1704 (.Q(w1778), .D(HPLA12), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1705 (.Q(w1661), .D(HPLA11), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1706 (.Q(w1779), .D(HPLA2), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1707 (.Q(w1647), .D(w1892), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1708 (.Q(w1788), .D(HPLA16), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1709 (.Q(w1642), .D(HPLA26), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1710 (.Q(w1660), .D(HPLA27), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1711 (.Q(w1927), .D(w1931), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1712 (.Q(w1694), .D(w1689), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1713 (.Q(w1644), .D(w1791), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1714 (.Q(w8), .D(HPLA28), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1715 (.Q(w1658), .D(HPLA17), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1716 (.Q(w1655), .D(w1837), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1717 (.Q(w1674), .D(HPLA10), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1718 (.Q(w1666), .D(HPLA3), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1719 (.Q(w1722), .D(w1670), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1720 (.Q(w27), .D(HPLA36), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1721 (.Q(w21), .D(HPLA29), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1722 (.Q(w1688), .D(HPLA18), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1723 (.Q(w1894), .D(w1728), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1724 (.Q(w1724), .D(HPLA9), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1725 (.Q(w1684), .D(HPLA4), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1726 (.Q(w1709), .D(HPLA35), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1727 (.Q(w28), .D(HPLA34), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1728 (.Q(w1711), .D(HPLA19), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1729 (.Q(w1712), .D(HPLA20), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1730 (.Q(w1737), .D(HPLA8), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1731 (.Q(w1685), .D(HPLA5), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1732 (.Q(w1602), .D(w1921), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1733 (.Q(w1672), .D(w1920), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1734 (.Q(w1723), .D(HPLA7), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1735 (.Q(w1686), .D(HPLA6), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1736 (.Q(w1727), .D(HPLA21), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1737 (.Q(w1706), .D(HPLA32), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1738 (.Q(w24), .D(HPLA31), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1739 (.Q(w1707), .D(w1602), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1740 (.Q(w1738), .D(w1695), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1741 (.Q(w1782), .D(HPLA22), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_not g1742 (.nZ(w1629), .A(M5) );
	vdp_not g1743 (.nZ(w6), .A(w1865) );
	vdp_not g1744 (.nZ(w35), .A(w1609) );
	vdp_not g1745 (.nZ(w1789), .A(w1606) );
	vdp_not g1746 (.nZ(w1613), .A(w50) );
	vdp_not g1747 (.nZ(w1615), .A(w1860) );
	vdp_not g1748 (.nZ(w1874), .A(w1) );
	vdp_not g1749 (.nZ(w1652), .A(w1625) );
	vdp_not g1750 (.nZ(w1635), .A(w1634) );
	vdp_not g1751 (.nZ(w1645), .A(w1609) );
	vdp_not g1752 (.nZ(w1646), .A(VSCR) );
	vdp_not g1753 (.nZ(w7), .A(w1640) );
	vdp_not g1754 (.nZ(w1631), .A(w36) );
	vdp_not g1755 (.nZ(w1926), .A(w50) );
	vdp_not g1756 (.nZ(w12), .A(w1888) );
	vdp_not g1757 (.nZ(w1889), .A(w1655) );
	vdp_not g1758 (.nZ(w1892), .A(w1665) );
	vdp_not g1759 (.nZ(w1699), .A(w1626) );
	vdp_not g1760 (.nZ(w1911), .A(w1624) );
	vdp_not g1761 (.nZ(w1650), .A(H40) );
	vdp_not g1762 (.nZ(w13), .A(w1697) );
	vdp_not g1763 (.nZ(w1881), .A(w1612) );
	vdp_not g1764 (.nZ(w1734), .A(w1668) );
	vdp_not g1765 (.nZ(w1713), .A(w1700) );
	vdp_not g1766 (.nZ(w1729), .A(w49) );
	vdp_not g1767 (.nZ(w1676), .A(w1833) );
	vdp_not g1768 (.nZ(w11), .A(w1866) );
	vdp_not g1769 (.nZ(w1741), .A(w1738) );
	vdp_not g1770 (.nZ(w1643), .A(w39) );
	vdp_not g1771 (.nZ(w1659), .A(w48) );
	vdp_not g1772 (.nZ(w1610), .A(w38) );
	vdp_not g1773 (.nZ(w1849), .A(w18) );
	vdp_not g1774 (.nZ(w1912), .A(w42) );
	vdp_not g1775 (.nZ(w1915), .A(M5) );
	vdp_not g1776 (.nZ(w1907), .A(w1677) );
	vdp_not g1777 (.nZ(w1754), .A(w1873) );
	vdp_not g1778 (.nZ(w1885), .A(w1858) );
	vdp_not g1779 (.nZ(w1756), .A(w1739) );
	vdp_not g1780 (.nZ(w1773), .A(w1771) );
	vdp_not g1781 (.nZ(w1767), .A(M2) );
	vdp_not g1782 (.nZ(w1768), .A(PAL) );
	vdp_aon22 g1783 (.Z(w1936), .B1(w1758), .A1(w1757), .A2(DB[4]), .B2(w1756) );
	vdp_aon22 g1784 (.Z(w1872), .B1(w1758), .A1(w1757), .A2(DB[5]), .B2(w1745) );
	vdp_aon22 g1785 (.Z(w1875), .B1(w1758), .A1(w1757), .B2(w1885), .A2(DB[6]) );
	vdp_aon22 g1786 (.Z(w1869), .B2(1'b1), .A2(DB[7]), .B1(w1758), .A1(w1757) );
	vdp_aon22 g1787 (.Z(w1868), .B2(1'b1), .A2(DB[8]), .B1(w1758), .A1(w1757) );
	vdp_aon22 g1788 (.Z(w1748), .B2(1'b1), .B1(w1611), .A2(DB[8]), .A1(w1930) );
	vdp_aon22 g1789 (.Z(w1884), .B2(w1744), .A2(DB[3]), .B1(w1758), .A1(w1757) );
	vdp_aon22 g1790 (.Z(w1765), .A2(DB[2]), .B2(w1768), .B1(w1758), .A1(w1757) );
	vdp_aon22 g1791 (.Z(w1766), .A2(DB[1]), .B2(w1743), .B1(w1758), .A1(w1757) );
	vdp_aon22 g1792 (.Z(w1876), .A1(w1930), .B1(w1611), .B2(1'b1), .A2(DB[7]) );
	vdp_aon22 g1793 (.Z(w20), .A1(w1915), .B2(w1746), .B1(M5), .A2(w1722) );
	vdp_aon22 g1794 (.Z(w1715), .B1(w1611), .A1(w1930), .A2(DB[6]), .B2(1'b1) );
	vdp_aon22 g1795 (.Z(w1693), .B1(w1707), .B2(w1708), .A2(w1783), .A1(w1705) );
	vdp_not g1796 (.nZ(w1708), .A(w1705) );
	vdp_aon22 g1797 (.Z(w1877), .B1(w1611), .A1(w1930), .B2(1'b0), .A2(DB[5]) );
	vdp_not g1798 (.nZ(w1735), .A(w1732) );
	vdp_aon22 g1799 (.Z(w1922), .B1(w1611), .A1(w1930), .B2(w1881), .A2(DB[4]) );
	vdp_aon22 g1800 (.Z(w1878), .B2(w1880), .B1(w1611), .A2(DB[3]), .A1(w1930) );
	vdp_aon22 g1801 (.Z(w1691), .A2(w1629), .B2(M5), .A1(w1693), .B1(w1692) );
	vdp_aon22 g1802 (.Z(w1879), .A2(DB[2]), .B2(w1662), .A1(w1930), .B1(w1611) );
	vdp_aon22 g1803 (.Z(w1890), .B2(w1788), .B1(VSCR), .A2(w1646), .A1(w1645) );
	vdp_aon22 g1804 (.Z(w1913), .B1(w1864), .A1(HCLK2), .B2(w1631), .A2(w36) );
	vdp_aon22 g1805 (.Z(w1905), .A1(w1930), .B1(w1611), .B2(w1648), .A2(DB[1]) );
	vdp_aon22 g1806 (.Z(w1616), .A2(DB[0]), .B1(w1611), .B2(w1612), .A1(w1930) );
	vdp_not g1807 (.nZ(w4), .A(w1778) );
	vdp_not g1808 (.nZ(w3), .A(w1644) );
	vdp_rs_ff g1809 (.Q(w1687), .S(w1736), .R(w1852) );
	vdp_rs_ff g1810 (.Q(w1733), .R(w1724), .S(w1726) );
	vdp_rs_ff g1811 (.Q(w1670), .S(w1895), .R(w1686) );
	vdp_rs_ff g1812 (.Q(w1851), .R(w1925), .S(w1666) );
	vdp_rs_ff g1813 (.Q(w1671), .R(w1661), .S(w1919) );
	vdp_aon22 g1814 (.Z(w1770), .A2(DB[0]), .B2(w1742), .B1(w1758), .A1(w1757) );
	vdp_notif0 g1815 (.nZ(DB[1]), .A(VRAM_REFRESH), .nE(w1627) );
	vdp_notif0 g1816 (.nZ(DB[0]), .A(w30), .nE(w1627) );
	vdp_notif0 g1817 (.nZ(DB[7]), .A(w34), .nE(w1628) );
	vdp_notif0 g1818 (.A(w35), .nZ(DB[6]), .nE(w1628) );
	vdp_notif0 g1819 (.A(w6), .nZ(DB[2]), .nE(w1627) );
	vdp_notif0 g1820 (.A(w7), .nZ(DB[3]), .nE(w1627) );
	vdp_notif0 g1821 (.nZ(DB[5]), .A(w13), .nE(w1627) );
	vdp_notif0 g1822 (.A(w12), .nZ(DB[4]), .nE(w1627) );
	vdp_notif0 g1823 (.A(w15), .nZ(DB[5]), .nE(w1628) );
	vdp_notif0 g1824 (.nZ(DB[7]), .A(w8), .nE(w1627) );
	vdp_notif0 g1825 (.nZ(DB[6]), .A(w3), .nE(w1627) );
	vdp_notif0 g1826 (.nZ(DB[4]), .A(w16), .nE(w1628) );
	vdp_notif0 g1827 (.nZ(DB[9]), .A(w27), .nE(w1627) );
	vdp_notif0 g1828 (.nZ(DB[8]), .A(w21), .nE(w1627) );
	vdp_notif0 g1829 (.nZ(DB[3]), .A(w10), .nE(w1628) );
	vdp_notif0 g1830 (.nZ(DB[2]), .A(w26), .nE(w1628) );
	vdp_notif0 g1831 (.nZ(DB[10]), .A(w28), .nE(w1627) );
	vdp_notif0 g1832 (.nZ(DB[11]), .A(w11), .nE(w1627) );
	vdp_notif0 g1833 (.nZ(DB[12]), .A(w23), .nE(w1627) );
	vdp_notif0 g1834 (.nZ(DB[13]), .A(w24), .nE(w1627) );
	vdp_notif0 g1835 (.nZ(DB[1]), .A(w14), .nE(w1628) );
	vdp_notif0 g1836 (.nZ(DB[0]), .A(w9), .nE(w1628) );
	vdp_not g1837 (.nZ(VPOS[9]), .A(w1871) );
	vdp_not g1838 (.nZ(VPOS[8]), .A(w1870) );
	vdp_not g1839 (.nZ(VPOS[7]), .A(w1679) );
	vdp_not g1840 (.nZ(HPOS[7]), .A(w1907) );
	vdp_not g1841 (.nZ(HPOS[8]), .A(w1754) );
	vdp_not g1842 (.nZ(HPOS[6]), .A(w1676) );
	vdp_not g1843 (.nZ(VPOS[6]), .A(w1908) );
	vdp_not g1844 (.nZ(VPOS[5]), .A(w1909) );
	vdp_not g1845 (.nZ(HPOS[5]), .A(w1713) );
	vdp_not g1846 (.nZ(HPOS[4]), .A(w1734) );
	vdp_not g1847 (.nZ(VPOS[4]), .A(w1910) );
	vdp_not g1848 (.nZ(HPOS[3]), .A(w1911) );
	vdp_not g1849 (.nZ(VPOS[3]), .A(w1663) );
	vdp_not g1850 (.nZ(HPOS[2]), .A(w1699) );
	vdp_not g1851 (.nZ(VPOS[2]), .A(w1653) );
	vdp_not g1852 (.nZ(HPOS[1]), .A(w1652) );
	vdp_not g1853 (.nZ(VPOS[1]), .A(w1614) );
	vdp_not g1854 (.nZ(HPOS[0]), .A(w1615) );
	vdp_not g1855 (.nZ(VPOS[0]), .A(w1608) );
	vdp_aoi22 g1856 (.Z(w1864), .A1(w1603), .B1(w1630), .B2(M5), .A2(w1629) );
	vdp_aon22 g1857 (.Z(w1654), .A2(w1629), .B1(w1690), .B2(M5), .A1(w1695) );
	vdp_aoi22 g1858 (.Z(w1608), .B2(w1874), .B1(w1637), .A1(ODD_EVEN), .A2(w1) );
	vdp_aoi22 g1859 (.Z(w1614), .B2(w1874), .B1(w1775), .A1(w1637), .A2(w1) );
	vdp_aoi22 g1860 (.Z(w1653), .A2(w1), .A1(w1775), .B2(w1874), .B1(w1857) );
	vdp_aoi22 g1861 (.Z(w1663), .A1(w1857), .B2(w1874), .A2(w1), .B1(w1760) );
	vdp_aoi22 g1862 (.Z(w1910), .B1(w1856), .A1(w1760), .A2(w1), .B2(w1874) );
	vdp_aoi22 g1863 (.Z(w1909), .B1(w1855), .A1(w1856), .A2(w1), .B2(w1874) );
	vdp_aoi22 g1864 (.Z(w1908), .A2(w1), .B2(w1874), .B1(w1680), .A1(w1855) );
	vdp_aoi22 g1865 (.Z(w1679), .B2(w1874), .A1(w1680), .B1(w1854), .A2(w1) );
	vdp_aoi22 g1866 (.Z(w1870), .B2(w1874), .A2(w1), .A1(w1854), .B1(w1777) );
	vdp_aoi22 g1867 (.Z(w1871), .B1(1'b0), .A2(w1), .B2(w1874), .A1(w1777) );
	vdp_comp_dff g1868 (.Q(w1598), .D(w1632), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_comp_dff g1869 (.Q(w1730), .D(w1896), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_cnt_bit g1870 (.CI(w1898), .Q(w1783), .R(SYSRES), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g1871 (.nZ(w1867), .A(w52) );
	vdp_and g1872 (.Z(w1717), .A(w1732), .B(w1671) );
	vdp_and g1873 (.Z(w1718), .A(w1732), .B(w1671) );
	vdp_and g1874 (.Z(w1720), .A(w1924), .B(w1733) );
	vdp_and g1875 (.Z(w1721), .A(w1733), .B(w1735) );
	vdp_and g1876 (.Z(w1719), .A(w1781), .B(w1687) );
	vdp_and g1877 (.Z(w1924), .A(w1780), .B(w1669) );
	vdp_and g1878 (.Z(w1662), .A(w50), .B(w1650) );
	vdp_and g1879 (.Z(w15), .A(w1890), .B(w1641) );
	vdp_and g1880 (.Z(w1648), .A(w1613), .B(w1650) );
	vdp_and g1881 (.Z(w25), .A(w1583), .B(w1851) );
	vdp_and g1882 (.Z(w1649), .A(w49), .B(w1730) );
	vdp_and g1883 (.Z(w1673), .A(w1849), .B(w50) );
	vdp_and g1884 (.Z(w14), .A(w1641), .B(w1727) );
	vdp_and g1885 (.Z(w1862), .A(w1912), .B(w1673) );
	vdp_and g1886 (.Z(w9), .A(w1782), .B(w1641) );
	vdp_and g1887 (.Z(w1883), .A(w1740), .B(w4) );
	vdp_or g1888 (.Z(w1745), .A(w1853), .B(w1858) );
	vdp_or g1889 (.Z(w1744), .A(w1886), .B(w1858) );
	vdp_and g1890 (.Z(w1705), .A(M5), .B(w22) );
	vdp_and g1891 (.Z(w1898), .A(w1741), .B(w1695) );
	vdp_or g1892 (.Z(w1726), .A(w1725), .B(SYSRES) );
	vdp_or g1893 (.Z(w26), .A(w1712), .B(w1711) );
	vdp_or g1894 (.Z(w23), .A(w1706), .B(w1712) );
	vdp_or g1895 (.Z(w1921), .A(w1717), .B(w1721) );
	vdp_or g1896 (.Z(w1736), .A(w1723), .B(w1684) );
	vdp_or g1897 (.Z(w1852), .A(SYSRES), .B(w1725) );
	vdp_or g1898 (.Z(w1725), .A(w1674), .B(w1737) );
	vdp_or g1899 (.Z(w1895), .A(w1685), .B(SYSRES) );
	vdp_or g1900 (.Z(w1880), .A(w1612), .B(w1923) );
	vdp_or g1901 (.Z(w1925), .A(SYSRES), .B(w1684) );
	vdp_or g1902 (.Z(w1893), .A(w1649), .B(w1598) );
	vdp_or g1903 (.Z(w1837), .A(w1894), .B(w1728) );
	vdp_and g1904 (.Z(w10), .A(w1641), .B(w1688) );
	vdp_and g1905 (.Z(w1728), .A(w1604), .B(w1673) );
	vdp_or g1906 (.Z(w1919), .A(SYSRES), .B(w1674) );
	vdp_not g1907 (.nZ(w1628), .A(w51) );
	vdp_not g1908 (.nZ(w1627), .A(w45) );
	vdp_aon33 g1909 (.Z(w1772), .A3(w1771), .A2(w1867), .A1(w4), .B1(w52), .B3(1'b1), .B2(w1188) );
	vdp_aoi21 g1910 (.Z(w1865), .A1(w1633), .A2(w1641), .B(w1605) );
	vdp_aoi21 g1911 (.Z(w1640), .A1(w1638), .B(w1639), .A2(w1641) );
	vdp_aoi21 g1912 (.Z(w1606), .A1(w37), .A2(w47), .B(w1636) );
	vdp_aoi21 g1913 (.Z(w1665), .A1(w1647), .B(w1891), .A2(w1893) );
	vdp_aoi21 g1914 (.Z(w1888), .A1(w1641), .B(w1887), .A2(w1642) );
	vdp_aoi21 g1915 (.Z(w1697), .B(w1897), .A1(w1641), .A2(w1660) );
	vdp_aoi21 g1916 (.Z(w1866), .A1(w1641), .A2(w1709), .B(w1710) );
	vdp_xor g1917 (.Z(w1695), .B(w1603), .A(w1672) );
	vdp_xor g1918 (.Z(w1742), .A(ODD_EVEN), .B(w1768) );
	vdp_and3 g1919 (.Z(w1605), .A(w1659), .B(w39), .C(w1610) );
	vdp_and3 g1920 (.Z(w1929), .A(w1928), .B(w1787), .C(w1656) );
	vdp_and3 g1921 (.Z(w1639), .A(w1643), .B(w48), .C(w1610) );
	vdp_and3 g1922 (.Z(w1887), .A(w48), .B(w1610), .C(w39) );
	vdp_and3 g1923 (.Z(w1897), .A(w1643), .B(w1659), .C(w1712) );
	vdp_and3 g1924 (.Z(w1710), .A(w39), .B(w1659), .C(w38) );
	vdp_or3 g1925 (.Z(w1920), .A(w1719), .B(w1720), .C(w1718) );
	vdp_and3 g1926 (.Z(w1923), .A(w50), .B(w1650), .C(M5) );
	vdp_and3 g1927 (.Z(w1798), .A(w1647), .B(w50), .C(w1635) );
	vdp_and3 g1928 (.Z(w1612), .A(H40), .B(M5), .C(w1613) );
	vdp_nor4 g1929 (.Z(w1656), .A(HPLA33), .B(HPLA35), .C(HPLA29), .D(HPLA36) );
	vdp_nor4 g1930 (.Z(w1771), .A(w53), .B(w1774), .D(w1883), .C(SYSRES) );
	vdp_comp_we g1931 (.Z(w1755), .nZ(w1882), .A(w1773) );
	vdp_comp_we g1932 (.Z(w1757), .nZ(w1758), .A(w53) );
	vdp_comp_we g1933 (.Z(w1930), .nZ(w1611), .A(w54) );
	vdp_comp_we g1934 (.Z(w1618), .nZ(w1617), .A(w1604) );
	vdp_and3 g1935 (.Z(w17), .A(DISP), .B(w1851), .C(w29) );
	vdp_or4 g1936 (.Z(w1604), .A(w54), .B(SYSRES), .C(w1798), .D(w1914) );
	vdp_nor3 g1937 (.Z(w1787), .A(HPLA28), .B(HPLA30), .C(HPLA27) );
	vdp_nor3 g1938 (.Z(w1732), .A(w1669), .B(w1781), .C(w1780) );
	vdp_nand g1939 (.Z(w1689), .A(w1691), .B(w1729) );
	vdp_nand g1940 (.Z(w1931), .A(w1654), .B(w1926) );
	vdp_nand g1941 (.Z(w1791), .A(w1889), .B(HPLA30) );
	vdp_nor3 g1942 (.Z(w1641), .A(w39), .B(w48), .C(w38) );
	vdp_nor g1943 (.Z(w1858), .A(w1768), .B(M5) );
	vdp_nor g1944 (.Z(w1743), .A(ODD_EVEN), .B(w1768) );
	vdp_nor g1945 (.Z(w1853), .A(w1756), .B(PAL) );
	vdp_nor g1946 (.Z(w1886), .A(w1756), .B(w1768) );
	vdp_nor g1947 (.Z(w1891), .A(w1597), .B(SYSRES) );
	vdp_sdelay8 g1948 (.Q(w1746), .D(w1722), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2), .nC3(nHCLK1), .C3(HCLK1), .nC4(nHCLK2), .C4(HCLK2), .nC5(nHCLK1), .C5(HCLK1), .nC6(nHCLK2), .C6(HCLK2), .nC7(nHCLK1), .C7(HCLK1), .nC8(nHCLK2), .C8(HCLK2), .nC9(nHCLK1), .C9(HCLK1), .nC10(nHCLK2), .C10(HCLK2), .nC11(nHCLK1), .C11(HCLK1), .nC12(nHCLK2), .C12(HCLK2), .nC13(nHCLK1), .C13(HCLK1), .nC14(nHCLK2), .C14(HCLK2), .nC15(nHCLK1), .C15(HCLK1), .nC16(nHCLK2), .C16(HCLK2) );
	vdp_sdelay7 g1949 (.Q(w1692), .D(w1693), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .nC4(nHCLK2), .C5(HCLK1), .nC5(nHCLK1), .C6(HCLK2), .nC6(nHCLK2), .C7(HCLK1), .nC7(nHCLK1), .C8(HCLK2), .nC8(nHCLK2), .C9(HCLK1), .nC9(nHCLK1), .C10(HCLK2), .nC10(nHCLK2), .C11(HCLK1), .nC11(nHCLK1), .C12(HCLK2), .nC12(nHCLK2), .C13(HCLK1), .nC13(nHCLK1), .C14(HCLK2), .nC14(nHCLK2), .C3(HCLK1) );
	vdp_sdelay8 g1950 (.Q(w1690), .D(w1695), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2), .C3(HCLK1), .nC4(nHCLK2), .C4(HCLK2), .nC5(nHCLK1), .C5(HCLK1), .nC6(nHCLK2), .C6(HCLK2), .nC7(nHCLK1), .C7(HCLK1), .nC8(nHCLK2), .C8(HCLK2), .nC9(nHCLK1), .C9(HCLK1), .nC10(nHCLK2), .C10(HCLK2), .C11(HCLK1), .nC12(nHCLK2), .C12(HCLK2), .nC13(nHCLK1), .C13(HCLK1), .nC14(nHCLK2), .C14(HCLK2), .nC15(nHCLK1), .C15(HCLK1), .nC16(nHCLK2), .C16(HCLK2), .nC3(nHCLK1), .nC11(nHCLK1) );
	vdp_sdelay8 g1951 (.Q(w1630), .D(w1603), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2), .C3(HCLK1), .nC4(nHCLK2), .C4(HCLK2), .nC5(nHCLK1), .C5(HCLK1), .nC6(nHCLK2), .C6(HCLK2), .nC7(nHCLK1), .C7(HCLK1), .nC8(nHCLK2), .C8(HCLK2), .nC9(nHCLK1), .C9(HCLK1), .nC10(nHCLK2), .C10(HCLK2), .nC11(nHCLK1), .C11(HCLK1), .nC12(nHCLK2), .C12(HCLK2), .nC13(nHCLK1), .C13(HCLK1), .nC14(nHCLK2), .C14(HCLK2), .nC15(nHCLK1), .C15(HCLK1), .nC16(nHCLK2), .C16(HCLK2), .nC3(nHCLK1) );
	vdp_cnt_bit_load g1952 (.D(w1766), .Q(w1775), .nL(w1882), .L(w1755), .CI(w1848), .nC1(nHCLK1), .CO(w1933), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1953 (.D(w1765), .Q(w1857), .nL(w1882), .L(w1755), .CI(w1933), .nC1(nHCLK1), .CO(w1934), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1954 (.D(w1884), .Q(w1760), .nL(w1882), .L(w1755), .CI(w1934), .nC1(nHCLK1), .CO(w1935), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1955 (.D(w1936), .Q(w1856), .nL(w1882), .L(w1755), .CI(w1935), .nC1(nHCLK1), .CO(w1786), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1956 (.D(w1872), .Q(w1855), .nL(w1882), .L(w1755), .CI(w1786), .nC1(nHCLK1), .CO(w1785), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1957 (.D(w1875), .Q(w1680), .nL(w1882), .L(w1755), .CI(w1785), .nC1(nHCLK1), .CO(w1937), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1958 (.D(w1869), .Q(w1854), .nL(w1882), .L(w1755), .CI(w1937), .nC1(nHCLK1), .CO(w1784), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1959 (.D(w1868), .Q(w1777), .nL(w1882), .L(w1755), .CI(w1784), .nC1(nHCLK1), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1960 (.D(w1748), .Q(w1873), .nL(w1617), .L(w1618), .CI(w1749), .nC1(nHCLK1), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1961 (.D(w1876), .Q(w1677), .nL(w1617), .L(w1618), .CI(w1675), .nC1(nHCLK1), .CO(w1749), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1962 (.D(w1715), .Q(w1833), .nL(w1617), .L(w1618), .CI(w1714), .nC1(nHCLK1), .CO(w1675), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1963 (.D(w1877), .Q(w1700), .nL(w1617), .L(w1618), .CI(w1701), .nC1(nHCLK1), .CO(w1714), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1964 (.D(w1922), .Q(w1668), .nL(w1617), .L(w1618), .CI(w1667), .nC1(nHCLK1), .CO(w1701), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1965 (.D(w1878), .Q(w1624), .nL(w1617), .L(w1618), .CI(w1664), .nC1(nHCLK1), .CO(w1667), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1966 (.D(w1879), .Q(w1626), .nL(w1617), .L(w1618), .CI(w1651), .nC1(nHCLK1), .CO(w1664), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1967 (.D(w1905), .Q(w1625), .nL(w1617), .L(w1618), .CI(w1932), .nC1(nHCLK1), .CO(w1651), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1968 (.D(w1616), .Q(w1860), .nL(w1617), .L(w1618), .CI(w1789), .nC1(nHCLK1), .CO(w1932), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_or8 g1969 (.Z(VPLA7), .A(w1799), .B(w1800), .C(w1801), .D(w1802), .E(w1845), .F(w1846), .G(w1847), .H(w1803) );
	vdp_or8 g1970 (.Z(VPLA6), .A(w1804), .B(w1844), .C(w1843), .D(w1826), .E(w1842), .F(w1805), .G(w1806), .H(w1841) );
	vdp_or8 g1971 (.Z(VPLA5), .A(w1938), .B(w1917), .C(w1918), .D(w1903), .E(w1825), .F(w1824), .G(w1902), .H(w1823) );
	vdp_or5 g1972 (.Z(VPLA4), .A(w1819), .B(w1820), .C(w1821), .D(w1822), .E(w6537) );
	vdp_or7 g1973 (.Z(VPLA3), .A(w6614), .B(w6615), .C(w6613), .D(w1818), .E(w6534), .F(w6535), .G(w6536) );
	vdp_or7 g1974 (.Z(VPLA0), .A(w1807), .B(w1808), .C(w1809), .D(w1810), .E(w1811), .F(w1812), .G(w1813) );
	vdp_nor g1975 (.Z(w1636), .A(w1604), .B(w37) );
	vdp_and g1976 (.Z(w16), .A(w1641), .B(w1658) );
	vdp_not g1977 (.nZ(VPLA1), .A(w1814) );
	vdp_nor3 g1978 (.Z(VPLA2), .A(w1817), .B(w1816), .C(w1815) );
	vdp_rs_ff g1979 (.S(w1850), .R(w1579), .Q(w1577) );
	vdp_rs_ff g1980 (.S(w1591), .R(w1587), .Q(w1575) );
	vdp_and g1981 (.Z(w1780), .A(w1566), .B(M5) );
	vdp_nor4 g1982 (.Z(w1928), .A(HPLA23), .B(HPLA25), .C(HPLA24), .D(HPLA26) );
	vdp_nand3 g1983 (.A(w2059), .B(w2058), .C(w2056), .Z(w2052) );
	vdp_nand3 g1984 (.A(w2056), .B(w2058), .C(w2061), .Z(w2047) );
	vdp_nand3 g1985 (.A(w2056), .B(w2059), .C(w2060), .Z(w2048) );
	vdp_nand3 g1986 (.A(w2060), .B(w2056), .C(w2061), .Z(w2049) );
	vdp_nand3 g1987 (.A(w2060), .B(w2057), .C(w2061), .Z(w2044) );
	vdp_nand3 g1988 (.A(w2057), .B(w2059), .C(w2060), .Z(w2043) );
	vdp_nand3 g1989 (.A(w2058), .B(w2057), .C(w2061), .Z(w2051) );
	vdp_nand3 g1990 (.A(w2059), .B(w2058), .C(w2057), .Z(w2050) );
	vdp_nand3 g1991 (.A(w2032), .B(w2033), .C(w2028), .Z(w2042) );
	vdp_nand3 g1992 (.A(w2028), .B(w2033), .C(w2031), .Z(w2041) );
	vdp_nand3 g1993 (.A(w2030), .B(w2029), .C(w2031), .Z(w2035) );
	vdp_nand3 g1994 (.A(w2029), .B(w2032), .C(w2030), .Z(w2036) );
	vdp_nand3 g1995 (.A(w2033), .B(w2029), .C(w2031), .Z(w2037) );
	vdp_nand3 g1996 (.A(w2032), .B(w2033), .C(w2029), .Z(w2038) );
	vdp_nand3 g1997 (.A(w2030), .B(w2028), .C(w2031), .Z(w2039) );
	vdp_nand3 g1998 (.A(w2028), .B(w2032), .C(w2030), .Z(w2040) );
	vdp_nand3 g1999 (.A(w2020), .B(w2018), .C(w2016), .Z(w2013) );
	vdp_nand3 g2000 (.A(w2016), .B(w2018), .C(w2021), .Z(w2012) );
	vdp_nand3 g2001 (.A(w2019), .B(w2017), .C(w2021), .Z(w2006) );
	vdp_nand3 g2002 (.A(w2017), .B(w2020), .C(w2019), .Z(w2007) );
	vdp_nand3 g2003 (.A(w2018), .B(w2017), .C(w2021), .Z(w2008) );
	vdp_nand3 g2004 (.A(w2020), .B(w2018), .C(w2017), .Z(w2009) );
	vdp_nand3 g2005 (.A(w2019), .B(w2016), .C(w2021), .Z(w2010) );
	vdp_nand3 g2006 (.A(w2016), .B(w2020), .C(w2019), .Z(w2011) );
	vdp_nand3 g2007 (.A(w1959), .B(w1956), .C(w1960), .Z(w1953) );
	vdp_nand3 g2008 (.A(w1960), .B(w1956), .C(w1958), .Z(w1952) );
	vdp_nand3 g2009 (.A(w1957), .B(w1955), .C(w1958), .Z(w1946) );
	vdp_nand3 g2010 (.A(w1955), .B(w1959), .C(w1957), .Z(w1947) );
	vdp_nand3 g2011 (.A(w1956), .B(w1955), .C(w1958), .Z(w1948) );
	vdp_nand3 g2012 (.A(w1959), .B(w1956), .C(w1955), .Z(w1949) );
	vdp_nand3 g2013 (.A(w1957), .B(w1960), .C(w1958), .Z(w1950) );
	vdp_nand3 g2014 (.A(w1960), .B(w1959), .C(w1957), .Z(w1951) );
	vdp_not g2015 (.nZ(w1954), .A(w1941) );
	vdp_not g2016 (.nZ(w2014), .A(w1942) );
	vdp_not g2017 (.nZ(w2022), .A(w1939) );
	vdp_not g2018 (.nZ(w2053), .A(w1940) );
	vdp_nand g2019 (.Z(w1944), .B(w1945), .A(w1954) );
	vdp_nand g2020 (.Z(w1945), .B(w1954), .A(w1961) );
	vdp_nand g2021 (.Z(w2004), .B(w2005), .A(w2014) );
	vdp_nand g2022 (.Z(w2005), .B(w2014), .A(w1965) );
	vdp_comp_we g2023 (.A(w2015), .Z(w2017), .nZ(w2016) );
	vdp_comp_we g2024 (.A(w2075), .Z(w2019), .nZ(w2018) );
	vdp_comp_we g2025 (.A(w2074), .Z(w2021), .nZ(w2020) );
	vdp_comp_we g2026 (.A(w1962), .Z(w1955), .nZ(w1960) );
	vdp_comp_we g2027 (.A(w1963), .Z(w1957), .nZ(w1956) );
	vdp_comp_we g2028 (.A(w1964), .Z(w1958), .nZ(w1959) );
	vdp_nand g2029 (.Z(w2023), .B(w2022), .A(w2026) );
	vdp_comp_we g2030 (.A(w2025), .Z(w2029), .nZ(w2028) );
	vdp_comp_we g2031 (.A(w2027), .Z(w2030), .nZ(w2033) );
	vdp_comp_we g2032 (.A(w2034), .Z(w2031), .nZ(w2032) );
	vdp_nand g2033 (.Z(w2024), .B(w2023), .A(w2022) );
	vdp_nand g2034 (.Z(w2045), .B(w2053), .A(w2054) );
	vdp_comp_we g2035 (.A(w2055), .Z(w2057), .nZ(w2056) );
	vdp_comp_we g2036 (.A(w2062), .Z(w2060), .nZ(w2058) );
	vdp_comp_we g2037 (.A(w2063), .Z(w2061), .nZ(w2059) );
	vdp_nand g2038 (.Z(w2046), .B(w2045), .A(w2053) );
	vdp_comp_str g2039 (.A(w2086), .Z(w2087), .nZ(w2085) );
	vdp_comp_str g2040 (.A(w2103), .Z(w2076), .nZ(w2077) );
	vdp_comp_str g2041 (.A(w2112), .Z(w2067), .nZ(w2066) );
	vdp_comp_str g2042 (.A(w2113), .Z(w1968), .nZ(w1967) );
	vdp_comp_str g2043 (.A(w1976), .Z(w1977), .nZ(w1978) );
	vdp_comp_str g2044 (.A(w2150), .Z(w2336), .nZ(w2213) );
	vdp_comp_str g2045 (.A(w2361), .Z(w2329), .nZ(w2328) );
	vdp_comp_str g2046 (.A(w2332), .Z(w2342), .nZ(w2330) );
	vdp_comp_str g2047 (.A(w2121), .Z(w2333), .nZ(w2331) );
	vdp_comp_str g2048 (.A(w2241), .Z(w1984), .nZ(w1988) );
	vdp_comp_str g2049 (.A(w2362), .Z(w1985), .nZ(w1989) );
	vdp_comp_str g2050 (.A(w2119), .Z(w1987), .nZ(w1990) );
	vdp_slatch g2051 (.Q(w2346), .C(w1987), .D(w2114), .nC(w1990) );
	vdp_slatch g2052 (.Q(w2345), .C(w1985), .D(w2114), .nC(w1989) );
	vdp_slatch g2053 (.Q(w2308), .C(w1987), .D(w2248), .nC(w1990) );
	vdp_slatch g2054 (.Q(w2344), .C(w1984), .D(w2114), .nC(w1988) );
	vdp_slatch g2055 (.Q(w2349), .C(w1987), .D(w2249), .nC(w1990) );
	vdp_slatch g2056 (.Q(w2307), .C(w1984), .D(w2248), .nC(w1988) );
	vdp_slatch g2057 (.Q(w2309), .C(w1985), .D(w2248), .nC(w1989) );
	vdp_slatch g2058 (.Q(w2243), .C(w1987), .D(w2251), .nC(w1990) );
	vdp_slatch g2059 (.Q(w2347), .C(w1984), .D(w2249), .nC(w1988) );
	vdp_slatch g2060 (.Q(w2348), .C(w1985), .D(w2249), .nC(w1989) );
	vdp_slatch g2061 (.Q(w1997), .C(w1987), .D(w1986), .nC(w1990) );
	vdp_slatch g2062 (.Q(w2242), .C(w1984), .D(w2251), .nC(w1988) );
	vdp_slatch g2063 (.Q(w2244), .C(w1985), .D(w2251), .nC(w1989) );
	vdp_slatch g2064 (.Q(w1994), .C(w1984), .D(w1986), .nC(w1988) );
	vdp_slatch g2065 (.Q(w1996), .C(w1985), .D(w1986), .nC(w1989) );
	vdp_slatch g2066 (.Q(w1991), .C(w1987), .D(w1983), .nC(w1990) );
	vdp_slatch g2067 (.Q(w2003), .C(w1984), .D(w1983), .nC(w1988) );
	vdp_slatch g2068 (.Q(w1992), .C(w1985), .D(w1983), .nC(w1989) );
	vdp_slatch g2069 (.Q(w2322), .C(w2333), .D(w2114), .nC(w2331) );
	vdp_slatch g2070 (.Q(w2321), .C(w2342), .D(w2114), .nC(w2330) );
	vdp_slatch g2071 (.Q(w2327), .C(w2333), .D(w2248), .nC(w2331) );
	vdp_slatch g2072 (.Q(w2323), .C(w2329), .D(w2114), .nC(w2328) );
	vdp_slatch g2073 (.Q(w2315), .C(w2333), .D(w2249), .nC(w2331) );
	vdp_slatch g2074 (.Q(w2325), .C(w2329), .D(w2248), .nC(w2328) );
	vdp_slatch g2075 (.Q(w2326), .C(w2342), .D(w2248), .nC(w2330) );
	vdp_slatch g2076 (.Q(w2312), .C(w2333), .D(w2251), .nC(w2331) );
	vdp_slatch g2077 (.Q(w2313), .C(w2329), .D(w2249), .nC(w2328) );
	vdp_slatch g2078 (.Q(w2314), .C(w2342), .D(w2249), .nC(w2330) );
	vdp_slatch g2079 (.Q(w2310), .C(w2329), .D(w2251), .nC(w2328) );
	vdp_slatch g2080 (.Q(w2311), .C(w2342), .D(w2251), .nC(w2330) );
	vdp_slatch g2081 (.Q(w2197), .C(w2336), .D(w2249), .nC(w2213) );
	vdp_slatch g2082 (.Q(w2339), .C(w2336), .D(w2248), .nC(w2213) );
	vdp_slatch g2083 (.Q(w2340), .C(w2336), .D(w2114), .nC(w2213) );
	vdp_and g2084 (.Z(w2157), .A(w2340), .B(w2339) );
	vdp_and g2085 (.Z(w2324), .A(w2339), .B(w2337) );
	vdp_and g2086 (.Z(w2306), .A(w2340), .B(w2338) );
	vdp_and g2087 (.Z(w2252), .A(w2337), .B(w2338) );
	vdp_slatch g2088 (.Q(w2089), .C(w2087), .D(w2083), .nC(w2085) );
	vdp_or g2089 (.Z(w2063), .A(w2088), .B(w2089) );
	vdp_notif0 g2090 (.A(w2063), .nZ(DB[0]), .nE(w1969) );
	vdp_slatch g2091 (.Q(w2364), .C(w2087), .D(w2080), .nC(w2085) );
	vdp_or g2092 (.Z(w2062), .A(w2088), .B(w2364) );
	vdp_notif0 g2093 (.A(w2062), .nZ(DB[1]), .nE(w1969) );
	vdp_slatch g2094 (.Q(w2365), .C(w2087), .D(w2082), .nC(w2085) );
	vdp_or g2095 (.Z(w2055), .A(w2088), .B(w2365) );
	vdp_notif0 g2096 (.A(w2055), .nZ(DB[2]), .nE(w1969) );
	vdp_slatch g2097 (.Q(w2093), .C(w2087), .D(w2094), .nC(w2085) );
	vdp_or g2098 (.Z(w2054), .A(w2088), .B(w2093) );
	vdp_notif0 g2099 (.A(w2054), .nZ(DB[3]), .nE(w1969) );
	vdp_slatch g2100 (.Q(w2084), .C(w2076), .D(w2083), .nC(w2077) );
	vdp_or g2101 (.Z(w2034), .A(w2081), .B(w2084) );
	vdp_notif0 g2102 (.A(w2034), .nZ(DB[4]), .nE(w1969) );
	vdp_slatch g2103 (.Q(w2079), .C(w2076), .D(w2080), .nC(w2077) );
	vdp_or g2104 (.Z(w2027), .A(w2081), .B(w2079) );
	vdp_notif0 g2105 (.A(w2027), .nZ(DB[5]), .nE(w1969) );
	vdp_slatch g2106 (.Q(w2078), .C(w2076), .D(w2082), .nC(w2077) );
	vdp_or g2107 (.Z(w2025), .A(w2081), .B(w2078) );
	vdp_notif0 g2108 (.A(w2025), .nZ(DB[6]), .nE(w1969) );
	vdp_slatch g2109 (.Q(w2073), .C(w2076), .D(w2094), .nC(w2077) );
	vdp_or g2110 (.Z(w2026), .A(w2081), .B(w2073) );
	vdp_notif0 g2111 (.A(w2026), .nZ(DB[7]), .nE(w1969) );
	vdp_slatch g2112 (.Q(w2363), .C(w2067), .D(w2083), .nC(w2066) );
	vdp_or g2113 (.Z(w2074), .A(w2068), .B(w2363) );
	vdp_notif0 g2114 (.A(w2074), .nZ(DB[8]), .nE(w1969) );
	vdp_slatch g2115 (.Q(w2072), .C(w2067), .D(w2080), .nC(w2066) );
	vdp_or g2116 (.Z(w2075), .A(w2068), .B(w2072) );
	vdp_notif0 g2117 (.A(w2075), .nZ(DB[9]), .nE(w1969) );
	vdp_slatch g2118 (.Q(w2065), .C(w2067), .D(w2082), .nC(w2066) );
	vdp_or g2119 (.Z(w2015), .A(w2068), .B(w2065) );
	vdp_notif0 g2120 (.A(w2015), .nZ(DB[10]), .nE(w1969) );
	vdp_slatch g2121 (.Q(w2064), .C(w2067), .D(w2094), .nC(w2066) );
	vdp_or g2122 (.Z(w1965), .A(w2068), .B(w2064) );
	vdp_notif0 g2123 (.A(w1965), .nZ(DB[11]), .nE(w1969) );
	vdp_slatch g2124 (.Q(w1970), .C(w1968), .D(w2083), .nC(w1967) );
	vdp_or g2125 (.Z(w1964), .A(w1966), .B(w1970) );
	vdp_notif0 g2126 (.A(w1964), .nZ(DB[12]), .nE(w1969) );
	vdp_slatch g2127 (.Q(w1971), .C(w1968), .D(w2080), .nC(w1967) );
	vdp_or g2128 (.Z(w1963), .A(w1966), .B(w1971) );
	vdp_notif0 g2129 (.A(w1963), .nZ(DB[13]), .nE(w1969) );
	vdp_slatch g2130 (.Q(w1972), .C(w1968), .D(w2082), .nC(w1967) );
	vdp_or g2131 (.Z(w1962), .A(w1966), .B(w1972) );
	vdp_notif0 g2132 (.A(w1962), .nZ(DB[14]), .nE(w1969) );
	vdp_slatch g2133 (.Q(w1973), .C(w1968), .D(w2094), .nC(w1967) );
	vdp_or g2134 (.Z(w1961), .A(w1966), .B(w1973) );
	vdp_notif0 g2135 (.A(w1961), .nZ(DB[15]), .nE(w1969) );
	vdp_not g2136 (.A(PSG_TEST_OE), .nZ(w1969) );
	vdp_not g2137 (.nZ(w2142), .A(PSG_Z80_CLK) );
	vdp_clkgen g2138 (.PH(w2142), .CLK1(w2143), .nCLK1(w2144), .CLK2(w2145), .nCLK2(w2146) );
	vdp_comp_dff g2139 (.D(SYSRES), .nC1(w2144), .C1(w2143), .C2(w2145), .nC2(w2146), .Q(w2174) );
	vdp_sr_bit g2140 (.D(w2174), .nC1(w2144), .nC2(w2146), .C1(w2143), .C2(w2145), .Q(w2176) );
	vdp_sr_bit g2141 (.D(w2149), .nC1(w2144), .nC2(w2146), .C1(w2143), .C2(w2145), .Q(w2148) );
	vdp_not g2142 (.nZ(w2175), .A(w2176) );
	vdp_and g2143 (.Z(w2147), .A(w2174), .B(w2175) );
	vdp_nor g2144 (.Z(w2149), .A(w2148), .B(w2147) );
	vdp_cnt_bit g2145 (.CI(w2148), .R(w2147), .C1(w2143), .nC1(w2144), .nC2(w2146), .C2(w2145), .Q(w2173) );
	vdp_dlatch_inv g2146 (.nQ(w2172), .D(w2173), .nC(w2144), .C(w2143) );
	vdp_not g2147 (.nZ(w2171), .A(w2172) );
	vdp_nand g2148 (.Z(w2170), .A(w2148), .B(w2172) );
	vdp_not g2149 (.nZ(w2169), .A(w2170) );
	vdp_not g2150 (.nZ(w2168), .A(w2167) );
	vdp_not g2151 (.nZ(PSG_CLK1), .A(w2170) );
	vdp_not g2152 (.nZ(PSG_nCLK1), .A(w2169) );
	vdp_not g2153 (.nZ(PSG_nCLK2), .A(w2168) );
	vdp_not g2154 (.nZ(PSG_CLK2), .A(w2167) );
	vdp_nand g2155 (.Z(w2167), .A(w2148), .B(w2171) );
	vdp_sr_bit g2156 (.D(w2277), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2133) );
	vdp_sr_bit g2157 (.D(w2278), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2277) );
	vdp_sr_bit g2158 (.D(w2276), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2278) );
	vdp_sr_bit g2159 (.D(w2137), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2276) );
	vdp_sr_bit g2160 (.D(w2275), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2136) );
	vdp_sr_bit g2161 (.D(w2274), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2275) );
	vdp_sr_bit g2162 (.D(w2273), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2274) );
	vdp_sr_bit g2163 (.D(w2141), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2273) );
	vdp_sr_bit g2164 (.D(w2272), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2140) );
	vdp_sr_bit g2165 (.D(w2271), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2272) );
	vdp_sr_bit g2166 (.D(w2270), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2271) );
	vdp_sr_bit g2167 (.D(w2203), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2270) );
	vdp_sr_bit g2168 (.D(w2268), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2202) );
	vdp_sr_bit g2169 (.D(w2269), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2268) );
	vdp_sr_bit g2170 (.D(w2267), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2269) );
	vdp_sr_bit g2171 (.D(w2201), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2267) );
	vdp_sr_bit g2172 (.D(w2266), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2200) );
	vdp_sr_bit g2173 (.D(w2265), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2266) );
	vdp_sr_bit g2174 (.D(w2264), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2265) );
	vdp_sr_bit g2175 (.D(w2189), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2264) );
	vdp_sr_bit g2176 (.D(w2263), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2188) );
	vdp_sr_bit g2177 (.D(w2262), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2263) );
	vdp_sr_bit g2178 (.D(w2259), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2262) );
	vdp_sr_bit g2179 (.D(w2186), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2259) );
	vdp_sr_bit g2180 (.D(w2260), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2187) );
	vdp_sr_bit g2181 (.D(w2261), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2260) );
	vdp_sr_bit g2182 (.D(w2287), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2261) );
	vdp_sr_bit g2183 (.D(w2255), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2287) );
	vdp_sr_bit g2184 (.D(w2286), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2256) );
	vdp_sr_bit g2185 (.D(w2288), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2286) );
	vdp_sr_bit g2186 (.D(w2289), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2288) );
	vdp_sr_bit g2187 (.D(w2224), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2289) );
	vdp_sr_bit g2188 (.D(w2214), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2223) );
	vdp_sr_bit g2189 (.D(w2215), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2214) );
	vdp_sr_bit g2190 (.D(w2216), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2215) );
	vdp_sr_bit g2191 (.D(w2225), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2216) );
	vdp_sr_bit g2192 (.D(w2131), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2221) );
	vdp_sr_bit g2193 (.D(w2130), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2131) );
	vdp_sr_bit g2194 (.D(w2129), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2130) );
	vdp_sr_bit g2195 (.D(w2127), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2129) );
	vdp_aon2222 g2196 (.Z(w1999), .D2(1'b0), .C2(w2003), .C1(w1995), .D1(w2002), .B1(w1992), .A2(w1991), .A1(w1993), .B2(w2001) );
	vdp_cgi2a g2197 (.Z(w2341), .A(w1999), .C(w2353), .B(w2133) );
	vdp_aon2222 g2198 (.Z(w2000), .D2(1'b0), .C2(w1994), .C1(w1995), .D1(w2002), .B1(w1996), .A2(w1997), .A1(w1993), .B2(w2001) );
	vdp_cgi2a g2199 (.Z(w2353), .A(w2000), .C(w2352), .B(w2136) );
	vdp_aon2222 g2200 (.Z(w2247), .D2(1'b0), .C2(w2242), .C1(w1995), .D1(w2002), .B1(w2244), .A2(w2243), .A1(w1993), .B2(w2001) );
	vdp_cgi2a g2201 (.Z(w2352), .A(w2247), .C(w2351), .B(w2140) );
	vdp_aon2222 g2202 (.Z(w2246), .D2(w2324), .C2(w2347), .C1(w1995), .D1(w2002), .B1(w2348), .A2(w2349), .A1(w1993), .B2(w2001) );
	vdp_cgi2a g2203 (.Z(w2351), .A(w2246), .C(w2253), .B(w2202) );
	vdp_aon2222 g2204 (.Z(w2245), .D2(w2306), .C2(w2307), .C1(w1995), .D1(w2002), .B1(w2309), .A2(w2308), .A1(w1993), .B2(w2001) );
	vdp_cgi2a g2205 (.Z(w2253), .A(w2245), .C(w2254), .B(w2200) );
	vdp_aon2222 g2206 (.Z(w2317), .D2(w2252), .C2(w2344), .C1(w1995), .D1(w2002), .B1(w2345), .A2(w2346), .A1(w1993), .B2(w2001) );
	vdp_cgi2a g2207 (.Z(w2254), .A(w2317), .C(w2350), .B(w2188) );
	vdp_aon2222 g2208 (.Z(w2316), .D2(1'b0), .C2(w2310), .C1(w1995), .D1(w2002), .B1(w2311), .A2(w2312), .A1(w1993), .B2(w2001) );
	vdp_cgi2a g2209 (.Z(w2350), .A(w2316), .C(w2343), .B(w2187) );
	vdp_aon2222 g2210 (.Z(w2318), .D2(1'b0), .C2(w2313), .C1(w1995), .D1(w2002), .B1(w2314), .A2(w2315), .A1(w1993), .B2(w2001) );
	vdp_cgi2a g2211 (.Z(w2343), .A(w2318), .C(w2217), .B(w2256) );
	vdp_aon2222 g2212 (.Z(w2319), .D2(1'b0), .C2(w2325), .C1(w1995), .D1(w2002), .B1(w2326), .A2(w2327), .A1(w1993), .B2(w2001) );
	vdp_cgi2a g2213 (.Z(w2217), .A(w2319), .C(w2218), .B(w2223) );
	vdp_aon2222 g2214 (.Z(w2220), .D2(1'b0), .C2(w2323), .C1(w1995), .D1(w2002), .B1(w2321), .A2(w2322), .A1(w1993), .B2(w2001) );
	vdp_cgi2a g2215 (.Z(w2218), .A(w2220), .C(1'b1), .B(w2221) );
	vdp_not g2216 (.nZ(w2002), .A(w2320) );
	vdp_sr_bit g2217 (.D(w2301), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .Q(w2222) );
	vdp_nand g2218 (.Z(w2320), .A(w2296), .B(w2222) );
	vdp_not g2219 (.nZ(w1995), .A(w2302) );
	vdp_sr_bit g2220 (.D(w2297), .Q(w2301), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_nand g2221 (.Z(w2302), .A(w2296), .B(w2301) );
	vdp_not g2222 (.nZ(w2001), .A(w2300) );
	vdp_sr_bit g2223 (.D(w2233), .Q(w2297), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_nand g2224 (.Z(w2300), .A(w2296), .B(w2297) );
	vdp_not g2225 (.nZ(w1993), .A(w2298) );
	vdp_sr_bit g2226 (.D(w2299), .Q(w2233), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_nand g2227 (.Z(w2298), .A(w2296), .B(w2233) );
	vdp_sr_bit g2228 (.D(w2123), .Q(w2204), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_sr_bit g2229 (.D(w2305), .Q(w2303), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_sr_bit g2230 (.D(w2304), .Q(w2305), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_sr_bit g2231 (.D(w2232), .Q(w2304), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_sr_bit g2232 (.D(w2341), .Q(w2232), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2) );
	vdp_not g2233 (.nZ(w2296), .A(w2204) );
	vdp_nor4 g2234 (.Z(w2299), .A(w2301), .B(w2297), .D(w2233), .C(w2123) );
	vdp_nor4 g2235 (.Z(w2194), .A(w2236), .B(w2237), .D(w2234), .C(w2235) );
	vdp_nor4 g2236 (.Z(w2196), .A(w2229), .B(w2230), .D(w2209), .C(w2210) );
	vdp_nor3 g2237 (.Z(w2195), .A(w2205), .B(w2206), .C(w2207) );
	vdp_not g2238 (.nZ(w1981), .A(w2204) );
	vdp_nand4 g2239 (.Z(w2193), .A(w2194), .B(w2196), .D(w2164), .C(w2195) );
	vdp_nand g2240 (.Z(w2198), .A(w2132), .B(w2197) );
	vdp_nand g2241 (.Z(w2199), .A(w2193), .B(w2198) );
	vdp_lfsr_bit g2242 (.Q(w2229), .A(w2199), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2227), .B(w2228) );
	vdp_lfsr_bit g2243 (.Q(w2230), .A(w2229), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2227), .B(w2228) );
	vdp_lfsr_bit g2244 (.Q(w2210), .A(w2230), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2227), .B(w2228) );
	vdp_lfsr_bit g2245 (.Q(w2209), .A(w2210), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2227), .B(w2228) );
	vdp_lfsr_bit g2246 (.Q(w2205), .A(w2209), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2227), .B(w2228) );
	vdp_lfsr_bit g2247 (.Q(w2206), .A(w2205), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2227), .B(w2228) );
	vdp_lfsr_bit g2248 (.Q(w2207), .A(w2206), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2227), .B(w2228) );
	vdp_lfsr_bit g2249 (.Q(w2234), .A(w2207), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2227), .B(w2228) );
	vdp_lfsr_bit g2250 (.Q(w2235), .A(w2234), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2227), .B(w2228) );
	vdp_lfsr_bit g2251 (.Q(w2236), .A(w2235), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2227), .B(w2228) );
	vdp_lfsr_bit g2252 (.Q(w2237), .A(w2236), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2227), .B(w2228) );
	vdp_lfsr_bit g2253 (.Q(w2238), .A(w2237), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2227), .B(w2228) );
	vdp_lfsr_bit g2254 (.Q(w2239), .A(w2238), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2227), .B(w2228) );
	vdp_lfsr_bit g2255 (.Q(w2226), .A(w2239), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2227), .B(w2228) );
	vdp_lfsr_bit g2256 (.Q(w2126), .A(w2226), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2227), .B(w2228) );
	vdp_lfsr_bit g2257 (.Q(w2240), .A(w2126), .C2(PSG_CLK2), .C1(PSG_CLK1), .nC2(PSG_nCLK2), .nC1(PSG_nCLK1), .C(w2227), .B(w2228) );
	vdp_xor g2258 (.Z(w2132), .A(w2239), .B(w2240) );
	vdp_and g2259 (.Z(w2285), .A(w2128), .B(w2221) );
	vdp_ha g2260 (.SUM(w2127), .CO(w2183), .B(w2285), .A(1'b1) );
	vdp_and g2261 (.Z(w2258), .A(w2128), .B(w2223) );
	vdp_ha g2262 (.SUM(w2225), .CO(w2182), .B(w2258), .A(w2183) );
	vdp_and g2263 (.Z(w2257), .A(w2128), .B(w2256) );
	vdp_ha g2264 (.SUM(w2224), .CO(w2181), .B(w2257), .A(w2182) );
	vdp_and g2265 (.Z(w2185), .A(w2128), .B(w2187) );
	vdp_ha g2266 (.SUM(w2255), .CO(w2180), .B(w2185), .A(w2181) );
	vdp_and g2267 (.Z(w2284), .A(w2128), .B(w2188) );
	vdp_ha g2268 (.SUM(w2186), .CO(w2179), .B(w2284), .A(w2180) );
	vdp_and g2269 (.Z(w2283), .A(w2128), .B(w2200) );
	vdp_ha g2270 (.SUM(w2189), .CO(w2178), .B(w2283), .A(w2179) );
	vdp_and g2271 (.Z(w2282), .A(w2128), .B(w2202) );
	vdp_ha g2272 (.SUM(w2201), .CO(w2177), .B(w2282), .A(w2178) );
	vdp_and g2273 (.Z(w2281), .A(w2128), .B(w2140) );
	vdp_ha g2274 (.SUM(w2203), .CO(w2139), .B(w2281), .A(w2177) );
	vdp_and g2275 (.Z(w2280), .A(w2128), .B(w2136) );
	vdp_ha g2276 (.SUM(w2141), .CO(w2138), .B(w2280), .A(w2139) );
	vdp_and g2277 (.Z(w2279), .A(w2128), .B(w2133) );
	vdp_ha g2278 (.SUM(w2137), .B(w2279), .A(w2138) );
	vdp_and g2279 (.Z(w2208), .A(w2233), .B(w2303) );
	vdp_cnt_bit g2280 (.CI(w2208), .R(w2204), .C1(PSG_CLK1), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C2(PSG_CLK2), .Q(w2334) );
	vdp_and g2281 (.Z(w2212), .A(w2233), .B(w2305) );
	vdp_cnt_bit g2282 (.CI(w2212), .R(w2204), .C1(PSG_CLK1), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C2(PSG_CLK2), .Q(w2335) );
	vdp_and g2283 (.Z(w2211), .A(w2233), .B(w2304) );
	vdp_cnt_bit g2284 (.CI(w2211), .R(w2204), .C1(PSG_CLK1), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C2(PSG_CLK2), .Q(w2158) );
	vdp_and g2285 (.Z(w2231), .A(w2233), .B(w2232) );
	vdp_cnt_bit g2286 (.CI(w2231), .R(w2204), .C1(PSG_CLK1), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C2(PSG_CLK2), .Q(w2151) );
	vdp_nor g2287 (.Z(w2128), .A(w2341), .B(w2204) );
	vdp_slatch g2288 (.Q(w1982), .C(w1979), .D(DB[7]), .nC(w1980) );
	vdp_comp_str g2289 (.A(nPSGWRITE), .Z(w1979), .nZ(w1980) );
	vdp_and g2290 (.Z(w1974), .A(w1981), .B(w1982) );
	vdp_and g2291 (.Z(w1976), .A(w1975), .B(w1974) );
	vdp_and g2292 (.Z(w2360), .A(w1981), .B(w2359) );
	vdp_slatch g2293 (.Q(w2359), .C(w1979), .D(DB[6]), .nC(w1980) );
	vdp_slatch g2294 (.Q(w2102), .C(w1977), .D(w2360), .nC(w1978) );
	vdp_and g2295 (.Z(w1983), .A(w1981), .B(w2070) );
	vdp_slatch g2296 (.Q(w2070), .C(w1979), .D(DB[5]), .nC(w1980) );
	vdp_slatch g2297 (.Q(w2071), .C(w1977), .D(w1983), .nC(w1978) );
	vdp_and g2298 (.Z(w1986), .A(w1981), .B(w2069) );
	vdp_slatch g2299 (.Q(w2069), .C(w1979), .D(DB[4]), .nC(w1980) );
	vdp_slatch g2300 (.Q(w2101), .C(w1977), .D(w1986), .nC(w1978) );
	vdp_and g2301 (.Z(w2251), .A(w1981), .B(w2108) );
	vdp_slatch g2302 (.Q(w2108), .C(w1979), .D(DB[3]), .nC(w1980) );
	vdp_or g2303 (.Z(w2094), .A(w2109), .B(w2251) );
	vdp_and g2304 (.Z(w2249), .A(w1981), .B(w2358) );
	vdp_or g2305 (.Z(w2082), .A(w2109), .B(w2249) );
	vdp_slatch g2306 (.Q(w2358), .C(w1979), .D(DB[2]), .nC(w1980) );
	vdp_not g2307 (.nZ(w2109), .A(w1981) );
	vdp_and g2308 (.Z(w2248), .A(w1981), .B(w2250) );
	vdp_or g2309 (.Z(w2080), .A(w2109), .B(w2248) );
	vdp_slatch g2310 (.Q(w2250), .C(w1979), .D(DB[1]), .nC(w1980) );
	vdp_and g2311 (.Z(w2114), .A(w1981), .B(w2115) );
	vdp_or g2312 (.Z(w2083), .A(w2109), .B(w2114) );
	vdp_slatch g2313 (.Q(w2115), .C(w1979), .D(DB[0]), .nC(w1980) );
	vdp_not g2314 (.nZ(w2113), .A(w2111) );
	vdp_aoi21 g2315 (.Z(w2111), .B(w2123), .A1(w2116), .A2(w2110) );
	vdp_and3 g2316 (.Z(w2110), .A(w2091), .B(w2090), .C(w2101) );
	vdp_not g2317 (.nZ(w2112), .A(w2356) );
	vdp_aoi21 g2318 (.Z(w2356), .B(w2123), .A1(w2116), .A2(w2357) );
	vdp_and3 g2319 (.Z(w2357), .A(w2091), .B(w2071), .C(w2101) );
	vdp_not g2320 (.nZ(w2366), .A(w2355) );
	vdp_aoi21 g2321 (.Z(w2355), .B(w2123), .A1(w2116), .A2(w2354) );
	vdp_and3 g2322 (.Z(w2354), .A(w2102), .B(w2090), .C(w2092) );
	vdp_not g2323 (.nZ(w2120), .A(w1974) );
	vdp_or g2324 (.Z(w2122), .A(w1974), .B(w2123) );
	vdp_and g2325 (.Z(w2361), .A(w2122), .B(w2366) );
	vdp_and g2326 (.Z(w2241), .A(w2120), .B(w2366) );
	vdp_and g2327 (.Z(w2332), .A(w2122), .B(w2107) );
	vdp_and g2328 (.Z(w2362), .A(w2120), .B(w2107) );
	vdp_not g2329 (.nZ(w2107), .A(w2106) );
	vdp_aoi21 g2330 (.Z(w2106), .B(w2123), .A1(w2116), .A2(w2105) );
	vdp_and3 g2331 (.Z(w2105), .A(w2091), .B(w2071), .C(w2092) );
	vdp_not g2332 (.nZ(w2103), .A(w2104) );
	vdp_aoi21 g2333 (.Z(w2104), .B(w2123), .A1(w2116), .A2(w2118) );
	vdp_and3 g2334 (.Z(w2118), .A(w2102), .B(w2090), .C(w2101) );
	vdp_and g2335 (.Z(w2121), .A(w2122), .B(w2117) );
	vdp_and g2336 (.Z(w2119), .A(w2120), .B(w2117) );
	vdp_not g2337 (.nZ(w2117), .A(w2100) );
	vdp_aoi21 g2338 (.Z(w2100), .B(w2123), .A1(w2116), .A2(w2099) );
	vdp_and3 g2339 (.Z(w2099), .A(w2091), .B(w2090), .C(w2092) );
	vdp_and3 g2340 (.Z(w2098), .A(w2102), .B(w2071), .C(w2101) );
	vdp_not g2341 (.nZ(w2086), .A(w2097) );
	vdp_aoi21 g2342 (.Z(w2097), .B(w2123), .A1(w2116), .A2(w2098) );
	vdp_and3 g2343 (.Z(w2095), .A(w2102), .B(w2071), .C(w2092) );
	vdp_not g2344 (.nZ(w2150), .A(w2096) );
	vdp_aoi21 g2345 (.Z(w2096), .B(w2123), .A1(w2116), .A2(w2095) );
	vdp_not g2346 (.nZ(w2337), .A(w2340) );
	vdp_not g2347 (.nZ(w2338), .A(w2339) );
	vdp_not g2348 (.nZ(w2092), .A(w2101) );
	vdp_not g2349 (.nZ(w2090), .A(w2071) );
	vdp_not g2350 (.nZ(w2091), .A(w2102) );
	vdp_nor g2351 (.Z(w1966), .A(w2334), .B(PSG_TEST9) );
	vdp_nor g2352 (.Z(w2068), .A(w2335), .B(PSG_TEST9) );
	vdp_nor g2353 (.Z(w2081), .A(w2158), .B(PSG_TEST9) );
	vdp_nor g2354 (.Z(w2088), .A(w2126), .B(PSG_TEST9) );
	vdp_aon22 g2355 (.Z(w2153), .A2(w2158), .A1(w2157), .B2(w2152), .B1(w2151) );
	vdp_sr_bit g2356 (.D(w2153), .nC1(PSG_nCLK1), .nC2(PSG_nCLK2), .C1(PSG_CLK1), .C2(PSG_CLK2), .Q(w2154) );
	vdp_not g2357 (.nZ(w2152), .A(w2157) );
	vdp_not g2358 (.nZ(w2155), .A(w2154) );
	vdp_not g2359 (.nZ(w2291), .A(PSG_TEST10) );
	vdp_not g2360 (.nZ(w2290), .A(PSG_TEST11) );
	vdp_not g2361 (.nZ(w2191), .A(w2190) );
	vdp_sr_bit g2362 (.D(w1975), .nC1(w2144), .nC2(w2146), .C1(w2143), .C2(w2145), .Q(w2116) );
	vdp_nand g2363 (.Z(w2292), .A(PSG_TEST10), .B(w2290) );
	vdp_nand g2364 (.Z(w2156), .A(PSG_TEST11), .B(PSG_TEST10) );
	vdp_nand g2365 (.Z(w2293), .A(w2290), .B(w2291) );
	vdp_nand g2366 (.Z(w2294), .A(PSG_TEST11), .B(w2291) );
	vdp_and g2367 (.Z(w2160), .A(w2153), .B(w2155) );
	vdp_and g2368 (.Z(w1940), .A(PSG_TEST9), .B(w2156) );
	vdp_and g2369 (.Z(w1942), .A(PSG_TEST9), .B(w2292) );
	vdp_and g2370 (.Z(w1941), .A(PSG_TEST9), .B(w2293) );
	vdp_and g2371 (.Z(w1939), .A(PSG_TEST9), .B(w2294) );
	vdp_nor4 g2372 (.Z(w2164), .A(w2226), .B(w2239), .D(w2238), .C(w2126) );
	vdp_not g2373 (.nZ(w2161), .A(w2160) );
	vdp_not g2374 (.nZ(w2228), .A(w2162) );
	vdp_not g2375 (.nZ(w2227), .A(w2295) );
	vdp_not g2376 (.nZ(w2123), .A(w2191) );
	vdp_nand g2377 (.Z(w2162), .A(w2159), .B(w2161) );
	vdp_nand g2378 (.Z(w2295), .A(w2159), .B(w2160) );
	vdp_nor g2379 (.Z(w2159), .A(w2123), .B(w2163) );
	vdp_rs_ff g2380 (.S(w2150), .R(w2163), .Q(w2192) );
	vdp_rs_ff g2381 (.S(w1975), .R(nPSGWRITE), .Q(w2165) );
	vdp_nor g2382 (.Z(w2166), .A(nPSGWRITE), .B(w2165) );
	vdp_comp_dff g2383 (.D(w2166), .nC1(w2144), .C1(w2143), .C2(w2145), .nC2(w2146), .Q(w1975) );
	vdp_comp_dff g2384 (.D(SYSRES), .nC1(PSG_nCLK1), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC2(PSG_nCLK2), .Q(w2190) );
	vdp_comp_dff g2385 (.D(w2192), .nC1(PSG_nCLK1), .C1(PSG_CLK1), .C2(PSG_CLK2), .nC2(PSG_nCLK2), .Q(w2163) );
	vdp_sr_bit g2386 (.Q(w2534), .D(w2528), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2387 (.nZ(AD_RD_DIR), .A(w2527) );
	vdp_sr_bit g2388 (.Q(w2535), .D(w2398), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2389 (.Q(w2463), .D(w2411), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2390 (.Q(w2518), .D(w760), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2391 (.Q(w2390), .D(w517), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2392 (.nZ(w2530), .A(w2388) );
	vdp_or g2393 (.Z(w2398), .A(w517), .B(w2390) );
	vdp_sr_bit g2394 (.Q(w2407), .D(w2409), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_sr_bit g2395 (.Q(w2531), .D(w2520), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2396 (.nZ(w2462), .A(w2531) );
	vdp_or g2397 (.Z(w2386), .A(w2390), .B(w2389) );
	vdp_sr_bit g2398 (.Q(w2389), .D(w518), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2399 (.Q(w2387), .D(w30), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2400 (.Q(w2522), .D(w2387), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2401 (.Q(w2521), .D(w2399), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2402 (.Q(w2516), .D(w2518), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2403 (.Q(w2533), .D(w2538), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_not g2404 (.nZ(w2512), .A(w2578) );
	vdp_not g2405 (.nZ(w2410), .A(VRAM128k) );
	vdp_sr_bit g2406 (.Q(w2399), .D(VRAM_REFRESH), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2407 (.nZ(w2470), .A(w2385) );
	vdp_not g2408 (.nZ(w2536), .A(w2523) );
	vdp_not g2409 (.nZ(w2405), .A(w2397) );
	vdp_oai21 g2410 (.Z(w2385), .B(w2405), .A1(w2536), .A2(w2524) );
	vdp_or g2411 (.Z(w2397), .A(w2530), .B(w2529) );
	vdp_or g2412 (.Z(w2528), .A(w2389), .B(w518) );
	vdp_not g2413 (.nZ(w2537), .A(w2391) );
	vdp_not g2414 (.nZ(w2570), .A(w2538) );
	vdp_dlatch_inv g2415 (.nQ(w2538), .D(w3), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2416 (.nQ(w2532), .D(w2406), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g2417 (.nQ(w2406), .D(w2533), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g2418 (.nQ(w2388), .D(w2386), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2419 (.nQ(w2529), .D(w2388), .C(HCLK2), .nC(nHCLK2) );
	vdp_dlatch_inv g2420 (.nQ(w2526), .D(w2525), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2421 (.nQ(w2523), .D(w2522), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2422 (.nQ(w2524), .D(w2523), .C(HCLK2), .nC(nHCLK2) );
	vdp_aon22 g2423 (.Z(nCAS1), .A1(w2406), .B1(w2395), .B2(1'b1), .A2(w2531) );
	vdp_and3 g2424 (.Z(nWE1), .A(w2394), .B(w2535), .C(w2395) );
	vdp_and3 g2425 (.Z(nWE0), .A(w2395), .B(w2394), .C(w2534) );
	vdp_aoi222 g2426 (.Z(w2527), .A1(1'b1), .B1(w2392), .B2(1'b1), .A2(w85), .C1(w2397), .C2(w2395) );
	vdp_aon333 g2427 (.Z(nOE1), .A1(w2470), .A2(w2533), .A3(w2395), .B1(w2526), .B2(w2526), .B3(w2537), .C1(w2526), .C2(w2526), .C3(w2392) );
	vdp_or3 g2428 (.Z(w2525), .A(w2520), .B(w2522), .C(w2387) );
	vdp_sr_bit g2429 (.Q(w2392), .D(w2570), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_dlatch_inv g2430 (.nQ(w2394), .D(w2392), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g2431 (.nQ(w2519), .D(w2394), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g2432 (.nQ(w2395), .D(w2393), .C(DCLK1), .nC(nDCLK1) );
	vdp_not g2433 (.nZ(w2393), .A(w2519) );
	vdp_nand g2434 (.Z(w2604), .A(w2519), .B(w2392) );
	vdp_nand g2435 (.Z(w2603), .A(w2392), .B(w2532) );
	vdp_nand g2436 (.Z(w2401), .A(w2533), .B(1'b1) );
	vdp_aoi33 g2437 (.Z(w2584), .A1(w2516), .A2(w561), .A3(w561), .B1(w2412), .B2(w2413), .B3(w3) );
	vdp_and g2438 (.Z(w2408), .A(w2395), .B(w2394) );
	vdp_not g2439 (.nZ(w2402), .A(w2463) );
	vdp_comp_strong g2440 (.nZ(w2419), .Z(w2418), .A(w2425) );
	vdp_comp_strong g2441 (.nZ(w2485), .Z(w2507), .A(w2508) );
	vdp_comp_strong g2442 (.nZ(w2420), .Z(w2464), .A(w2508) );
	vdp_comp_strong g2443 (.nZ(w2468), .Z(w2467), .A(w2425) );
	vdp_comp_strong g2444 (.nZ(w2426), .Z(w2469), .A(w2422) );
	vdp_comp_strong g2445 (.nZ(w2472), .Z(w2513), .A(w2422) );
	vdp_not g2446 (.nZ(w2428), .A(w2392) );
	vdp_not g2447 (.nZ(w2413), .A(w561) );
	vdp_not g2448 (.nZ(w2412), .A(w31) );
	vdp_comp_strong g2449 (.nZ(w2466), .Z(w6533), .A(w2408) );
	vdp_comp_strong g2450 (.nZ(w2403), .Z(w2509), .A(w2408) );
	vdp_or g2451 (.Z(w2520), .A(w2399), .B(w2521) );
	vdp_and g2452 (.Z(w2409), .A(VRAM128k), .B(HCLK1) );
	vdp_comp_we g2453 (.nZ(w2510), .Z(w2511), .A(w85) );
	vdp_comp_we g2454 (.nZ(w2421), .Z(w2582), .A(w2429) );
	vdp_not g2455 (.nZ(w2583), .A(w2463) );
	vdp_not g2456 (.nZ(w2424), .A(w2604) );
	vdp_not g2457 (.nZ(w6538), .A(w2603) );
	vdp_not g2458 (.nZ(w6539), .A(w2401) );
	vdp_comp_we g2459 (.nZ(w6540), .Z(w2515), .A(M5) );
	vdp_comp_we g2460 (.nZ(w2471), .Z(w2427), .A(VRAM128k) );
	vdp_and g2461 (.Z(w2411), .A(w95), .B(w3) );
	vdp_and g2462 (.Z(w2422), .A(w3), .B(HCLK1) );
	vdp_and g2463 (.Z(w2425), .A(HCLK2), .B(w2517) );
	vdp_and g2464 (.Z(w2508), .A(w3), .B(HCLK1) );
	vdp_oai21 g2465 (.Z(w2578), .A1(HCLK2), .A2(w2410), .B(DCLK1) );
	vdp_notif0 g2466 (.nZ(AD_DATA[0]), .A(w2416), .nE(w2402) );
	vdp_aon22 g2467 (.Z(nYS), .A1(VRAMA[16]), .A2(w2511), .B1(w2510), .B2(w2567) );
	vdp_aon22 g2468 (.Z(w2552), .A1(VRAMA[15]), .B1(w2510), .A2(w2511), .B2(w2491) );
	vdp_aon22 g2469 (.Z(w2550), .A1(VRAMA[14]), .B1(w2510), .A2(w2511), .B2(w2377) );
	vdp_aon22 g2470 (.Z(w2600), .A1(VRAMA[6]), .B1(w2510), .A2(w2511), .B2(w2551) );
	vdp_aon22 g2471 (.Z(w2490), .A1(VRAMA[7]), .B1(w2510), .A2(w2511), .B2(w2369) );
	vdp_aon22 g2472 (.Z(w2568), .A1(VRAMA[13]), .B1(w2510), .A2(w2511), .B2(w2384) );
	vdp_aon22 g2473 (.Z(w2589), .A1(VRAMA[5]), .B1(w2510), .A2(w2511), .B2(w2586) );
	vdp_aon22 g2474 (.Z(w2554), .A1(VRAMA[12]), .B1(w2510), .A2(w2511), .B2(w2452) );
	vdp_aon22 g2475 (.Z(w2602), .A1(VRAMA[4]), .B1(w2510), .A2(w2511), .B2(w2459) );
	vdp_aon22 g2476 (.Z(w2553), .A1(VRAMA[11]), .B1(w2510), .A2(w2511), .B2(w2593) );
	vdp_aon22 g2477 (.Z(w2594), .A1(VRAMA[3]), .B1(w2510), .A2(w2511), .B2(w2587) );
	vdp_aon22 g2478 (.Z(w2569), .A1(VRAMA[10]), .B1(w2510), .A2(w2511), .B2(w2503) );
	vdp_aon22 g2479 (.Z(w2592), .A1(VRAMA[2]), .B1(w2510), .A2(w2511), .B2(w2448) );
	vdp_aon22 g2480 (.Z(w2414), .A1(VRAMA[8]), .B1(w2510), .A2(w2511), .B2(w2417) );
	vdp_aon22 g2481 (.Z(w2590), .A1(VRAMA[0]), .B1(w2510), .A2(w2511), .B2(w2440) );
	vdp_aon22 g2482 (.Z(w2591), .A1(VRAMA[9]), .B1(w2510), .A2(w2511), .B2(w2486) );
	vdp_aon22 g2483 (.Z(w2601), .A1(VRAMA[1]), .B1(w2510), .A2(w2511), .B2(w2444) );
	vdp_notif0 g2484 (.nZ(AD_DATA[1]), .A(w2435), .nE(w2402) );
	vdp_notif0 g2485 (.nZ(AD_DATA[2]), .A(w2488), .nE(w2402) );
	vdp_notif0 g2486 (.nZ(AD_DATA[3]), .A(w2445), .nE(w2402) );
	vdp_notif0 g2487 (.nZ(AD_DATA[5]), .A(w2383), .nE(w2402) );
	vdp_notif0 g2488 (.nZ(AD_DATA[4]), .A(w2465), .nE(w2402) );
	vdp_notif0 g2489 (.nZ(AD_DATA[6]), .A(w2378), .nE(w2402) );
	vdp_notif0 g2490 (.nZ(AD_DATA[7]), .A(w2376), .nE(w2402) );
	vdp_slatch g2491 (.nQ(w2416), .D(w2415), .nC(w2403), .C(w2509) );
	vdp_slatch g2492 (.nQ(w2435), .D(w2434), .nC(w2403), .C(w2509) );
	vdp_slatch g2493 (.nQ(w2488), .D(w2442), .nC(w2403), .C(w2509) );
	vdp_slatch g2494 (.nQ(w2445), .D(w2446), .nC(w2403), .C(w2509) );
	vdp_slatch g2495 (.nQ(w2465), .D(w2400), .nC(w2403), .C(w2509) );
	vdp_slatch g2496 (.nQ(w2383), .D(w2606), .nC(w2403), .C(w2509) );
	vdp_slatch g2497 (.nQ(w2378), .D(w2454), .nC(w2403), .C(w2509) );
	vdp_slatch g2498 (.nQ(w2376), .D(w2607), .nC(w2403), .C(w2509) );
	vdp_slatch g2499 (.nQ(w2371), .D(w2370), .nC(w2466), .C(w6533) );
	vdp_slatch g2500 (.nQ(w2457), .D(w2453), .nC(w2466), .C(w6533) );
	vdp_slatch g2501 (.nQ(w2494), .D(w2579), .nC(w2466), .C(w6533) );
	vdp_slatch g2502 (.nQ(w2495), .D(w2382), .nC(w2466), .C(w6533) );
	vdp_slatch g2503 (.nQ(w2555), .D(w2455), .nC(w2466), .C(w6533) );
	vdp_slatch g2504 (.nQ(w2449), .D(w2447), .nC(w2466), .C(w6533) );
	vdp_slatch g2505 (.nQ(w2443), .D(w2489), .nC(w2466), .C(w6533) );
	vdp_slatch g2506 (.nQ(w2473), .D(w2612), .nC(w2466), .C(w6533) );
	vdp_slatch g2507 (.Q(w2417), .D(w2476), .nC(w2419), .C(w2418) );
	vdp_slatch g2508 (.Q(w2486), .D(w2596), .nC(w2419), .C(w2418) );
	vdp_slatch g2509 (.Q(w2593), .D(w2558), .nC(w2419), .C(w2418) );
	vdp_slatch g2510 (.Q(w2503), .D(w2487), .nC(w2419), .C(w2418) );
	vdp_slatch g2511 (.Q(w2384), .D(w2475), .nC(w2419), .C(w2418) );
	vdp_slatch g2512 (.Q(w2452), .D(w2559), .nC(w2419), .C(w2418) );
	vdp_slatch g2513 (.Q(w2491), .D(w2562), .nC(w2419), .C(w2418) );
	vdp_slatch g2514 (.Q(w2377), .D(w2474), .nC(w2419), .C(w2418) );
	vdp_slatch g2515 (.nQ(w2561), .D(w334), .nC(w2485), .C(w2507) );
	vdp_slatch g2516 (.nQ(w2563), .D(RD_DATA[6]), .nC(w2485), .C(w2507) );
	vdp_slatch g2517 (.nQ(w2560), .D(RD_DATA[5]), .nC(w2485), .C(w2507) );
	vdp_slatch g2518 (.nQ(w2598), .D(RD_DATA[4]), .nC(w2485), .C(w2507) );
	vdp_slatch g2519 (.nQ(w2557), .D(w300), .nC(w2485), .C(w2507) );
	vdp_slatch g2520 (.nQ(w2599), .D(RD_DATA[2]), .nC(w2485), .C(w2507) );
	vdp_slatch g2521 (.nQ(w2597), .D(RD_DATA[0]), .nC(w2485), .C(w2507) );
	vdp_slatch g2522 (.nQ(w2556), .D(RD_DATA[1]), .nC(w2485), .C(w2507) );
	vdp_notif0 g2523 (.nZ(w334), .A(w2371), .nE(w2583) );
	vdp_notif0 g2524 (.nZ(RD_DATA[6]), .A(w2457), .nE(w2583) );
	vdp_notif0 g2525 (.nZ(RD_DATA[5]), .A(w2494), .nE(w2583) );
	vdp_notif0 g2526 (.nZ(RD_DATA[4]), .A(w2495), .nE(w2583) );
	vdp_notif0 g2527 (.nZ(w300), .A(w2555), .nE(w2583) );
	vdp_notif0 g2528 (.nZ(RD_DATA[2]), .A(w2449), .nE(w2583) );
	vdp_notif0 g2529 (.nZ(RD_DATA[1]), .A(w2443), .nE(w2583) );
	vdp_notif0 g2530 (.nZ(RD_DATA[0]), .A(w2473), .nE(w2583) );
	vdp_slatch g2531 (.nQ(w2572), .D(AD_DATA[7]), .nC(w2420), .C(w2464) );
	vdp_slatch g2532 (.nQ(w2571), .D(AD_DATA[6]), .nC(w2420), .C(w2464) );
	vdp_slatch g2533 (.nQ(w2595), .D(AD_DATA[5]), .nC(w2420), .C(w2464) );
	vdp_slatch g2534 (.nQ(w2574), .D(AD_DATA[3]), .nC(w2420), .C(w2464) );
	vdp_slatch g2535 (.nQ(w2575), .D(AD_DATA[2]), .nC(w2420), .C(w2464) );
	vdp_slatch g2536 (.nQ(w2577), .D(AD_DATA[1]), .nC(w2420), .C(w2464) );
	vdp_slatch g2537 (.nQ(w2576), .D(AD_DATA[0]), .nC(w2420), .C(w2464) );
	vdp_slatch g2538 (.Q(w2375), .D(w2484), .nC(w2468), .C(w2467) );
	vdp_slatch g2539 (.Q(w2381), .D(w2483), .nC(w2468), .C(w2467) );
	vdp_slatch g2540 (.Q(w2456), .D(w2482), .nC(w2468), .C(w2467) );
	vdp_slatch g2541 (.Q(w2580), .D(w2479), .nC(w2468), .C(w2467) );
	vdp_slatch g2542 (.Q(w2506), .D(w2480), .nC(w2468), .C(w2467) );
	vdp_slatch g2543 (.Q(w2441), .D(w2478), .nC(w2468), .C(w2467) );
	vdp_slatch g2544 (.Q(w2493), .D(w2374), .nC(w2426), .C(w2469) );
	vdp_slatch g2545 (.Q(w2585), .D(w2380), .nC(w2426), .C(w2469) );
	vdp_slatch g2546 (.Q(w2565), .D(w2433), .nC(w2426), .C(w2469) );
	vdp_slatch g2547 (.Q(w2497), .D(w2432), .nC(w2426), .C(w2469) );
	vdp_slatch g2548 (.Q(w2504), .D(w2505), .nC(w2426), .C(w2469) );
	vdp_slatch g2549 (.Q(w2581), .D(w2438), .nC(w2426), .C(w2469) );
	vdp_slatch g2550 (.Q(w2502), .D(w2404), .nC(w2426), .C(w2469) );
	vdp_slatch g2551 (.Q(w2588), .D(w2439), .nC(w2426), .C(w2469) );
	vdp_slatch g2552 (.Q(w2514), .D(w2437), .nC(w2472), .C(w2513) );
	vdp_slatch g2553 (.Q(w2501), .D(w2611), .nC(w2472), .C(w2513) );
	vdp_slatch g2554 (.Q(w2450), .D(w2431), .nC(w2472), .C(w2513) );
	vdp_slatch g2555 (.Q(w2498), .D(w2605), .nC(w2472), .C(w2513) );
	vdp_slatch g2556 (.Q(w2460), .D(w2379), .nC(w2472), .C(w2513) );
	vdp_slatch g2557 (.Q(w2496), .D(w2430), .nC(w2472), .C(w2513) );
	vdp_slatch g2558 (.Q(w2458), .D(w2373), .nC(w2472), .C(w2513) );
	vdp_slatch g2559 (.Q(w2492), .D(w2372), .nC(w2472), .C(w2513) );
	vdp_sr_bit g2560 (.Q(w2429), .D(w561), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2561 (.nZ(w2618), .A(w113) );
	vdp_not g2562 (.nZ(w2499), .A(w2500) );
	vdp_not g2563 (.nZ(w6541), .A(M5) );
	vdp_not g2564 (.nZ(w2436), .A(w2428) );
	vdp_not g2565 (.nZ(w2391), .A(w2436) );
	vdp_aoi21 g2566 (.Z(w2500), .B(w2566), .A2(VRAMA[9]), .A1(w6541) );
	vdp_aoi22 g2567 (.Z(w2596), .A1(w2443), .B1(w2421), .B2(w2556), .A2(w2582) );
	vdp_aoi22 g2568 (.Z(w2558), .A1(w2555), .B1(w2421), .B2(w2557), .A2(w2582) );
	vdp_aoi22 g2569 (.Z(w2487), .A1(w2449), .B1(w2421), .B2(w2599), .A2(w2582) );
	vdp_aoi22 g2570 (.Z(w2475), .A1(w2494), .B1(w2421), .B2(w2560), .A2(w2582) );
	vdp_aoi22 g2571 (.Z(w2559), .A1(w2495), .B1(w2421), .B2(w2598), .A2(w2582) );
	vdp_aoi22 g2572 (.Z(w2562), .A1(w2371), .B1(w2421), .B2(w2561), .A2(w2582) );
	vdp_aoi22 g2573 (.Z(w2474), .A1(w2457), .B1(w2421), .B2(w2563), .A2(w2582) );
	vdp_slatch g2574 (.Q(w2423), .D(w2477), .nC(w2468), .C(w2467) );
	vdp_slatch g2575 (.nQ(w2573), .D(AD_DATA[4]), .nC(w2420), .C(w2464) );
	vdp_slatch g2576 (.Q(w2451), .D(w2481), .nC(w2468), .C(w2467) );
	vdp_aoi22 g2577 (.Z(w2477), .A1(w2416), .B1(w2421), .B2(w2576), .A2(w2582) );
	vdp_aoi22 g2578 (.Z(w2478), .A1(w2435), .B1(w2421), .B2(w2577), .A2(w2582) );
	vdp_aoi22 g2579 (.Z(w2479), .A1(w2488), .B1(w2421), .B2(w2575), .A2(w2582) );
	vdp_aoi22 g2580 (.Z(w2480), .A1(w2445), .B1(w2421), .B2(w2574), .A2(w2582) );
	vdp_aoi22 g2581 (.Z(w2481), .A1(w2465), .B1(w2421), .B2(w2573), .A2(w2582) );
	vdp_aoi22 g2582 (.Z(w2482), .A1(w2383), .B1(w2421), .B2(w2595), .A2(w2582) );
	vdp_aoi22 g2583 (.Z(w2484), .A1(w2376), .B1(w2421), .B2(w2572), .A2(w2582) );
	vdp_aoi22 g2584 (.Z(w2483), .A1(w2378), .B1(w2421), .B2(w2571), .A2(w2582) );
	vdp_aon22 g2585 (.Z(w2439), .A1(VRAMA[2]), .B1(w6540), .B2(VRAMA[1]), .A2(w2515) );
	vdp_aon22 g2586 (.Z(w2438), .A1(VRAMA[3]), .B1(w6540), .B2(VRAMA[2]), .A2(w2515) );
	vdp_aon22 g2587 (.Z(w2404), .A1(VRAMA[4]), .B1(w6540), .B2(VRAMA[3]), .A2(w2515) );
	vdp_aon22 g2588 (.Z(w2505), .A1(VRAMA[5]), .B1(w6540), .B2(VRAMA[4]), .A2(w2515) );
	vdp_aon22 g2589 (.Z(w2432), .A1(VRAMA[6]), .B1(w6540), .B2(VRAMA[5]), .A2(w2515) );
	vdp_aon22 g2590 (.Z(w2433), .A1(VRAMA[7]), .B1(w6540), .B2(VRAMA[6]), .A2(w2515) );
	vdp_aon22 g2591 (.Z(w2380), .A1(VRAMA[8]), .B1(w6540), .B2(VRAMA[7]), .A2(w2515) );
	vdp_aon22 g2592 (.Z(w2374), .A1(VRAMA[9]), .B1(w6540), .B2(VRAMA[8]), .A2(w2515) );
	vdp_and g2593 (.Z(w2566), .A(VRAMA[1]), .B(M5) );
	vdp_aon22 g2594 (.Z(w2372), .A1(w2564), .B1(w2471), .B2(VRAMA[15]), .A2(w2427) );
	vdp_aon22 g2595 (.Z(w2373), .A1(VRAMA[15]), .B1(w2471), .B2(VRAMA[14]), .A2(w2427) );
	vdp_aon22 g2596 (.Z(w2379), .A1(VRAMA[14]), .B1(w2471), .B2(VRAMA[13]), .A2(w2427) );
	vdp_aon22 g2597 (.Z(w2605), .A1(VRAMA[12]), .B1(w2471), .B2(VRAMA[11]), .A2(w2427) );
	vdp_aon22 g2598 (.Z(w2430), .A1(VRAMA[13]), .B1(w2471), .B2(VRAMA[12]), .A2(w2427) );
	vdp_aon22 g2599 (.Z(w2431), .A1(VRAMA[11]), .B1(w2471), .B2(VRAMA[10]), .A2(w2427) );
	vdp_aon22 g2600 (.Z(w2611), .A1(VRAMA[10]), .B1(w2471), .B2(w2499), .A2(w2427) );
	vdp_aon22 g2601 (.Z(w2437), .A1(w2566), .B1(w2471), .B2(VRAMA[0]), .A2(w2427) );
	vdp_aon22 g2602 (.Z(w2564), .A1(w2618), .B1(w113), .B2(w79), .A2(VRAMA[16]) );
	vdp_aon222 g2603 (.Z(w2440), .A1(w2424), .A2(w2423), .B1(w6538), .B2(w2588), .C1(w6539), .C2(w2514) );
	vdp_aon222 g2604 (.Z(w2444), .A1(w2424), .A2(w2441), .B1(w6538), .B2(w2581), .C1(w6539), .C2(w2501) );
	vdp_aon222 g2605 (.Z(w2448), .A1(w2424), .A2(w2580), .B1(w6538), .B2(w2502), .C1(w6539), .C2(w2450) );
	vdp_aon222 g2606 (.Z(w2587), .A1(w2424), .A2(w2506), .B1(w6538), .B2(w2504), .C1(w6539), .C2(w2498) );
	vdp_aon222 g2607 (.Z(w2459), .A1(w2424), .A2(w2451), .B1(w6538), .B2(w2497), .C1(w6539), .C2(w2496) );
	vdp_aon222 g2608 (.Z(w2586), .A1(w2424), .A2(w2456), .B1(w6538), .B2(w2565), .C1(w6539), .C2(w2460) );
	vdp_aon222 g2609 (.Z(w2551), .A1(w2424), .A2(w2381), .B1(w6538), .B2(w2585), .C1(w6539), .C2(w2458) );
	vdp_aon222 g2610 (.Z(w2369), .A1(w2424), .A2(w2375), .B1(w6538), .B2(w2493), .C1(w6539), .C2(w2492) );
	vdp_dlatch_inv g2611 (.nQ(w2517), .D(w2584), .C(HCLK1), .nC(nHCLK1) );
	vdp_comp_we g2612 (.Z(w2461), .A(w2519) );
	vdp_aon22 g2613 (.Z(nRAS1), .A1(1'b1), .B1(w2462), .B2(w2406), .A2(w2461) );
	vdp_aoi22 g2614 (.Z(w2476), .A1(w2473), .B1(w2421), .B2(w2597), .A2(w2582) );
	vdp_and g2615 (.Z(w2539), .B(w2617), .A(DCLK2) );
	vdp_nor g2616 (.Z(w2613), .A(w2541), .B(RES) );
	vdp_sr_bit g2617 (.Q(w2541), .D(w2613), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_dlatch_inv g2618 (.nQ(w2614), .D(w2542), .C(DCLK1), .nC(nDCLK1) );
	vdp_and g2619 (.Z(w2615), .A(DCLK2), .B(w2614) );
	vdp_dlatch_inv g2620 (.nQ(w2617), .D(w2541), .C(DCLK1), .nC(nDCLK1) );
	vdp_not g2621 (.nZ(w2545), .A(w2547) );
	vdp_not g2622 (.nZ(w2544), .A(w2616) );
	vdp_neg_dff g2623 (.Q(w2547), .C(DCLK1), .D(1'b1), .R(w2539) );
	vdp_not g2624 (.A(w2541), .nZ(w2542) );
	vdp_neg_dff g2625 (.Q(w2616), .R(w2615), .C(DCLK1), .D(1'b1) );
	vdp_sr_bit g2626 (.Q(w2693), .D(w2685), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2627 (.Q(w2689), .D(w2688), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2628 (.Q(w2877), .D(w2689), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2629 (.Q(w2707), .D(w2877), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2630 (.Q(w2662), .D(RD_DATA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2631 (.Q(w2663), .D(RD_DATA[2]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2632 (.Q(w2664), .D(w300), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2633 (.Q(w2856), .D(w2880), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2634 (.Q(w2880), .D(w2881), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2635 (.Q(w2881), .D(w2882), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2636 (.Q(w2882), .D(w2883), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2637 (.Q(w2883), .D(w2884), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2638 (.Q(w2884), .D(w2885), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2639 (.Q(w2885), .D(w2886), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2640 (.Q(w2886), .D(w17), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2641 (.Q(w2671), .D(w2699), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2642 (.Q(w2669), .D(w2889), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2643 (.Q(w2913), .D(w2891), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2644 (.Q(w2891), .D(w2645), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2645 (.Q(w2645), .D(w93), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2646 (.Q(w2620), .D(w2619), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2647 (.Q(w2625), .D(w2759), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2648 (.Q(w2683), .D(w2871), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2649 (.Q(w2687), .D(w2888), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2650 (.Q(w2703), .D(w2695), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2651 (.Q(w2619), .D(w2698), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2652 (.Q(w2724), .D(w2701), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2653 (.Q(w2723), .D(w2760), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2654 (.Q(PLANE_A_PRIO), .D(w2715), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2655 (.Q(PLANE_B_PRIO), .D(w2716), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2656 (.Q(w2679), .D(w2717), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2657 (.Q(w2722), .D(w2721), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2658 (.Q(w2641), .D(w2720), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2659 (.Q(w2720), .D(COL[7]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2660 (.Q(w2642), .D(w2915), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2661 (.Q(w2915), .D(w114), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2662 (.Q(w2733), .D(w2706), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2663 (.Q(w2719), .D(w2718), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2664 (.Q(SPR_PRIO), .D(w2863), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2665 (.Q(w2730), .D(w1434), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2666 (.Q(w2729), .D(w1435), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2667 (.Q(w2634), .D(w2650), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2668 (.Q(w2639), .D(w2651), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2669 (.Q(w2636), .D(w2661), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2670 (.Q(w2627), .D(w2652), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2671 (.Q(w2646), .D(w2658), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2672 (.Q(w2626), .D(w2653), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2673 (.Q(w2621), .D(w2756), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2674 (.Q(w2631), .D(w2654), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2675 (.Q(w2637), .D(w2648), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_slatch g2676 (.nQ(w2911), .D(w2650), .C(w2647), .nC(w2644) );
	vdp_slatch g2677 (.nQ(w2912), .D(w2648), .C(w2647), .nC(w2644) );
	vdp_slatch g2678 (.nQ(w2910), .D(w2651), .C(w2647), .nC(w2644) );
	vdp_slatch g2679 (.nQ(w2909), .D(w2661), .C(w2647), .nC(w2644) );
	vdp_slatch g2680 (.nQ(w2908), .D(w2652), .C(w2647), .nC(w2644) );
	vdp_slatch g2681 (.nQ(w2907), .D(w2658), .C(w2647), .nC(w2644) );
	vdp_slatch g2682 (.nQ(w2906), .D(w2653), .C(w2647), .nC(w2644) );
	vdp_slatch g2683 (.nQ(w2905), .D(w2756), .C(w2647), .nC(w2644) );
	vdp_slatch g2684 (.nQ(w2904), .D(w2654), .C(w2647), .nC(w2644) );
	vdp_slatch g2685 (.Q(w2705), .D(REG_BUS[7]), .nC(w2682), .C(w2692) );
	vdp_slatch g2686 (.Q(w2702), .D(REG_BUS[5]), .nC(w2682), .C(w2692) );
	vdp_slatch g2687 (.Q(w2694), .D(REG_BUS[4]), .nC(w2682), .C(w2692) );
	vdp_slatch g2688 (.Q(w2690), .D(REG_BUS[3]), .nC(w2682), .C(w2692) );
	vdp_slatch g2689 (.Q(w2686), .D(REG_BUS[2]), .nC(w2682), .C(w2692) );
	vdp_slatch g2690 (.Q(w2876), .D(REG_BUS[1]), .nC(w2682), .C(w2692) );
	vdp_slatch g2691 (.Q(w2684), .D(REG_BUS[0]), .nC(w2682), .C(w2692) );
	vdp_slatch g2692 (.Q(w2849), .D(REG_BUS[6]), .nC(w2682), .C(w2692) );
	vdp_aon2222 g2693 (.Z(w2826), .B2(w2765), .B1(w2770), .A2(w2899), .A1(w2765), .D2(w2761), .D1(w2770), .C2(w2770), .C1(HIGHLIGHT) );
	vdp_aon22 g2694 (.Z(w2791), .B2(w2761), .B1(w2775), .A2(w2900), .A1(w2766) );
	vdp_aon22 g2695 (.Z(w2796), .B2(w2761), .B1(w2771), .A2(w2899), .A1(w2766) );
	vdp_not g2696 (.nZ(w2779), .A(w2825) );
	vdp_not g2697 (.nZ(w2773), .A(w2774) );
	vdp_not g2698 (.nZ(w2778), .A(w2777) );
	vdp_not g2699 (.nZ(w2797), .A(w2826) );
	vdp_not g2700 (.nZ(w2790), .A(w2783) );
	vdp_comp_we g2701 (.Z(w2765), .A(w2669) );
	vdp_not g2702 (.nZ(w2860), .A(w2818) );
	vdp_not g2703 (.nZ(w2821), .A(w2819) );
	vdp_not g2704 (.nZ(w2822), .A(w2823) );
	vdp_not g2705 (.nZ(w2786), .A(HIGHLIGHT) );
	vdp_sr_bit g2706 (.Q(SHADOW), .D(w2642), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2707 (.Q(w2823), .D(w2640), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2708 (.Q(HIGHLIGHT), .D(w2641), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2709 (.Q(w2818), .D(w2820), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2710 (.Q(w2819), .D(w2665), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g2711 (.Z(w2895), .A(w2822), .B(w2860), .C(w2819) );
	vdp_and3 g2712 (.Z(w2897), .A(w2821), .B(w2823), .C(w2860) );
	vdp_and3 g2713 (.Z(w2896), .A(w2822), .B(w2860), .C(w2821) );
	vdp_and3 g2714 (.Z(w2784), .A(w2860), .B(w2819), .C(w2823) );
	vdp_and3 g2715 (.Z(w2782), .A(w2822), .B(w2818), .C(w2821) );
	vdp_and3 g2716 (.Z(w2780), .A(w2818), .B(w2819), .C(w2823) );
	vdp_and3 g2717 (.Z(w2898), .A(w2822), .B(w2819), .C(w2818) );
	vdp_and3 g2718 (.Z(w2781), .A(w2821), .B(w2823), .C(w2818) );
	vdp_sr_bit g2719 (.Q(w2777), .D(w2824), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2720 (.Q(w2774), .D(w2630), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2721 (.Q(w2825), .D(w2666), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g2722 (.Z(w2776), .A(w2778), .B(w2779), .C(w2773) );
	vdp_and3 g2723 (.Z(w2775), .A(w2773), .B(w2777), .C(w2779) );
	vdp_and3 g2724 (.Z(w2900), .A(w2778), .B(w2779), .C(w2774) );
	vdp_and3 g2725 (.Z(w2771), .A(w2779), .B(w2774), .C(w2777) );
	vdp_and3 g2726 (.Z(w2772), .A(w2773), .B(w2777), .C(w2825) );
	vdp_and3 g2727 (.Z(w2769), .A(w2778), .B(w2825), .C(w2773) );
	vdp_and3 g2728 (.Z(w2899), .A(w2778), .B(w2774), .C(w2825) );
	vdp_and3 g2729 (.Z(w2770), .A(w2825), .B(w2774), .C(w2777) );
	vdp_not g2730 (.nZ(w2859), .A(w2914) );
	vdp_not g2731 (.nZ(w2814), .A(w2816) );
	vdp_not g2732 (.nZ(w2815), .A(w2817) );
	vdp_sr_bit g2733 (.Q(w2816), .D(w2855), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2734 (.Q(w2817), .D(w2853), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2735 (.Q(w2914), .D(w2628), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g2736 (.Z(w2768), .A(w2815), .B(w2859), .C(w2814) );
	vdp_and3 g2737 (.Z(w2767), .A(w2814), .B(w2817), .C(w2859) );
	vdp_and3 g2738 (.A(w2815), .B(w2859), .C(w2816), .Z(w2764) );
	vdp_and3 g2739 (.Z(w2901), .A(w2859), .B(w2816), .C(w2817) );
	vdp_and3 g2740 (.Z(w2763), .A(w2815), .B(w2914), .C(w2814) );
	vdp_and3 g2741 (.Z(w2903), .A(w2814), .B(w2817), .C(w2914) );
	vdp_and3 g2742 (.Z(w2858), .A(w2914), .B(w2816), .C(w2817) );
	vdp_and3 g2743 (.Z(w2902), .A(w2815), .B(w2816), .C(w2914) );
	vdp_aon22 g2744 (.nZ(w2848), .B2(w2761), .B1(w2902), .A2(w2903), .A1(HIGHLIGHT) );
	vdp_aon22 g2745 (.nZ(w2813), .B2(w2761), .B1(w2763), .A2(w2767), .A1(HIGHLIGHT) );
	vdp_aon22 g2746 (.nZ(w2847), .B2(HIGHLIGHT), .B1(w2768), .A2(w2858), .A1(w2766) );
	vdp_and g2747 (.nZ(w2812), .B(HIGHLIGHT), .A(w2763) );
	vdp_and g2748 (.nZ(w2846), .B(HIGHLIGHT), .A(w2902) );
	vdp_and g2749 (.nZ(w2845), .B(HIGHLIGHT), .A(w2764) );
	vdp_aon22 g2750 (.nZ(w2844), .B2(w2765), .B1(w2903), .A2(w2763), .A1(w2765) );
	vdp_aon22 g2751 (.nZ(w2843), .B2(w2761), .B1(w2903), .A2(w2901), .A1(HIGHLIGHT) );
	vdp_aon2222 g2752 (.Z(w2827), .B2(w2765), .B1(w2858), .A2(w2902), .A1(w2765), .D2(w2761), .D1(w2858), .C2(w2858), .C1(HIGHLIGHT) );
	vdp_aon22 g2753 (.Z(w2810), .B2(w2761), .B1(w2767), .A2(w2764), .A1(w2766) );
	vdp_aon22 g2754 (.Z(w2807), .B2(w2761), .B1(w2901), .A2(w2902), .A1(w2766) );
	vdp_and g2755 (.Z(w2811), .B(w2903), .A(w2766) );
	vdp_and g2756 (.Z(w2806), .B(w2766), .A(w2901) );
	vdp_and g2757 (.Z(w2808), .B(w2767), .A(w2766) );
	vdp_aon22 g2758 (.Z(w2805), .B2(w2765), .B1(w2901), .A2(w2764), .A1(w2765) );
	vdp_aon22 g2759 (.Z(w2804), .B2(w2761), .B1(w2764), .A2(w2763), .A1(w2766) );
	vdp_aon2222 g2760 (.Z(w2842), .B2(w2765), .B1(w2767), .A2(w2768), .A1(w2765), .D2(w2761), .D1(w2768), .C2(w2768), .C1(w2766) );
	vdp_not g2761 (.nZ(w2809), .A(w2827) );
	vdp_aon22 g2762 (.nZ(w2841), .B2(w2761), .B1(w2899), .A2(w2772), .A1(HIGHLIGHT) );
	vdp_aon22 g2763 (.nZ(w2840), .B2(w2761), .B1(w2769), .A2(w2775), .A1(HIGHLIGHT) );
	vdp_aon22 g2764 (.nZ(w2803), .B2(HIGHLIGHT), .B1(w2776), .A2(w2770), .A1(w2766) );
	vdp_and g2765 (.nZ(w2802), .B(HIGHLIGHT), .A(w2769) );
	vdp_and g2766 (.nZ(w2801), .B(HIGHLIGHT), .A(w2899) );
	vdp_and g2767 (.nZ(w2800), .B(HIGHLIGHT), .A(w2900) );
	vdp_aon22 g2768 (.nZ(w2799), .B2(w2765), .B1(w2772), .A2(w2769), .A1(w2765) );
	vdp_aon22 g2769 (.nZ(w2798), .B2(w2761), .B1(w2772), .A2(w2771), .A1(HIGHLIGHT) );
	vdp_and g2770 (.Z(w2795), .B(w2772), .A(w2766) );
	vdp_and g2771 (.Z(w2892), .B(w2766), .A(w2771) );
	vdp_and g2772 (.Z(w2794), .B(w2775), .A(w2766) );
	vdp_aon22 g2773 (.Z(w2793), .B2(w2765), .B1(w2771), .A2(w2900), .A1(w2765) );
	vdp_aon22 g2774 (.Z(w2792), .B2(w2761), .B1(w2900), .A2(w2769), .A1(w2766) );
	vdp_aon2222 g2775 (.Z(w2893), .B2(w2765), .B1(w2775), .A2(w2776), .A1(w2765), .D2(w2761), .D1(w2776), .C2(w2776), .C1(w2766) );
	vdp_aon22 g2776 (.nZ(w2789), .B2(w2761), .B1(w2898), .A2(w2781), .A1(HIGHLIGHT) );
	vdp_aon22 g2777 (.nZ(w2839), .B2(w2761), .B1(w2782), .A2(w2897), .A1(HIGHLIGHT) );
	vdp_aon22 g2778 (.nZ(w2835), .B2(HIGHLIGHT), .B1(w2896), .A2(w2780), .A1(w2766) );
	vdp_and g2779 (.nZ(w2836), .B(HIGHLIGHT), .A(w2782) );
	vdp_and g2780 (.nZ(w2837), .B(HIGHLIGHT), .A(w2898) );
	vdp_and g2781 (.nZ(w2834), .B(HIGHLIGHT), .A(w2895) );
	vdp_aon22 g2782 (.nZ(w2838), .B2(w2765), .B1(w2781), .A2(w2782), .A1(w2765) );
	vdp_aon22 g2783 (.nZ(w2894), .B2(w2761), .B1(w2781), .A2(w2784), .A1(HIGHLIGHT) );
	vdp_aon2222 g2784 (.Z(w2783), .B2(w2765), .B1(w2780), .A2(w2898), .A1(w2765), .D2(w2761), .D1(w2780), .C2(w2780), .C1(HIGHLIGHT) );
	vdp_aon22 g2785 (.Z(w2787), .B2(w2761), .B1(w2897), .A2(w2895), .A1(w2766) );
	vdp_aon22 g2786 (.Z(w2788), .B2(w2765), .B1(w2784), .A2(w2895), .A1(w2765) );
	vdp_aon22 g2787 (.Z(w2833), .B2(w2761), .B1(w2784), .A2(w2898), .A1(w2766) );
	vdp_and g2788 (.Z(w2832), .B(w2766), .A(w2784) );
	vdp_and g2789 (.Z(w2831), .B(w2897), .A(w2766) );
	vdp_and g2790 (.Z(w2830), .B(w2766), .A(w2781) );
	vdp_aon22 g2791 (.Z(w2828), .B2(w2761), .B1(w2895), .A2(w2782), .A1(w2766) );
	vdp_aon2222 g2792 (.Z(w2829), .B2(w2765), .B1(w2897), .A2(w2896), .A1(w2765), .D2(w2761), .D1(w2896), .C2(w2896), .C1(w2766) );
	vdp_nor3 g2793 (.Z(w2761), .A(w2765), .B(SHADOW), .C(HIGHLIGHT) );
	vdp_and g2794 (.Z(w2766), .A(SHADOW), .B(w2786) );
	vdp_bufif0 g2795 (.A(w2684), .nE(w2691), .Z(COL[0]) );
	vdp_bufif0 g2796 (.A(w2876), .nE(w2691), .Z(COL[1]) );
	vdp_bufif0 g2797 (.A(w2686), .nE(w2691), .Z(COL[2]) );
	vdp_bufif0 g2798 (.A(w2690), .nE(w2691), .Z(COL[3]) );
	vdp_bufif0 g2799 (.A(w2704), .nE(w2691), .Z(COL[4]) );
	vdp_bufif0 g2800 (.A(w2875), .nE(w2691), .Z(COL[5]) );
	vdp_and g2801 (.Z(w2875), .A(M5), .B(w2702) );
	vdp_or g2802 (.Z(w2704), .A(w2674), .B(w2694) );
	vdp_not g2803 (.nZ(w2567), .A(M5) );
	vdp_not g2804 (.nZ(w2672), .A(w2874) );
	vdp_not g2805 (.nZ(w2673), .A(w2675) );
	vdp_not g2806 (.nZ(w2674), .A(M5) );
	vdp_not g2807 (.nZ(w2670), .A(w2676) );
	vdp_not g2808 (.nZ(w2691), .A(w2679) );
	vdp_comp_strong g2809 (.nZ(w2682), .Z(w2692), .A(w811) );
	vdp_not g2810 (.nZ(w2680), .A(w86) );
	vdp_not g2811 (.nZ(w2887), .A(w18) );
	vdp_aon222 g2812 (.Z(w2871), .B2(w2672), .A2(w2673), .A1(VRAMA[0]), .B1(VRAMA[1]), .C2(w2670), .C1(COL[0]) );
	vdp_aon222 g2813 (.Z(w2888), .B2(w2672), .A2(w2673), .A1(VRAMA[1]), .B1(VRAMA[2]), .C2(w2670), .C1(COL[1]) );
	vdp_aon222 g2814 (.Z(w2685), .B2(w2672), .A2(w2673), .A1(VRAMA[2]), .B1(VRAMA[3]), .C2(w2670), .C1(COL[2]) );
	vdp_aon222 g2815 (.Z(w2695), .B2(w2672), .A2(w2673), .A1(VRAMA[3]), .B1(VRAMA[4]), .C2(w2670), .C1(COL[3]) );
	vdp_aon222 g2816 (.Z(w2701), .B2(w2672), .A2(w2673), .A1(VRAMA[4]), .B1(VRAMA[5]), .C2(w2670), .C1(COL[4]) );
	vdp_aon222 g2817 (.Z(w2760), .B2(w2672), .A2(w2673), .A1(1'b0), .B1(VRAMA[6]), .C2(w2670), .C1(COL[5]) );
	vdp_nand g2818 (.Z(w2874), .A(w2676), .B(M5) );
	vdp_nand g2819 (.Z(w2675), .A(w2676), .B(w2674) );
	vdp_and g2820 (.Z(w2706), .A(w2707), .B(w2922) );
	vdp_aon222 g2821 (.Z(w2922), .B2(w2917), .A2(w2712), .A1(w2667), .B1(w2714), .C2(w2916), .C1(w2735) );
	vdp_not g2822 (.nZ(w2917), .A(w2870) );
	vdp_not g2823 (.nZ(w2916), .A(w2668) );
	vdp_not g2824 (.nZ(w2740), .A(w2725) );
	vdp_nor g2825 (.Z(w2714), .A(w2668), .B(w2863) );
	vdp_nor g2826 (.Z(w2870), .A(w2735), .B(w2734) );
	vdp_and g2827 (.Z(w2713), .A(w2708), .B(w2748) );
	vdp_and g2828 (.Z(w2712), .A(w2725), .B(w2739) );
	vdp_and g2829 (.Z(w2742), .A(w2739), .B(w2740) );
	vdp_or g2830 (.Z(w2863), .A(w2743), .B(w2742) );
	vdp_or g2831 (.Z(w2711), .A(w2667), .B(w2668) );
	vdp_and g2832 (.Z(w2681), .A(w2707), .B(w2680) );
	vdp_and g2833 (.Z(w2852), .A(w2708), .B(w2745) );
	vdp_and g2834 (.Z(w2862), .A(w2709), .B(w2747) );
	vdp_not g2835 (.nZ(w2753), .A(w86) );
	vdp_or g2836 (.Z(w2715), .A(w2746), .B(w2732) );
	vdp_not g2837 (.nZ(w2920), .A(w2709) );
	vdp_not g2838 (.nZ(w2850), .A(w2609) );
	vdp_not g2839 (.nZ(w2737), .A(w2726) );
	vdp_not g2840 (.nZ(w2736), .A(w2727) );
	vdp_not g2841 (.nZ(w2741), .A(w2610) );
	vdp_and g2842 (.Z(w2758), .A(w2709), .B(w2744) );
	vdp_and g2843 (.Z(w2738), .A(w2710), .B(w2750) );
	vdp_not g2844 (.nZ(w2861), .A(w83) );
	vdp_not g2845 (.nZ(w2868), .A(w84) );
	vdp_and g2846 (.Z(w2743), .A(w2868), .B(w83) );
	vdp_and g2847 (.Z(w2746), .A(w2861), .B(w84) );
	vdp_and g2848 (.Z(w2757), .A(w83), .B(w84) );
	vdp_or3 g2849 (.Z(w2676), .A(w93), .B(w1435), .C(w1434) );
	vdp_and3 g2850 (.Z(w2867), .A(w2710), .B(w2709), .C(w2747) );
	vdp_and3 g2851 (.Z(w2745), .A(w2736), .B(w2726), .C(w2610) );
	vdp_and3 g2852 (.Z(w2744), .A(w2737), .B(w2727), .C(w2741) );
	vdp_and3 g2853 (.Z(w2750), .A(w2736), .B(w2726), .C(w2741) );
	vdp_and3 g2854 (.Z(w2747), .A(w2726), .B(w2727), .C(w2741) );
	vdp_and g2855 (.Z(w2857), .A(M5), .B(S_TE) );
	vdp_or g2856 (.Z(w2708), .A(w2850), .B(w2725) );
	vdp_and3 g2857 (.Z(w2718), .A(w2712), .B(w2668), .C(w2870) );
	vdp_and3 g2858 (.Z(w2866), .A(w2710), .B(w2708), .C(w2745) );
	vdp_and3 g2859 (.Z(w2865), .A(w2710), .B(w2708), .C(w2750) );
	vdp_and3 g2860 (.Z(w2732), .A(w2731), .B(w2681), .C(w2920) );
	vdp_and3 g2861 (.Z(w2725), .A(w2711), .B(w2728), .C(w2857) );
	vdp_and3 g2862 (.Z(w2754), .A(w2709), .B(w2708), .C(w2748) );
	vdp_and3 g2863 (.Z(w2919), .A(w2709), .B(w2708), .C(w2744) );
	vdp_and3 g2864 (.Z(w2751), .A(w2710), .B(w2709), .C(w2708) );
	vdp_and3 g2865 (.Z(w2752), .A(w2681), .B(w2749), .C(w2918) );
	vdp_and g2866 (.Z(w2717), .A(w2851), .B(w2864) );
	vdp_not g2867 (.nZ(w2755), .A(w2681) );
	vdp_not g2868 (.nZ(w2918), .A(w2710) );
	vdp_or g2869 (.Z(w2716), .A(w2757), .B(w2752) );
	vdp_or g2870 (.Z(w2864), .A(w2755), .B(w2751) );
	vdp_not g2871 (.nZ(w2879), .A(M5) );
	vdp_notif0 g2872 (.A(w2912), .nE(w2649), .nZ(w300) );
	vdp_notif0 g2873 (.nZ(RD_DATA[2]), .A(w2911), .nE(w2649) );
	vdp_notif0 g2874 (.nZ(RD_DATA[1]), .A(w2910), .nE(w2649) );
	vdp_notif0 g2875 (.nZ(AD_DATA[7]), .A(w2909), .nE(w2649) );
	vdp_notif0 g2876 (.nZ(AD_DATA[6]), .A(w2908), .nE(w2649) );
	vdp_notif0 g2877 (.nZ(AD_DATA[5]), .A(w2907), .nE(w2649) );
	vdp_notif0 g2878 (.nZ(AD_DATA[3]), .A(w2906), .nE(w2649) );
	vdp_notif0 g2879 (.nZ(AD_DATA[2]), .A(w2905), .nE(w2649) );
	vdp_notif0 g2880 (.nZ(AD_DATA[1]), .A(w2904), .nE(w2649) );
	vdp_notif0 g2881 (.nZ(DB[1]), .A(w2642), .nE(w2633) );
	vdp_notif0 g2882 (.nZ(DB[0]), .A(w2641), .nE(w2633) );
	vdp_notif0 g2883 (.nZ(DB[2]), .A(w2853), .nE(w2633) );
	vdp_notif0 g2884 (.nZ(DB[5]), .A(w2824), .nE(w2633) );
	vdp_notif0 g2885 (.nZ(DB[8]), .A(w2640), .nE(w2633) );
	vdp_notif0 g2886 (.nZ(DB[10]), .A(w2820), .nE(w2633) );
	vdp_notif0 g2887 (.nZ(DB[9]), .A(w2665), .nE(w2633) );
	vdp_notif0 g2888 (.nZ(DB[7]), .A(w2666), .nE(w2633) );
	vdp_notif0 g2889 (.nZ(DB[6]), .A(w2630), .nE(w2633) );
	vdp_notif0 g2890 (.nZ(DB[4]), .A(w2628), .nE(w2633) );
	vdp_comp_we g2891 (.A(M5), .nZ(w2623), .Z(w2622) );
	vdp_notif0 g2892 (.nZ(DB[3]), .A(w2855), .nE(w2633) );
	vdp_not g2893 (.A(w73), .nZ(w2633) );
	vdp_and g2894 (.Z(w2624), .A(w2625), .B(w2620) );
	vdp_and3 g2895 (.Z(w2855), .A(w82), .B(w2625), .C(w2854) );
	vdp_and3 g2896 (.Z(w2628), .A(w82), .B(w2625), .C(w2890) );
	vdp_and3 g2897 (.Z(w2630), .A(w82), .B(w2625), .C(w2629) );
	vdp_and3 g2898 (.Z(w2666), .A(w82), .B(w2625), .C(w2632) );
	vdp_and3 g2899 (.Z(w2665), .A(w82), .B(w2625), .C(w2635) );
	vdp_and3 g2900 (.Z(w2820), .A(w82), .B(w2625), .C(w2638) );
	vdp_and3 g2901 (.Z(w2640), .A(M5), .B(w2625), .C(w2639) );
	vdp_and3 g2902 (.Z(w2824), .A(M5), .B(w2625), .C(w2646) );
	vdp_and3 g2903 (.Z(w2853), .A(M5), .B(w2625), .C(w2631) );
	vdp_comp_strong g2904 (.nZ(w2644), .A(w2643), .Z(w2647) );
	vdp_and g2905 (.Z(w2643), .A(w2645), .B(HCLK1) );
	vdp_not g2906 (.nZ(w2649), .A(w2913) );
	vdp_aon22 g2907 (.Z(w2878), .B2(FIFOo[5]), .A2(FIFOo[7]), .A1(w2697), .B1(w2696) );
	vdp_aon22 g2908 (.Z(w2660), .B2(FIFOo[4]), .A2(FIFOo[6]), .A1(w2697), .B1(w2696) );
	vdp_aon22 g2909 (.Z(w2657), .B2(FIFOo[3]), .A2(FIFOo[5]), .A1(w2697), .B1(w2696) );
	vdp_aon22 g2910 (.Z(w2656), .B2(FIFOo[2]), .A2(FIFOo[3]), .A1(w2697), .B1(w2696) );
	vdp_aon22 g2911 (.Z(w2655), .B2(FIFOo[1]), .A2(FIFOo[2]), .A1(w2697), .B1(w2696) );
	vdp_aon22 g2912 (.Z(w2659), .B2(FIFOo[0]), .A2(FIFOo[1]), .A1(w2697), .B1(w2696) );
	vdp_comp_we g2913 (.Z(w2697), .nZ(w2696), .A(M5) );
	vdp_aon22 g2914 (.Z(w2688), .B2(w2879), .A2(M5), .A1(w2856), .B1(w17) );
	vdp_aon22 g2915 (.Z(COL[7]), .B2(w2719), .A2(w2705), .A1(w86), .B1(w2753) );
	vdp_aon22 g2916 (.Z(w114), .B2(w2733), .A2(w2849), .A1(w86), .B1(w2753) );
	vdp_and3 g2917 (.Z(w2739), .A(w2681), .B(w2609), .C(w2921) );
	vdp_aon22 g2918 (.Z(w2748), .B2(w2736), .A2(w2727), .A1(w2610), .B1(w2737) );
	vdp_aon22 g2919 (.Z(w2632), .B2(w2646), .A2(w2636), .A1(w2622), .B1(w2623) );
	vdp_aon22 g2920 (.Z(w2629), .B2(w2626), .A2(w2627), .A1(w2622), .B1(w2623) );
	vdp_aon22 g2921 (.Z(w2854), .B2(w2631), .A2(w2621), .A1(w2622), .B1(w2623) );
	vdp_aon22 g2922 (.Z(w2890), .B2(w2621), .A2(w2626), .A1(w2622), .B1(w2623) );
	vdp_aon22 g2923 (.Z(w2635), .B2(w2627), .A2(w2634), .A1(w2622), .B1(w2623) );
	vdp_aon22 g2924 (.Z(w2638), .B2(w2636), .A2(w2637), .A1(w2622), .B1(w2623) );
	vdp_and4 g2925 (.Z(w2734), .A(w2737), .B(w2610), .C(w2857), .D(w2736) );
	vdp_or5 g2926 (.Z(w2731), .A(w2713), .B(w2744), .C(w2747), .D(w2866), .E(w2865) );
	vdp_or5 g2927 (.Z(w2749), .A(w2754), .B(w2750), .C(w2852), .D(w2862), .E(w2919) );
	vdp_or5 g2928 (.Z(w2921), .A(w2745), .B(w2748), .C(w2758), .D(w2738), .E(w2867) );
	vdp_nor4 g2929 (.Z(w2698), .A(COL[2]), .B(COL[3]), .C(COL[1]), .D(COL[0]) );
	vdp_nor g2930 (.Z(w2851), .A(w83), .B(w84) );
	vdp_nor g2931 (.Z(w2709), .A(w2869), .B(w2873) );
	vdp_nor g2932 (.Z(w2869), .A(w2609), .B(M5) );
	vdp_nand g2933 (.Z(w2710), .A(M5), .B(w2872) );
	vdp_nand g2934 (.Z(w2721), .A(SPR_PRIO), .B(w18) );
	vdp_and4 g2935 (.Z(w2735), .A(w2736), .B(w2857), .C(w2737), .D(w2741) );
	vdp_aoi21 g2936 (.Z(w2889), .B(w2624), .A2(w2887), .A1(w2671) );
	vdp_nor g2937 (.Z(w2759), .A(w20), .B(w19) );
	vdp_n_fet g2938 (.A(w2679), .Z(COL[6]) );
	vdp_slatch g2939 (.Q(w3997), .D(S[3]), .C(w3049), .nC(w3039) );
	vdp_slatch g2940 (.Q(w3999), .D(S[3]), .C(w3030), .nC(w3029) );
	vdp_slatch g2941 (.Q(w4001), .D(S[3]), .C(w3031), .nC(w3027) );
	vdp_slatch g2942 (.Q(w4003), .D(S[3]), .C(w3048), .nC(w3040) );
	vdp_slatch g2943 (.Q(w4005), .D(S[7]), .C(w3049), .nC(w3039) );
	vdp_slatch g2944 (.Q(w4008), .D(S[7]), .C(w3030), .nC(w3029) );
	vdp_slatch g2945 (.Q(w4007), .D(S[7]), .C(w3031), .nC(w3027) );
	vdp_slatch g2946 (.Q(w4012), .D(S[7]), .C(w3048), .nC(w3040) );
	vdp_slatch g2947 (.Q(w4011), .D(S[2]), .C(w3049), .nC(w3039) );
	vdp_slatch g2948 (.Q(w4018), .D(S[2]), .C(w3030), .nC(w3029) );
	vdp_slatch g2949 (.Q(w4017), .D(S[2]), .C(w3031), .nC(w3027) );
	vdp_slatch g2950 (.Q(w4020), .D(S[2]), .C(w3048), .nC(w3040) );
	vdp_slatch g2951 (.Q(w4019), .D(S[6]), .C(w3049), .nC(w3039) );
	vdp_slatch g2952 (.Q(w4024), .D(S[6]), .C(w3030), .nC(w3029) );
	vdp_slatch g2953 (.Q(w4023), .D(S[6]), .C(w3031), .nC(w3027) );
	vdp_slatch g2954 (.Q(w4028), .D(S[6]), .C(w3048), .nC(w3040) );
	vdp_slatch g2955 (.Q(w4027), .D(S[1]), .C(w3049), .nC(w3039) );
	vdp_slatch g2956 (.Q(w4032), .D(S[1]), .C(w3030), .nC(w3029) );
	vdp_slatch g2957 (.Q(w4031), .D(S[1]), .C(w3031), .nC(w3027) );
	vdp_slatch g2958 (.Q(w4036), .D(S[1]), .C(w3048), .nC(w3040) );
	vdp_slatch g2959 (.Q(w4035), .D(S[5]), .C(w3049), .nC(w3039) );
	vdp_slatch g2960 (.Q(w4040), .D(S[5]), .C(w3030), .nC(w3029) );
	vdp_slatch g2961 (.Q(w4039), .D(S[5]), .C(w3031), .nC(w3027) );
	vdp_slatch g2962 (.Q(w4044), .D(S[5]), .C(w3048), .nC(w3040) );
	vdp_slatch g2963 (.Q(w4043), .D(S[0]), .C(w3049), .nC(w3039) );
	vdp_slatch g2964 (.Q(w4048), .D(S[0]), .C(w3030), .nC(w3029) );
	vdp_slatch g2965 (.Q(w4047), .D(S[0]), .C(w3031), .nC(w3027) );
	vdp_slatch g2966 (.Q(w4052), .D(S[0]), .C(w3048), .nC(w3040) );
	vdp_slatch g2967 (.Q(w4051), .D(S[4]), .C(w3049), .nC(w3039) );
	vdp_slatch g2968 (.Q(w4056), .D(S[4]), .C(w3030), .nC(w3029) );
	vdp_slatch g2969 (.Q(w4055), .D(S[4]), .C(w3031), .nC(w3027) );
	vdp_slatch g2970 (.Q(w4059), .D(S[4]), .C(w3048), .nC(w3040) );
	vdp_slatch g2971 (.Q(w3998), .D(w3997), .C(w3018), .nC(w3036) );
	vdp_slatch g2972 (.Q(w4000), .D(w3999), .C(w3037), .nC(w3028) );
	vdp_slatch g2973 (.Q(w4002), .D(w4001), .C(w3038), .nC(w3026) );
	vdp_slatch g2974 (.Q(w4004), .D(w4003), .C(w3034), .nC(w3035) );
	vdp_slatch g2975 (.Q(w4006), .D(w4005), .C(w3018), .nC(w3036) );
	vdp_slatch g2976 (.Q(w4010), .D(w4008), .C(w3037), .nC(w3028) );
	vdp_slatch g2977 (.Q(w4009), .D(w4007), .C(w3038), .nC(w3026) );
	vdp_slatch g2978 (.Q(w4014), .D(w4012), .C(w3034), .nC(w3035) );
	vdp_slatch g2979 (.Q(w4013), .D(w4011), .C(w3018), .nC(w3036) );
	vdp_slatch g2980 (.Q(w4016), .D(w4018), .C(w3037), .nC(w3028) );
	vdp_slatch g2981 (.Q(w4015), .D(w4017), .C(w3038), .nC(w3026) );
	vdp_slatch g2982 (.Q(w4022), .D(w4020), .C(w3034), .nC(w3035) );
	vdp_slatch g2983 (.Q(w4021), .D(w4019), .C(w3018), .nC(w3036) );
	vdp_slatch g2984 (.Q(w4026), .D(w4024), .C(w3037), .nC(w3028) );
	vdp_slatch g2985 (.Q(w4025), .D(w4023), .C(w3038), .nC(w3026) );
	vdp_slatch g2986 (.Q(w4030), .D(w4028), .C(w3034), .nC(w3035) );
	vdp_slatch g2987 (.Q(w4029), .D(w4027), .C(w3018), .nC(w3036) );
	vdp_slatch g2988 (.Q(w4034), .D(w4032), .C(w3037), .nC(w3028) );
	vdp_slatch g2989 (.Q(w4033), .D(w4031), .C(w3038), .nC(w3026) );
	vdp_slatch g2990 (.Q(w4038), .D(w4036), .C(w3034), .nC(w3035) );
	vdp_slatch g2991 (.Q(w4037), .D(w4035), .C(w3018), .nC(w3036) );
	vdp_slatch g2992 (.Q(w4042), .D(w4040), .C(w3037), .nC(w3028) );
	vdp_slatch g2993 (.Q(w4041), .D(w4039), .C(w3038), .nC(w3026) );
	vdp_slatch g2994 (.Q(w4046), .D(w4044), .C(w3034), .nC(w3035) );
	vdp_slatch g2995 (.Q(w4045), .D(w4043), .C(w3018), .nC(w3036) );
	vdp_slatch g2996 (.Q(w4050), .D(w4048), .C(w3037), .nC(w3028) );
	vdp_slatch g2997 (.Q(w4049), .D(w4047), .C(w3038), .nC(w3026) );
	vdp_slatch g2998 (.Q(w4054), .D(w4052), .C(w3034), .nC(w3035) );
	vdp_slatch g2999 (.Q(w4053), .D(w4051), .C(w3018), .nC(w3036) );
	vdp_slatch g3000 (.Q(w4058), .D(w4056), .C(w3037), .nC(w3028) );
	vdp_slatch g3001 (.Q(w4057), .D(w4055), .C(w3038), .nC(w3026) );
	vdp_slatch g3002 (.Q(w4060), .D(w4059), .C(w3034), .nC(w3035) );
	vdp_slatch g3003 (.Q(w3076), .D(w3998), .C(w3041), .nC(w3067) );
	vdp_slatch g3004 (.Q(w3075), .D(w4000), .C(w3019), .nC(w3077) );
	vdp_slatch g3005 (.Q(w3074), .D(w4002), .C(w3032), .nC(w3078) );
	vdp_slatch g3006 (.Q(w3073), .D(w4004), .C(w3033), .nC(w3006) );
	vdp_slatch g3007 (.Q(w3072), .D(w4006), .C(w3041), .nC(w3067) );
	vdp_slatch g3008 (.Q(w3071), .D(w4010), .C(w3019), .nC(w3077) );
	vdp_slatch g3009 (.Q(w3070), .D(w4009), .C(w3032), .nC(w3078) );
	vdp_slatch g3010 (.Q(w3069), .D(w4014), .C(w3033), .nC(w3006) );
	vdp_slatch g3011 (.Q(w3068), .D(w4013), .C(w3041), .nC(w3067) );
	vdp_slatch g3012 (.Q(w3081), .D(w4016), .C(w3019), .nC(w3077) );
	vdp_slatch g3013 (.Q(w3085), .D(w4015), .C(w3032), .nC(w3078) );
	vdp_slatch g3014 (.Q(w3084), .D(w4022), .C(w3033), .nC(w3006) );
	vdp_slatch g3015 (.Q(w3083), .D(w4021), .C(w3041), .nC(w3067) );
	vdp_slatch g3016 (.Q(w3079), .D(w4026), .C(w3019), .nC(w3077) );
	vdp_slatch g3017 (.Q(w3080), .D(w4025), .C(w3032), .nC(w3078) );
	vdp_slatch g3018 (.D(w4030), .Q(w3082), .C(w3033), .nC(w3006) );
	vdp_slatch g3019 (.Q(w3086), .D(w4029), .C(w3041), .nC(w3067) );
	vdp_slatch g3020 (.Q(w3087), .D(w4034), .C(w3019), .nC(w3077) );
	vdp_slatch g3021 (.Q(w3089), .D(w4033), .C(w3032), .nC(w3078) );
	vdp_slatch g3022 (.Q(w3088), .D(w4038), .C(w3033), .nC(w3006) );
	vdp_slatch g3023 (.Q(w3130), .D(w4037), .C(w3041), .nC(w3067) );
	vdp_slatch g3024 (.Q(w3131), .D(w4042), .C(w3019), .nC(w3077) );
	vdp_slatch g3025 (.Q(w3127), .D(w4041), .C(w3032), .nC(w3078) );
	vdp_slatch g3026 (.Q(w3122), .D(w4046), .C(w3033), .nC(w3006) );
	vdp_slatch g3027 (.Q(w3134), .D(w4045), .C(w3041), .nC(w3067) );
	vdp_slatch g3028 (.Q(w3133), .D(w4050), .C(w3019), .nC(w3077) );
	vdp_slatch g3029 (.Q(w3132), .D(w4049), .C(w3032), .nC(w3078) );
	vdp_slatch g3030 (.Q(w3129), .D(w4054), .C(w3033), .nC(w3006) );
	vdp_slatch g3031 (.Q(w3115), .D(w4053), .C(w3041), .nC(w3067) );
	vdp_slatch g3032 (.Q(w3114), .D(w4058), .C(w3019), .nC(w3077) );
	vdp_slatch g3033 (.Q(w3116), .D(w4057), .C(w3032), .nC(w3078) );
	vdp_slatch g3034 (.Q(w3117), .D(w4060), .C(w3033), .nC(w3006) );
	vdp_slatch g3035 (.Q(w3193), .D(w4281), .C(w3189), .nC(w3191) );
	vdp_slatch g3036 (.Q(w3194), .D(w4282), .C(w3188), .nC(w3199) );
	vdp_slatch g3037 (.Q(w3195), .D(w4284), .C(w3187), .nC(w3200) );
	vdp_slatch g3038 (.Q(w3196), .D(w4283), .C(w3186), .nC(w3192) );
	vdp_slatch g3039 (.Q(w3197), .D(w4116), .C(w3189), .nC(w3191) );
	vdp_slatch g3040 (.Q(w3198), .D(w4115), .C(w3188), .nC(w3199) );
	vdp_slatch g3041 (.Q(w3204), .D(w4110), .C(w3187), .nC(w3200) );
	vdp_slatch g3042 (.Q(w3205), .D(w4109), .C(w3186), .nC(w3192) );
	vdp_slatch g3043 (.Q(w3206), .D(w4106), .C(w3189), .nC(w3191) );
	vdp_slatch g3044 (.Q(w3207), .D(w4105), .C(w3188), .nC(w3199) );
	vdp_slatch g3045 (.Q(w3208), .D(w4104), .C(w3187), .nC(w3200) );
	vdp_slatch g3046 (.Q(w3203), .D(w4101), .C(w3186), .nC(w3192) );
	vdp_slatch g3047 (.Q(w3209), .D(w4098), .C(w3189), .nC(w3191) );
	vdp_slatch g3048 (.Q(w3210), .D(w4099), .C(w3188), .nC(w3199) );
	vdp_slatch g3049 (.Q(w3211), .D(w4094), .C(w3187), .nC(w3200) );
	vdp_slatch g3050 (.Q(w3212), .D(w4095), .C(w3186), .nC(w3192) );
	vdp_slatch g3051 (.Q(w3138), .D(w4092), .C(w3189), .nC(w3191) );
	vdp_slatch g3052 (.Q(w3885), .D(w4091), .C(w3188), .nC(w3199) );
	vdp_slatch g3053 (.Q(w3140), .D(w4088), .C(w3187), .nC(w3200) );
	vdp_slatch g3054 (.Q(w3141), .D(w4087), .C(w3186), .nC(w3192) );
	vdp_slatch g3055 (.Q(w3213), .D(w4084), .C(w3189), .nC(w3191) );
	vdp_slatch g3056 (.Q(w3139), .D(w4083), .C(w3188), .nC(w3199) );
	vdp_slatch g3057 (.Q(w3119), .D(w4080), .C(w3187), .nC(w3200) );
	vdp_slatch g3058 (.Q(w3142), .D(w4079), .C(w3186), .nC(w3192) );
	vdp_slatch g3059 (.Q(w3145), .D(w4076), .C(w3189), .nC(w3191) );
	vdp_slatch g3060 (.Q(w3153), .D(w4075), .C(w3188), .nC(w3199) );
	vdp_slatch g3061 (.Q(w3152), .D(w4072), .C(w3187), .nC(w3200) );
	vdp_slatch g3062 (.Q(w3151), .D(w4071), .C(w3186), .nC(w3192) );
	vdp_slatch g3063 (.Q(w3149), .D(w4068), .C(w3189), .nC(w3191) );
	vdp_slatch g3064 (.Q(w3143), .D(w4067), .C(w3188), .nC(w3199) );
	vdp_slatch g3065 (.Q(w3150), .D(w4064), .C(w3187), .nC(w3200) );
	vdp_slatch g3066 (.Q(w3144), .D(w4063), .C(w3186), .nC(w3192) );
	vdp_slatch g3067 (.Q(w4281), .D(w4119), .C(w3190), .nC(w3177) );
	vdp_slatch g3068 (.Q(w4282), .D(w4120), .C(w2998), .nC(w3178) );
	vdp_slatch g3069 (.Q(w4284), .D(w4118), .C(w3184), .nC(w2986) );
	vdp_slatch g3070 (.Q(w4283), .D(w4117), .C(w3185), .nC(w2987) );
	vdp_slatch g3071 (.Q(w4116), .D(w4114), .C(w3190), .nC(w3177) );
	vdp_slatch g3072 (.Q(w4115), .D(w4113), .C(w2998), .nC(w3178) );
	vdp_slatch g3073 (.Q(w4110), .D(w4112), .C(w3184), .nC(w2986) );
	vdp_slatch g3074 (.Q(w4109), .D(w4111), .C(w3185), .nC(w2987) );
	vdp_slatch g3075 (.Q(w4106), .D(w4108), .C(w3190), .nC(w3177) );
	vdp_slatch g3076 (.Q(w4105), .D(w4107), .C(w2998), .nC(w3178) );
	vdp_slatch g3077 (.Q(w4104), .D(w4102), .C(w3184), .nC(w2986) );
	vdp_slatch g3078 (.Q(w4101), .D(w4103), .C(w3185), .nC(w2987) );
	vdp_slatch g3079 (.Q(w4098), .D(w4100), .C(w3190), .nC(w3177) );
	vdp_slatch g3080 (.Q(w4099), .D(w4097), .C(w2998), .nC(w3178) );
	vdp_slatch g3081 (.Q(w4094), .D(w4096), .C(w3184), .nC(w2986) );
	vdp_slatch g3082 (.Q(w4095), .D(w4093), .C(w3185), .nC(w2987) );
	vdp_slatch g3083 (.Q(w4092), .D(w4090), .C(w3190), .nC(w3177) );
	vdp_slatch g3084 (.Q(w4091), .D(w4089), .C(w2998), .nC(w3178) );
	vdp_slatch g3085 (.Q(w4088), .D(w4086), .C(w3184), .nC(w2986) );
	vdp_slatch g3086 (.Q(w4087), .D(w4085), .C(w3185), .nC(w2987) );
	vdp_slatch g3087 (.Q(w4084), .D(w4082), .C(w3190), .nC(w3177) );
	vdp_slatch g3088 (.Q(w4083), .D(w4081), .C(w2998), .nC(w3178) );
	vdp_slatch g3089 (.Q(w4080), .D(w4078), .C(w3184), .nC(w2986) );
	vdp_slatch g3090 (.Q(w4079), .D(w4077), .C(w3185), .nC(w2987) );
	vdp_slatch g3091 (.Q(w4076), .D(w4074), .C(w3190), .nC(w3177) );
	vdp_slatch g3092 (.Q(w4075), .D(w4073), .C(w2998), .nC(w3178) );
	vdp_slatch g3093 (.Q(w4072), .D(w4070), .C(w3184), .nC(w2986) );
	vdp_slatch g3094 (.Q(w4071), .D(w4069), .C(w3185), .nC(w2987) );
	vdp_slatch g3095 (.Q(w4068), .D(w4066), .C(w3190), .nC(w3177) );
	vdp_slatch g3096 (.Q(w4067), .D(w4065), .C(w2998), .nC(w3178) );
	vdp_slatch g3097 (.Q(w4064), .D(w4062), .C(w3184), .nC(w2986) );
	vdp_slatch g3098 (.Q(w4063), .D(w4061), .C(w3185), .nC(w2987) );
	vdp_slatch g3099 (.Q(w4119), .D(S[3]), .C(w2951), .nC(w2984) );
	vdp_slatch g3100 (.Q(w4120), .D(S[3]), .C(w2955), .nC(w2988) );
	vdp_slatch g3101 (.Q(w4118), .D(S[3]), .C(w2958), .nC(w2985) );
	vdp_slatch g3102 (.Q(w4117), .D(S[3]), .C(w2960), .nC(w2983) );
	vdp_slatch g3103 (.Q(w4114), .D(S[7]), .C(w2951), .nC(w2984) );
	vdp_slatch g3104 (.Q(w4113), .D(S[7]), .C(w2955), .nC(w2988) );
	vdp_slatch g3105 (.Q(w4112), .D(S[7]), .C(w2958), .nC(w2985) );
	vdp_slatch g3106 (.Q(w4111), .D(S[7]), .C(w2960), .nC(w2983) );
	vdp_slatch g3107 (.Q(w4108), .D(S[2]), .C(w2951), .nC(w2984) );
	vdp_slatch g3108 (.Q(w4107), .D(S[2]), .C(w2955), .nC(w2988) );
	vdp_slatch g3109 (.Q(w4102), .D(S[2]), .C(w2958), .nC(w2985) );
	vdp_slatch g3110 (.Q(w4103), .D(S[2]), .C(w2960), .nC(w2983) );
	vdp_slatch g3111 (.Q(w4100), .D(S[6]), .C(w2951), .nC(w2984) );
	vdp_slatch g3112 (.Q(w4097), .D(S[6]), .C(w2955), .nC(w2988) );
	vdp_slatch g3113 (.Q(w4096), .D(S[6]), .C(w2958), .nC(w2985) );
	vdp_slatch g3114 (.Q(w4093), .D(S[6]), .C(w2960), .nC(w2983) );
	vdp_slatch g3115 (.Q(w4090), .D(S[1]), .C(w2951), .nC(w2984) );
	vdp_slatch g3116 (.Q(w4089), .D(S[1]), .C(w2955), .nC(w2988) );
	vdp_slatch g3117 (.Q(w4086), .D(S[1]), .C(w2958), .nC(w2985) );
	vdp_slatch g3118 (.Q(w4085), .D(S[1]), .C(w2960), .nC(w2983) );
	vdp_slatch g3119 (.Q(w4082), .D(S[5]), .C(w2951), .nC(w2984) );
	vdp_slatch g3120 (.Q(w4081), .D(S[5]), .C(w2955), .nC(w2988) );
	vdp_slatch g3121 (.Q(w4078), .D(S[5]), .C(w2958), .nC(w2985) );
	vdp_slatch g3122 (.Q(w4077), .D(S[5]), .C(w2960), .nC(w2983) );
	vdp_slatch g3123 (.Q(w4074), .D(S[0]), .C(w2951), .nC(w2984) );
	vdp_slatch g3124 (.Q(w4073), .D(S[0]), .C(w2955), .nC(w2988) );
	vdp_slatch g3125 (.Q(w4070), .D(S[0]), .C(w2958), .nC(w2985) );
	vdp_slatch g3126 (.Q(w4069), .D(S[0]), .C(w2960), .nC(w2983) );
	vdp_slatch g3127 (.Q(w4066), .D(S[4]), .C(w2951), .nC(w2984) );
	vdp_slatch g3128 (.Q(w4065), .D(S[4]), .C(w2955), .nC(w2988) );
	vdp_slatch g3129 (.Q(w4062), .D(S[4]), .C(w2958), .nC(w2985) );
	vdp_slatch g3130 (.Q(w4061), .D(S[4]), .C(w2960), .nC(w2983) );
	vdp_slatch g3131 (.Q(w4124), .D(S[3]), .C(w2952), .nC(w2976) );
	vdp_slatch g3132 (.Q(w4123), .D(S[3]), .C(w2956), .nC(w2981) );
	vdp_slatch g3133 (.Q(w4128), .D(S[3]), .C(w2957), .nC(w2982) );
	vdp_slatch g3134 (.Q(w4127), .D(S[3]), .C(w2959), .nC(w2977) );
	vdp_slatch g3135 (.Q(w4132), .D(S[7]), .C(w2952), .nC(w2976) );
	vdp_slatch g3136 (.Q(w4131), .D(S[7]), .C(w2956), .nC(w2981) );
	vdp_slatch g3137 (.Q(w4136), .D(S[7]), .C(w2957), .nC(w2982) );
	vdp_slatch g3138 (.Q(w4135), .D(S[7]), .C(w2959), .nC(w2977) );
	vdp_slatch g3139 (.Q(w4140), .D(S[2]), .C(w2952), .nC(w2976) );
	vdp_slatch g3140 (.Q(w4139), .D(S[2]), .C(w2956), .nC(w2981) );
	vdp_slatch g3141 (.Q(w4144), .D(S[2]), .C(w2957), .nC(w2982) );
	vdp_slatch g3142 (.Q(w4143), .D(S[2]), .C(w2959), .nC(w2977) );
	vdp_slatch g3143 (.Q(w4146), .D(S[6]), .C(w2952), .nC(w2976) );
	vdp_slatch g3144 (.Q(w4147), .D(S[6]), .C(w2956), .nC(w2981) );
	vdp_slatch g3145 (.Q(w4183), .D(S[6]), .C(w2957), .nC(w2982) );
	vdp_slatch g3146 (.Q(w4182), .D(S[6]), .C(w2959), .nC(w2977) );
	vdp_slatch g3147 (.Q(w4179), .D(S[1]), .C(w2952), .nC(w2976) );
	vdp_slatch g3148 (.Q(w4178), .D(S[1]), .C(w2956), .nC(w2981) );
	vdp_slatch g3149 (.Q(w4175), .D(S[1]), .C(w2957), .nC(w2982) );
	vdp_slatch g3150 (.Q(w4174), .D(S[1]), .C(w2959), .nC(w2977) );
	vdp_slatch g3151 (.Q(w4171), .D(S[5]), .C(w2952), .nC(w2976) );
	vdp_slatch g3152 (.Q(w4170), .D(S[5]), .C(w2956), .nC(w2981) );
	vdp_slatch g3153 (.Q(w4167), .D(S[5]), .C(w2957), .nC(w2982) );
	vdp_slatch g3154 (.Q(w4166), .D(S[5]), .C(w2959), .nC(w2977) );
	vdp_slatch g3155 (.Q(w4163), .D(S[0]), .C(w2952), .nC(w2976) );
	vdp_slatch g3156 (.Q(w4162), .D(S[0]), .C(w2956), .nC(w2981) );
	vdp_slatch g3157 (.Q(w4159), .D(S[0]), .C(w2957), .nC(w2982) );
	vdp_slatch g3158 (.Q(w4158), .D(S[0]), .C(w2959), .nC(w2977) );
	vdp_slatch g3159 (.Q(w4155), .D(S[4]), .C(w2952), .nC(w2976) );
	vdp_slatch g3160 (.Q(w4154), .D(S[4]), .C(w2956), .nC(w2981) );
	vdp_slatch g3161 (.Q(w4151), .D(S[4]), .C(w2957), .nC(w2982) );
	vdp_slatch g3162 (.Q(w4150), .D(S[4]), .C(w2959), .nC(w2977) );
	vdp_slatch g3163 (.Q(w4122), .D(w4124), .C(w2939), .nC(w2978) );
	vdp_slatch g3164 (.Q(w4121), .D(w4123), .C(w2942), .nC(w2979) );
	vdp_slatch g3165 (.Q(w4126), .D(w4128), .C(w2947), .nC(w2980) );
	vdp_slatch g3166 (.Q(w4125), .D(w4127), .C(w2944), .nC(w2949) );
	vdp_slatch g3167 (.Q(w4130), .D(w4132), .C(w2939), .nC(w2978) );
	vdp_slatch g3168 (.Q(w4129), .D(w4131), .C(w2942), .nC(w2979) );
	vdp_slatch g3169 (.Q(w4134), .D(w4136), .C(w2947), .nC(w2980) );
	vdp_slatch g3170 (.Q(w4133), .D(w4135), .C(w2944), .nC(w2949) );
	vdp_slatch g3171 (.Q(w4138), .D(w4140), .C(w2939), .nC(w2978) );
	vdp_slatch g3172 (.Q(w4137), .D(w4139), .C(w2942), .nC(w2979) );
	vdp_slatch g3173 (.Q(w4248), .D(w4144), .C(w2947), .nC(w2980) );
	vdp_slatch g3174 (.Q(w4142), .D(w4143), .C(w2944), .nC(w2949) );
	vdp_slatch g3175 (.Q(w4141), .D(w4146), .C(w2939), .nC(w2978) );
	vdp_slatch g3176 (.Q(w4145), .D(w4147), .C(w2942), .nC(w2979) );
	vdp_slatch g3177 (.Q(w4181), .D(w4183), .C(w2947), .nC(w2980) );
	vdp_slatch g3178 (.Q(w4180), .D(w4182), .C(w2944), .nC(w2949) );
	vdp_slatch g3179 (.Q(w4177), .D(w4179), .C(w2939), .nC(w2978) );
	vdp_slatch g3180 (.Q(w4176), .D(w4178), .C(w2942), .nC(w2979) );
	vdp_slatch g3181 (.Q(w4173), .D(w4175), .C(w2947), .nC(w2980) );
	vdp_slatch g3182 (.Q(w4172), .D(w4174), .C(w2944), .nC(w2949) );
	vdp_slatch g3183 (.Q(w4169), .D(w4171), .C(w2939), .nC(w2978) );
	vdp_slatch g3184 (.Q(w4168), .D(w4170), .C(w2942), .nC(w2979) );
	vdp_slatch g3185 (.Q(w4165), .D(w4167), .C(w2947), .nC(w2980) );
	vdp_slatch g3186 (.Q(w4164), .D(w4166), .C(w2944), .nC(w2949) );
	vdp_slatch g3187 (.D(w4163), .Q(w4161), .C(w2939), .nC(w2978) );
	vdp_slatch g3188 (.Q(w4160), .D(w4162), .C(w2942), .nC(w2979) );
	vdp_slatch g3189 (.Q(w4157), .D(w4159), .C(w2947), .nC(w2980) );
	vdp_slatch g3190 (.Q(w4156), .D(w4158), .C(w2944), .nC(w2949) );
	vdp_slatch g3191 (.Q(w4153), .D(w4155), .C(w2939), .nC(w2978) );
	vdp_slatch g3192 (.Q(w4152), .D(w4154), .C(w2942), .nC(w2979) );
	vdp_slatch g3193 (.Q(w4149), .D(w4151), .C(w2947), .nC(w2980) );
	vdp_slatch g3194 (.Q(w4148), .D(w4150), .C(w2944), .nC(w2949) );
	vdp_slatch g3195 (.Q(w3259), .D(w4122), .C(w2940), .nC(w2941) );
	vdp_slatch g3196 (.Q(w3258), .D(w4121), .C(w2948), .nC(w2943) );
	vdp_slatch g3197 (.Q(w3246), .D(w4126), .C(w2945), .nC(w2946) );
	vdp_slatch g3198 (.Q(w3244), .D(w4125), .C(w2938), .nC(w2937) );
	vdp_slatch g3199 (.Q(w3257), .D(w4130), .C(w2940), .nC(w2941) );
	vdp_slatch g3200 (.Q(w3256), .D(w4129), .C(w2948), .nC(w2943) );
	vdp_slatch g3201 (.D(w4134), .C(w2945), .nC(w2946), .Q(w3255) );
	vdp_slatch g3202 (.Q(w3243), .D(w4133), .C(w2938), .nC(w2937) );
	vdp_slatch g3203 (.Q(w3254), .D(w4138), .C(w2940), .nC(w2941) );
	vdp_slatch g3204 (.Q(w3253), .D(w4137), .C(w2948), .nC(w2943) );
	vdp_slatch g3205 (.Q(w3252), .D(w4248), .C(w2945), .nC(w2946) );
	vdp_slatch g3206 (.Q(w3251), .D(w4142), .C(w2938), .nC(w2937) );
	vdp_slatch g3207 (.Q(w3250), .D(w4141), .C(w2940), .nC(w2941) );
	vdp_slatch g3208 (.Q(w3249), .D(w4145), .C(w2948), .nC(w2943) );
	vdp_slatch g3209 (.Q(w3248), .D(w4181), .C(w2945), .nC(w2946) );
	vdp_slatch g3210 (.Q(w3247), .D(w4180), .C(w2938), .nC(w2937) );
	vdp_slatch g3211 (.Q(w3239), .D(w4177), .C(w2940), .nC(w2941) );
	vdp_slatch g3212 (.Q(w3285), .D(w4176), .C(w2948), .nC(w2943) );
	vdp_slatch g3213 (.Q(w3240), .D(w4173), .C(w2945), .nC(w2946) );
	vdp_slatch g3214 (.Q(w3241), .D(w4172), .C(w2938), .nC(w2937) );
	vdp_slatch g3215 (.Q(w3289), .D(w4169), .C(w2940), .nC(w2941) );
	vdp_slatch g3216 (.Q(w3298), .D(w4168), .C(w2948), .nC(w2943) );
	vdp_slatch g3217 (.Q(w3290), .D(w4165), .C(w2945), .nC(w2946) );
	vdp_slatch g3218 (.Q(w3297), .D(w4164), .nC(w2937), .C(w2938) );
	vdp_slatch g3219 (.Q(w3296), .D(w4161), .C(w2940), .nC(w2941) );
	vdp_slatch g3220 (.Q(w3295), .D(w4160), .C(w2948), .nC(w2943) );
	vdp_slatch g3221 (.Q(w3291), .D(w4157), .C(w2945), .nC(w2946) );
	vdp_slatch g3222 (.Q(w3294), .D(w4156), .C(w2938), .nC(w2937) );
	vdp_slatch g3223 (.Q(w3293), .D(w4153), .C(w2940), .nC(w2941) );
	vdp_slatch g3224 (.Q(w3292), .D(w4152), .C(w2948), .nC(w2943) );
	vdp_slatch g3225 (.Q(w3245), .D(w4149), .C(w2945), .nC(w2946) );
	vdp_slatch g3226 (.Q(w3242), .D(w4148), .C(w2938), .nC(w2937) );
	vdp_slatch g3227 (.Q(w3277), .D(w4187), .nC(w3336), .C(w3335) );
	vdp_slatch g3228 (.Q(w3384), .D(w4186), .nC(w3339), .C(w3340) );
	vdp_slatch g3229 (.Q(w3279), .D(w4191), .nC(w3338), .C(w3337) );
	vdp_slatch g3230 (.Q(w3278), .D(w4190), .nC(w3342), .C(w3341) );
	vdp_slatch g3231 (.Q(w3383), .D(w4195), .nC(w3336), .C(w3335) );
	vdp_slatch g3232 (.Q(w3387), .D(w4194), .nC(w3339), .C(w3340) );
	vdp_slatch g3233 (.Q(w3386), .D(w4199), .nC(w3338), .C(w3337) );
	vdp_slatch g3234 (.Q(w3385), .D(w4198), .nC(w3342), .C(w3341) );
	vdp_slatch g3235 (.Q(w3280), .D(w4203), .nC(w3336), .C(w3335) );
	vdp_slatch g3236 (.Q(w3388), .D(w4202), .nC(w3339), .C(w3340) );
	vdp_slatch g3237 (.Q(w3382), .D(w4207), .nC(w3338), .C(w3337) );
	vdp_slatch g3238 (.Q(w3389), .D(w4206), .nC(w3342), .C(w3341) );
	vdp_slatch g3239 (.Q(w3390), .D(w4211), .nC(w3336), .C(w3335) );
	vdp_slatch g3240 (.Q(w3391), .D(w4210), .nC(w3339), .C(w3340) );
	vdp_slatch g3241 (.Q(w3281), .D(w4215), .nC(w3338), .C(w3337) );
	vdp_slatch g3242 (.Q(w3282), .D(w4214), .nC(w3342), .C(w3341) );
	vdp_slatch g3243 (.Q(w3374), .D(w4219), .nC(w3336), .C(w3335) );
	vdp_slatch g3244 (.Q(w3375), .D(w4218), .nC(w3339), .C(w3340) );
	vdp_slatch g3245 (.Q(w3376), .D(w4223), .nC(w3338), .C(w3337) );
	vdp_slatch g3246 (.Q(w3377), .D(w4222), .nC(w3342), .C(w3341) );
	vdp_slatch g3247 (.Q(w3378), .D(w4227), .nC(w3336), .C(w3335) );
	vdp_slatch g3248 (.Q(w3379), .D(w4226), .nC(w3339), .C(w3340) );
	vdp_slatch g3249 (.Q(w3380), .D(w4231), .nC(w3338), .C(w3337) );
	vdp_slatch g3250 (.Q(w3381), .D(w4230), .nC(w3342), .C(w3341) );
	vdp_slatch g3251 (.Q(w3373), .D(w4235), .nC(w3336), .C(w3335) );
	vdp_slatch g3252 (.Q(w3372), .D(w4234), .nC(w3339), .C(w3340) );
	vdp_slatch g3253 (.Q(w3371), .D(w4239), .nC(w3338), .C(w3337) );
	vdp_slatch g3254 (.Q(w3370), .D(w4238), .nC(w3342), .C(w3341) );
	vdp_slatch g3255 (.Q(w3369), .D(w4243), .nC(w3336), .C(w3335) );
	vdp_slatch g3256 (.Q(w3368), .D(w4242), .nC(w3339), .C(w3340) );
	vdp_slatch g3257 (.Q(w3366), .D(w4247), .nC(w3338), .C(w3337) );
	vdp_slatch g3258 (.Q(w3367), .D(w4246), .nC(w3342), .C(w3341) );
	vdp_slatch g3259 (.Q(w4187), .D(w4185), .C(w3303), .nC(w3334) );
	vdp_slatch g3260 (.Q(w4186), .D(w4184), .C(w3326), .nC(w3328) );
	vdp_slatch g3261 (.Q(w4191), .D(w4189), .C(w3304), .nC(w3329) );
	vdp_slatch g3262 (.Q(w4190), .D(w4188), .C(w3333), .nC(w3332) );
	vdp_slatch g3263 (.Q(w4195), .D(w4193), .C(w3303), .nC(w3334) );
	vdp_slatch g3264 (.Q(w4194), .D(w4192), .C(w3326), .nC(w3328) );
	vdp_slatch g3265 (.Q(w4199), .D(w4197), .C(w3304), .nC(w3329) );
	vdp_slatch g3266 (.Q(w4198), .D(w4196), .C(w3333), .nC(w3332) );
	vdp_slatch g3267 (.Q(w4203), .D(w4201), .C(w3303), .nC(w3334) );
	vdp_slatch g3268 (.Q(w4202), .D(w4200), .C(w3326), .nC(w3328) );
	vdp_slatch g3269 (.Q(w4207), .D(w4205), .C(w3304), .nC(w3329) );
	vdp_slatch g3270 (.Q(w4206), .D(w4204), .C(w3333), .nC(w3332) );
	vdp_slatch g3271 (.Q(w4211), .D(w4209), .C(w3303), .nC(w3334) );
	vdp_slatch g3272 (.Q(w4210), .D(w4208), .C(w3326), .nC(w3328) );
	vdp_slatch g3273 (.Q(w4215), .D(w4213), .C(w3304), .nC(w3329) );
	vdp_slatch g3274 (.Q(w4214), .D(w4212), .C(w3333), .nC(w3332) );
	vdp_slatch g3275 (.Q(w4219), .D(w4217), .C(w3303), .nC(w3334) );
	vdp_slatch g3276 (.Q(w4218), .D(w4216), .C(w3326), .nC(w3328) );
	vdp_slatch g3277 (.Q(w4223), .D(w4221), .C(w3304), .nC(w3329) );
	vdp_slatch g3278 (.Q(w4222), .D(w4220), .C(w3333), .nC(w3332) );
	vdp_slatch g3279 (.Q(w4227), .D(w4225), .C(w3303), .nC(w3334) );
	vdp_slatch g3280 (.Q(w4226), .D(w4224), .C(w3326), .nC(w3328) );
	vdp_slatch g3281 (.Q(w4231), .D(w4229), .C(w3304), .nC(w3329) );
	vdp_slatch g3282 (.Q(w4230), .D(w4228), .C(w3333), .nC(w3332) );
	vdp_slatch g3283 (.Q(w4235), .D(w4233), .C(w3303), .nC(w3334) );
	vdp_slatch g3284 (.Q(w4234), .D(w4232), .C(w3326), .nC(w3328) );
	vdp_slatch g3285 (.Q(w4239), .D(w4237), .C(w3304), .nC(w3329) );
	vdp_slatch g3286 (.Q(w4238), .D(w4236), .C(w3333), .nC(w3332) );
	vdp_slatch g3287 (.Q(w4243), .D(w4241), .C(w3303), .nC(w3334) );
	vdp_slatch g3288 (.Q(w4242), .D(w4240), .C(w3326), .nC(w3328) );
	vdp_slatch g3289 (.Q(w4247), .D(w4245), .C(w3304), .nC(w3329) );
	vdp_slatch g3290 (.Q(w4246), .D(w4244), .C(w3333), .nC(w3332) );
	vdp_slatch g3291 (.Q(w4185), .D(S[3]), .nC(w3327), .C(w3356) );
	vdp_slatch g3292 (.Q(w4184), .D(S[3]), .nC(w3343), .C(w3357) );
	vdp_slatch g3293 (.Q(w4189), .D(S[3]), .nC(w3330), .C(w3355) );
	vdp_slatch g3294 (.Q(w4188), .D(S[3]), .nC(w3331), .C(w3354) );
	vdp_slatch g3295 (.Q(w4193), .D(S[7]), .nC(w3327), .C(w3356) );
	vdp_slatch g3296 (.Q(w4192), .D(S[7]), .nC(w3343), .C(w3357) );
	vdp_slatch g3297 (.Q(w4197), .D(S[7]), .nC(w3330), .C(w3355) );
	vdp_slatch g3298 (.Q(w4196), .D(S[7]), .nC(w3331), .C(w3354) );
	vdp_slatch g3299 (.Q(w4201), .D(S[2]), .nC(w3327), .C(w3356) );
	vdp_slatch g3300 (.Q(w4200), .D(S[2]), .nC(w3343), .C(w3357) );
	vdp_slatch g3301 (.Q(w4205), .D(S[2]), .nC(w3330), .C(w3355) );
	vdp_slatch g3302 (.Q(w4204), .D(S[2]), .nC(w3331), .C(w3354) );
	vdp_slatch g3303 (.Q(w4209), .D(S[6]), .nC(w3327), .C(w3356) );
	vdp_slatch g3304 (.Q(w4208), .D(S[6]), .nC(w3343), .C(w3357) );
	vdp_slatch g3305 (.Q(w4213), .D(S[6]), .nC(w3330), .C(w3355) );
	vdp_slatch g3306 (.Q(w4212), .D(S[6]), .nC(w3331), .C(w3354) );
	vdp_slatch g3307 (.Q(w4217), .D(S[1]), .nC(w3327), .C(w3356) );
	vdp_slatch g3308 (.Q(w4216), .D(S[1]), .nC(w3343), .C(w3357) );
	vdp_slatch g3309 (.Q(w4221), .D(S[1]), .nC(w3330), .C(w3355) );
	vdp_slatch g3310 (.Q(w4220), .D(S[1]), .nC(w3331), .C(w3354) );
	vdp_slatch g3311 (.Q(w4225), .D(S[5]), .nC(w3327), .C(w3356) );
	vdp_slatch g3312 (.Q(w4224), .D(S[5]), .nC(w3343), .C(w3357) );
	vdp_slatch g3313 (.Q(w4229), .D(S[5]), .nC(w3330), .C(w3355) );
	vdp_slatch g3314 (.Q(w4228), .D(S[5]), .nC(w3331), .C(w3354) );
	vdp_slatch g3315 (.Q(w4233), .D(S[0]), .nC(w3327), .C(w3356) );
	vdp_slatch g3316 (.Q(w4232), .D(S[0]), .nC(w3343), .C(w3357) );
	vdp_slatch g3317 (.Q(w4237), .D(S[0]), .nC(w3330), .C(w3355) );
	vdp_slatch g3318 (.Q(w4236), .D(S[0]), .nC(w3331), .C(w3354) );
	vdp_slatch g3319 (.Q(w4241), .D(S[4]), .nC(w3327), .C(w3356) );
	vdp_slatch g3320 (.Q(w4240), .D(S[4]), .nC(w3343), .C(w3357) );
	vdp_slatch g3321 (.Q(w4245), .D(S[4]), .nC(w3330), .C(w3355) );
	vdp_slatch g3322 (.Q(w4244), .D(S[4]), .nC(w3331), .C(w3354) );
	vdp_aon2x8 g3323 (.Z(w3884), .A1(w3076), .B1(w3075), .C1(w3074), .D2(w3073), .A2(w3120), .B2(w3121), .C2(w3126), .D1(w3125), .E2(w3123), .F1(w3124), .E1(w3072), .F2(w3071), .G1(w3070), .H2(w3069), .G2(w3128), .H1(w3118) );
	vdp_aon2x8 g3324 (.Z(w3100), .A1(w3193), .B1(w3121), .C1(w3195), .D2(w3125), .A2(w3120), .B2(w3194), .C2(w3126), .D1(w3196), .E2(w3123), .F1(w3124), .E1(w3197), .F2(w3198), .G1(w3204), .H2(w3205), .G2(w3128), .H1(w3118) );
	vdp_aon2x8 g3325 (.Z(w3103), .A1(w3068), .B1(w3081), .C1(w3085), .D2(w3084), .A2(w3120), .B2(w3121), .C2(w3126), .D1(w3125), .E2(w3123), .F1(w3124), .E1(w3083), .F2(w3079), .G1(w3080), .H2(w3082), .G2(w3128), .H1(w3118) );
	vdp_aon2x8 g3326 (.Z(w3104), .A1(w3206), .B1(w3121), .C1(w3208), .D2(w3125), .A2(w3120), .B2(w3207), .C2(w3126), .D1(w3203), .E2(w3123), .F1(w3124), .E1(w3209), .F2(w3210), .G1(w3211), .H2(w3212), .G2(w3128), .H1(w3118) );
	vdp_aon2x8 g3327 (.Z(w3102), .A1(w3138), .B1(w3121), .C1(w3140), .D2(w3141), .A2(w3120), .B2(w3885), .C2(w3126), .D1(w3125), .E2(w3123), .F1(w3124), .E1(w3213), .F2(w3139), .G1(w3119), .H2(w3142), .G2(w3128), .H1(w3118) );
	vdp_aon2x8 g3328 (.Z(w3105), .A1(w3145), .B1(w3121), .C1(w3152), .D2(w3151), .A2(w3120), .B2(w3153), .C2(w3126), .D1(w3125), .E2(w3123), .F1(w3124), .E1(w3149), .F2(w3143), .G1(w3150), .G2(w3128), .H1(w3118), .H2(w3144) );
	vdp_aon2x8 g3329 (.Z(w3101), .A1(w3086), .B1(w3087), .C1(w3089), .D2(w3088), .A2(w3120), .B2(w3121), .C2(w3126), .D1(w3125), .E2(w3123), .F1(w3124), .E1(w3130), .F2(w3131), .G1(w3127), .H2(w3122), .G2(w3128), .H1(w3118) );
	vdp_aon2x8 g3330 (.Z(w3106), .A1(w3134), .B1(w3133), .C1(w3132), .D2(w3129), .A2(w3120), .B2(w3121), .C2(w3126), .D1(w3125), .E2(w3123), .F1(w3124), .E1(w3115), .F2(w3114), .G1(w3116), .H2(w3117), .G2(w3128), .H1(w3118) );
	vdp_aon2x8 g3331 (.A1(w3259), .B1(w3258), .C1(w3246), .D2(w3244), .A2(w3276), .B2(w3275), .C2(w3274), .D1(w3273), .E2(w3272), .F1(w3271), .E1(w3257), .F2(w3256), .G1(w3255), .H2(w3243), .G2(w3269), .H1(w3270), .Z(w3288) );
	vdp_aon2x8 g3332 (.Z(w3314), .A1(w3254), .B1(w3253), .C1(w3252), .D2(w3251), .A2(w3276), .B2(w3275), .C2(w3274), .D1(w3273), .E2(w3272), .F1(w3271), .E1(w3250), .F2(w3249), .G1(w3248), .H2(w3247), .G2(w3269), .H1(w3270) );
	vdp_aon2x8 g3333 (.Z(w3287), .A1(w3246), .B1(w3255), .C1(w3252), .D2(w3248), .A2(w3271), .B2(w3270), .C2(w3275), .D1(w3273), .E2(w3272), .F1(w3269), .E1(w3240), .F2(w3290), .G1(w3291), .H2(w3245), .G2(w3276), .H1(w3274) );
	vdp_aon2x8 g3334 (.Z(w3317), .A1(w3239), .B1(w3285), .C1(w3240), .D2(w3241), .A2(w3276), .B2(w3275), .C2(w3274), .D1(w3273), .E2(w3272), .F1(w3271), .E1(w3289), .F2(w3298), .G1(w3290), .H2(w3297), .G2(w3269), .H1(w3270) );
	vdp_aon2x8 g3335 (.Z(w3286), .A1(w3296), .B1(w3295), .C1(w3291), .D2(w3294), .A2(w3276), .B2(w3275), .C2(w3274), .D1(w3273), .E2(w3272), .F1(w3271), .E1(w3293), .F2(w3292), .G1(w3245), .H2(w3242), .G2(w3269), .H1(w3270) );
	vdp_aon2x8 g3336 (.Z(w3319), .A1(w3373), .B1(w3275), .C1(w3371), .D2(w3273), .A2(w3276), .B2(w3372), .C2(w3274), .D1(w3370), .E2(w3272), .F1(w3271), .E1(w3369), .F2(w3368), .G1(w3366), .H2(w3367), .G2(w3269), .H1(w3270) );
	vdp_aon2x8 g3337 (.Z(w3320), .A1(w3374), .B1(w3275), .C1(w3376), .D2(w3273), .A2(w3276), .B2(w3375), .C2(w3274), .D1(w3377), .E2(w3272), .F1(w3271), .E1(w3378), .F2(w3379), .G1(w3380), .H2(w3381), .G2(w3269), .H1(w3270) );
	vdp_aon2x8 g3338 (.Z(w3318), .A1(w3244), .B1(w3243), .C1(w3251), .D2(w3247), .A2(w3271), .B2(w3270), .C2(w3275), .D1(w3273), .E2(w3272), .F1(w3269), .E1(w3241), .F2(w3297), .G1(w3294), .H2(w3242), .G2(w3276), .H1(w3274) );
	vdp_aon2x8 g3339 (.Z(w3313), .A1(w3278), .B1(w3270), .C1(w3389), .D2(w3273), .A2(w3271), .B2(w3385), .C2(w3275), .D1(w3282), .E2(w3272), .F1(w3269), .E1(w3377), .F2(w3381), .G1(w3370), .H2(w3367), .G2(w3276), .H1(w3274) );
	vdp_aon2x8 g3340 (.Z(w3316), .A1(w3279), .B1(w3270), .C1(w3382), .D2(w3273), .A2(w3271), .B2(w3386), .C2(w3275), .D1(w3281), .E2(w3272), .F1(w3269), .E1(w3376), .F2(w3380), .G1(w3371), .H2(w3366), .G2(w3276), .H1(w3274) );
	vdp_aon2x8 g3341 (.Z(w3315), .A1(w3280), .B1(w3275), .C1(w3382), .D2(w3273), .A2(w3276), .B2(w3388), .C2(w3274), .D1(w3389), .E2(w3272), .F1(w3271), .E1(w3390), .F2(w3391), .G1(w3281), .H2(w3282), .G2(w3269), .H1(w3270) );
	vdp_aon2x8 g3342 (.A1(w3277), .B1(w3275), .C1(w3279), .D2(w3273), .A2(w3276), .B2(w3384), .C2(w3274), .D1(w3278), .E2(w3272), .F1(w3271), .E1(w3383), .F2(w3387), .G1(w3386), .H2(w3385), .G2(w3269), .H1(w3270), .Z(w3321) );
	vdp_sr_bit g3343 (.Q(w3266), .D(w3408), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3344 (.Q(w3408), .D(w3886), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3345 (.Q(w3324), .D(w3409), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3346 (.Q(w3409), .D(w3325), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3347 (.Q(w3323), .D(w3302), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3348 (.Q(w3913), .D(w3323), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3349 (.Q(w3392), .D(w3322), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3350 (.Q(w3301), .D(w3392), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3351 (.Q(w3915), .D(w3407), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3352 (.Q(w3300), .D(w3915), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3353 (.Q(w3299), .D(w3267), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3354 (.Q(w3267), .D(w3310), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3355 (.Q(w2727), .D(w3311), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3356 (.Q(w3393), .D(w2727), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3357 (.Q(w3092), .D(w3110), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3358 (.Q(w3094), .D(w3092), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3359 (.Q(w3097), .D(w3093), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3360 (.Q(w3093), .D(w3109), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3361 (.Q(w3108), .D(w3090), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3362 (.Q(w3090), .D(w3111), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3363 (.Q(w3091), .D(w3107), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3364 (.Q(w3099), .D(w3091), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3365 (.Q(w3176), .D(w2726), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3366 (.Q(w2726), .D(w3175), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3367 (.Q(w3896), .D(w3112), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3368 (.Q(w3098), .D(w3896), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3369 (.Q(w3895), .D(w3174), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3370 (.Q(w3096), .D(w3895), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3371 (.Q(w3024), .D(VRAMA[1]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3372 (.Q(w3056), .D(VRAMA[2]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3373 (.Q(w3058), .D(VRAMA[3]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3374 (.Q(w3059), .D(VRAMA[4]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3375 (.Q(w3060), .D(VRAMA[5]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3376 (.Q(w3061), .D(VRAMA[6]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3377 (.Q(w3893), .D(w3047), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3378 (.Q(w3394), .D(w3893), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3379 (.Q(w3046), .D(w3395), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3380 (.Q(w3395), .D(w3394), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_dlatch_inv g3381 (.nQ(w3047), .D(w3011), .C(DCLK1), .nC(nDCLK1) );
	vdp_slatch g3382 (.Q(w3168), .D(w4249), .C(w3162), .nC(w2925) );
	vdp_slatch g3383 (.Q(w4286), .D(w4250), .C(w3162), .nC(w2925) );
	vdp_slatch g3384 (.Q(w3167), .D(w4251), .C(w3162), .nC(w2925) );
	vdp_slatch g3385 (.Q(w3166), .D(w4252), .C(w3162), .nC(w2925) );
	vdp_slatch g3386 (.Q(w3165), .D(w4253), .C(w3162), .nC(w2925) );
	vdp_slatch g3387 (.Q(w3164), .D(w4254), .C(w3162), .nC(w2925) );
	vdp_slatch g3388 (.Q(w3163), .D(w4256), .C(w3162), .nC(w2925) );
	vdp_slatch g3389 (.Q(w2926), .D(w4255), .C(w3162), .nC(w2925) );
	vdp_slatch g3390 (.Q(w4249), .D(w2992), .C(w3183), .nC(w3215) );
	vdp_slatch g3391 (.Q(w4250), .D(w2967), .C(w3183), .nC(w3215) );
	vdp_slatch g3392 (.Q(w4251), .D(w2969), .C(w3183), .nC(w3215) );
	vdp_slatch g3393 (.Q(w4252), .D(w2970), .C(w3183), .nC(w3215) );
	vdp_slatch g3394 (.Q(w4253), .D(w2971), .C(w3183), .nC(w3215) );
	vdp_slatch g3395 (.Q(w4254), .D(w2993), .C(w3183), .nC(w3215) );
	vdp_slatch g3396 (.Q(w4256), .D(w2997), .C(w3183), .nC(w3215) );
	vdp_slatch g3397 (.Q(w4255), .D(w2996), .C(w3183), .nC(w3215) );
	vdp_slatch g3398 (.Q(w4257), .D(w2933), .C(w2935), .nC(w2934) );
	vdp_slatch g3399 (.Q(w4258), .D(w2966), .C(w2935), .nC(w2934) );
	vdp_slatch g3400 (.Q(w4259), .D(w2932), .C(w2935), .nC(w2934) );
	vdp_slatch g3401 (.Q(w4260), .D(w3947), .C(w2935), .nC(w2934) );
	vdp_slatch g3402 (.Q(w4261), .D(w3403), .C(w2935), .nC(w2934) );
	vdp_slatch g3403 (.Q(w4262), .D(w2973), .C(w2935), .nC(w2934) );
	vdp_slatch g3404 (.Q(w4263), .D(w2929), .C(w2935), .nC(w2934) );
	vdp_slatch g3405 (.Q(w4264), .D(w2974), .C(w2935), .nC(w2934) );
	vdp_slatch g3406 (.Q(w3224), .D(w4257), .C(w2936), .nC(w3217) );
	vdp_slatch g3407 (.Q(w3223), .D(w4258), .C(w2936), .nC(w3217) );
	vdp_slatch g3408 (.Q(w3222), .D(w4259), .C(w2936), .nC(w3217) );
	vdp_slatch g3409 (.Q(w3221), .D(w4260), .C(w2936), .nC(w3217) );
	vdp_slatch g3410 (.Q(w3220), .D(w4261), .C(w2936), .nC(w3217) );
	vdp_slatch g3411 (.Q(w3219), .D(w4262), .C(w2936), .nC(w3217) );
	vdp_slatch g3412 (.Q(w3218), .D(w4263), .C(w2936), .nC(w3217) );
	vdp_slatch g3413 (.Q(w4287), .D(w4264), .C(w2936), .nC(w3217) );
	vdp_slatch g3414 (.Q(w3358), .D(w3352), .C(w3044), .nC(w3348) );
	vdp_slatch g3415 (.Q(w3350), .D(w3051), .C(w3044), .nC(w3348) );
	vdp_slatch g3416 (.Q(w3732), .D(w3349), .C(w3044), .nC(w3348) );
	vdp_slatch g3417 (.Q(w3344), .D(w3347), .C(w3044), .nC(w3348) );
	vdp_slatch g3418 (.Q(w2933), .D(w2992), .C(w2995), .nC(w2994) );
	vdp_slatch g3419 (.Q(w2966), .D(w2967), .C(w2995), .nC(w2994) );
	vdp_slatch g3420 (.Q(w2932), .D(w2969), .C(w2995), .nC(w2994) );
	vdp_slatch g3421 (.Q(w3947), .D(w2970), .C(w2995), .nC(w2994) );
	vdp_slatch g3422 (.Q(w3403), .D(w2971), .C(w2995), .nC(w2994) );
	vdp_slatch g3423 (.Q(w2973), .D(w2993), .C(w2995), .nC(w2994) );
	vdp_slatch g3424 (.Q(w2929), .D(w2997), .C(w2995), .nC(w2994) );
	vdp_slatch g3425 (.Q(w2974), .D(w2996), .C(w2995), .nC(w2994) );
	vdp_cnt_bit_load g3426 (.D(w3349), .nL(w3015), .L(w3012), .R(1'b0), .Q(w3014), .CI(w3399), .CO(w3400), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3427 (.D(w3051), .nL(w3015), .L(w3012), .R(1'b0), .Q(w3883), .CI(w3400), .CO(w3401), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3428 (.D(w3016), .nL(w3015), .L(w3012), .R(1'b0), .Q(w3000), .CI(w3401), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3429 (.CO(w3399), .CI(1'b1), .D(w3347), .nL(w3015), .L(w3012), .R(1'b0), .Q(w3010), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3430 (.CO(w3398), .CI(1'b1), .D(w3344), .nL(w3346), .L(w3043), .R(1'b0), .Q(w3365), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3431 (.CO(w3397), .CI(w3398), .D(w3732), .nL(w3346), .L(w3043), .R(1'b0), .Q(w3312), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3432 (.CO(w3396), .CI(w3397), .D(w3350), .nL(w3346), .L(w3043), .R(1'b0), .Q(w3353), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3433 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .CI(w3396), .D(w3358), .nL(w3346), .L(w3043), .R(1'b0), .Q(w3265) );
	vdp_xor g3434 (.Z(w3154), .B(w3883), .A(w3009) );
	vdp_xor g3435 (.B(w3014), .A(w3009), .Z(w3001) );
	vdp_xor g3436 (.Z(w3157), .B(w3010), .A(w3009) );
	vdp_sr_bit g3437 (.Q(w3008), .D(w3891), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3438 (.Q(w3890), .D(w3008), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3439 (.Q(w3173), .D(w3890), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3440 (.Q(w3899), .D(w3402), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3441 (.Q(w3402), .D(w3900), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3442 (.Q(w3900), .D(w3901), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3443 (.Q(w2931), .D(w2930), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3444 (.Q(w2930), .D(w2928), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3445 (.Q(w2928), .D(w2927), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3446 (.Q(w3903), .D(w3904), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3447 (.Q(w3871), .D(w3903), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3448 (.Q(w3902), .D(w3871), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3449 (.Q(w3907), .D(w3906), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3450 (.Q(w3908), .D(w3907), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3451 (.Q(w3905), .D(w3908), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3452 (.Q(w3022), .D(w3905), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3453 (.Q(w3989), .D(w3990), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3454 (.Q(w3990), .D(w3909), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_xor g3455 (.Z(w3227), .A(w3309), .B(w3353) );
	vdp_xor g3456 (.Z(w3232), .A(w3309), .B(w3364) );
	vdp_xor g3457 (.Z(w3226), .A(w3309), .B(w3365) );
	vdp_dlatch_inv g3458 (.nQ(w3889), .D(w3888), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g3459 (.nQ(w2927), .D(w2972), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g3460 (.nQ(w3904), .D(w2923), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g3461 (.nQ(w3363), .D(w3910), .nC(nHCLK1), .C(HCLK1) );
	vdp_xor g3462 (.Z(w3364), .A(w3312), .B(M5) );
	vdp_sr_bit g3463 (.Q(w3405), .D(w3351), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_dlatch_inv g3464 (.nQ(w3906), .D(w3020), .nC(nDCLK1), .C(DCLK1) );
	vdp_comp_strong g3465 (.Z(w2940), .nZ(w2941), .A(w3216) );
	vdp_comp_strong g3466 (.Z(w2948), .nZ(w2943), .A(w3216) );
	vdp_comp_strong g3467 (.Z(w2945), .nZ(w2946), .A(w3216) );
	vdp_comp_strong g3468 (.Z(w2938), .nZ(w2937), .A(w3216) );
	vdp_comp_strong g3469 (.Z(w2939), .nZ(w2978), .A(w3023) );
	vdp_comp_strong g3470 (.Z(w2942), .nZ(w2979), .A(w3023) );
	vdp_comp_strong g3471 (.Z(w2947), .nZ(w2980), .A(w3023) );
	vdp_comp_strong g3472 (.Z(w2944), .nZ(w2949), .A(w3023) );
	vdp_comp_strong g3473 (.Z(w2952), .nZ(w2976), .A(w2975) );
	vdp_comp_strong g3474 (.Z(w2956), .nZ(w2981), .A(w3284) );
	vdp_comp_strong g3475 (.Z(w2957), .nZ(w2982), .A(w3283) );
	vdp_comp_strong g3476 (.Z(w2959), .nZ(w2977), .A(w2968) );
	vdp_comp_strong g3477 (.Z(w2951), .nZ(w2984), .A(w3898) );
	vdp_comp_strong g3478 (.Z(w2955), .nZ(w2988), .A(w2989) );
	vdp_comp_strong g3479 (.Z(w2958), .nZ(w2985), .A(w2991) );
	vdp_comp_strong g3480 (.Z(w2960), .nZ(w2983), .A(w2990) );
	vdp_comp_strong g3481 (.Z(w3190), .nZ(w3177), .A(w2924) );
	vdp_comp_strong g3482 (.Z(w2998), .nZ(w3178), .A(w2924) );
	vdp_comp_strong g3483 (.Z(w3184), .nZ(w2986), .A(w2924) );
	vdp_comp_strong g3484 (.Z(w3185), .nZ(w2987), .A(w2924) );
	vdp_comp_strong g3485 (.Z(w3189), .nZ(w3191), .A(w2999) );
	vdp_comp_strong g3486 (.Z(w3188), .nZ(w3199), .A(w2999) );
	vdp_comp_strong g3487 (.Z(w3187), .nZ(w3200), .A(w2999) );
	vdp_comp_strong g3488 (.Z(w3186), .nZ(w3192), .A(w2999) );
	vdp_comp_strong g3489 (.Z(w3041), .nZ(w3067), .A(w2999) );
	vdp_comp_strong g3490 (.Z(w3019), .nZ(w3077), .A(w2999) );
	vdp_comp_strong g3491 (.Z(w3032), .nZ(w3078), .A(w2999) );
	vdp_comp_strong g3492 (.Z(w3033), .nZ(w3006), .A(w2999) );
	vdp_comp_strong g3493 (.Z(w3018), .nZ(w3036), .A(w2924) );
	vdp_comp_strong g3494 (.Z(w3037), .nZ(w3028), .A(w2924) );
	vdp_comp_strong g3495 (.Z(w3038), .nZ(w3026), .A(w2924) );
	vdp_comp_strong g3496 (.Z(w3034), .nZ(w3035), .A(w2924) );
	vdp_comp_strong g3497 (.Z(w3049), .nZ(w3039), .A(w3050) );
	vdp_comp_strong g3498 (.Z(w3030), .nZ(w3029), .A(w3052) );
	vdp_comp_strong g3499 (.Z(w3031), .nZ(w3027), .A(w3053) );
	vdp_comp_strong g3500 (.Z(w3048), .nZ(w3040), .A(w3054) );
	vdp_comp_strong g3501 (.Z(w3356), .nZ(w3327), .A(w3171) );
	vdp_comp_strong g3502 (.Z(w3357), .nZ(w3343), .A(w3359) );
	vdp_comp_strong g3503 (.Z(w3355), .nZ(w3330), .A(w3360) );
	vdp_comp_strong g3504 (.Z(w3354), .nZ(w3331), .A(w3361) );
	vdp_comp_strong g3505 (.Z(w3303), .nZ(w3334), .A(w3023) );
	vdp_comp_strong g3506 (.Z(w3326), .nZ(w3328), .A(w3023) );
	vdp_comp_strong g3507 (.Z(w3304), .nZ(w3329), .A(w3023) );
	vdp_comp_strong g3508 (.Z(w3333), .nZ(w3332), .A(w3023) );
	vdp_comp_strong g3509 (.Z(w3335), .nZ(w3336), .A(w3216) );
	vdp_comp_strong g3510 (.Z(w3340), .nZ(w3339), .A(w3216) );
	vdp_comp_strong g3511 (.Z(w3337), .nZ(w3338), .A(w3216) );
	vdp_comp_strong g3512 (.Z(w3341), .nZ(w3342), .A(w3216) );
	vdp_not g3513 (.nZ(w3016), .A(w3352) );
	vdp_not g3514 (.nZ(w3891), .A(w3135) );
	vdp_not g3515 (.nZ(w3137), .A(w88) );
	vdp_not g3516 (.nZ(w3136), .A(w406) );
	vdp_not g3517 (.nZ(w3002), .A(w3136) );
	vdp_comp_strong g3518 (.Z(w3162), .nZ(w2925), .A(w2999) );
	vdp_comp_strong g3519 (.Z(w3183), .nZ(w3215), .A(w2924) );
	vdp_comp_strong g3520 (.Z(w2995), .nZ(w2994), .A(w3171) );
	vdp_comp_strong g3521 (.Z(w2936), .nZ(w3217), .A(w3216) );
	vdp_comp_strong g3522 (.Z(w2935), .nZ(w2934), .A(w3023) );
	vdp_comp_strong g3523 (.Z(w3044), .nZ(w3348), .A(w3405) );
	vdp_not g3524 (.nZ(w3233), .A(w3226) );
	vdp_not g3525 (.nZ(w3225), .A(w3232) );
	vdp_not g3526 (.nZ(w3236), .A(w3227) );
	vdp_nand3 g3527 (.Z(w3230), .A(w3236), .B(w3232), .C(w3226) );
	vdp_not g3528 (.nZ(w3275), .A(w3229) );
	vdp_nand3 g3529 (.Z(w3229), .A(w3227), .B(w3225), .C(w3226) );
	vdp_nand3 g3530 (.Z(w3228), .A(w3227), .B(w3232), .C(w3226) );
	vdp_nand3 g3531 (.Z(w3234), .A(w3227), .B(w3232), .C(w3233) );
	vdp_nand3 g3532 (.Z(w3231), .A(w3236), .B(w3225), .C(w3226) );
	vdp_nand3 g3533 (.Z(w3237), .A(w3236), .B(w3232), .C(w3233) );
	vdp_nand3 g3534 (.Z(w3235), .A(w3227), .B(w3225), .C(w3233) );
	vdp_nand3 g3535 (.Z(w3238), .A(w3233), .B(w3236), .C(w3225) );
	vdp_not g3536 (.nZ(w3276), .A(w3228) );
	vdp_not g3537 (.nZ(w3274), .A(w3230) );
	vdp_not g3538 (.nZ(w3273), .A(w3231) );
	vdp_not g3539 (.nZ(w3271), .A(w3235) );
	vdp_not g3540 (.nZ(w3272), .A(w3234) );
	vdp_not g3541 (.nZ(w3270), .A(w3238) );
	vdp_not g3542 (.nZ(w3269), .A(w3237) );
	vdp_not g3543 (.nZ(w3147), .A(w3157) );
	vdp_not g3544 (.nZ(w3155), .A(w3007) );
	vdp_not g3545 (.nZ(w3146), .A(w3154) );
	vdp_nand3 g3546 (.Z(w3159), .A(w3146), .B(w3007), .C(w3157) );
	vdp_not g3547 (.nZ(w3121), .A(w3161) );
	vdp_nand3 g3548 (.Z(w3161), .A(w3154), .B(w3155), .C(w3157) );
	vdp_nand3 g3549 (.Z(w3160), .A(w3154), .B(w3007), .C(w3157) );
	vdp_nand3 g3550 (.Z(w3897), .A(w3154), .B(w3007), .C(w3147) );
	vdp_nand3 g3551 (.Z(w3158), .A(w3146), .B(w3155), .C(w3157) );
	vdp_nand3 g3552 (.Z(w3156), .A(w3154), .B(w3155), .C(w3147) );
	vdp_not g3553 (.nZ(w3120), .A(w3160) );
	vdp_not g3554 (.nZ(w3126), .A(w3159) );
	vdp_not g3555 (.nZ(w3125), .A(w3158) );
	vdp_not g3556 (.nZ(w3124), .A(w3156) );
	vdp_not g3557 (.nZ(w3123), .A(w3897) );
	vdp_aon22 g3558 (.Z(w3175), .A1(w3163), .B1(w3169), .A2(w3170), .B2(w2926) );
	vdp_aon22 g3559 (.Z(w3174), .A1(w3165), .B1(w3169), .A2(w3170), .B2(w3164) );
	vdp_aon22 g3560 (.Z(w3112), .A1(w3167), .B1(w3169), .A2(w3170), .B2(w3166) );
	vdp_aon22 g3561 (.Z(w3009), .A1(w3168), .B1(w3169), .A2(w3170), .B2(w4286) );
	vdp_sr_bit g3562 (.Q(w3005), .D(w3892), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3563 (.Q(w3892), .D(w3004), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_xor g3564 (.Z(w3007), .A(w3001), .B(1'b1) );
	vdp_xor g3565 (.A(HPOS[3]), .B(w3025), .Z(w3946) );
	vdp_aon22 g3566 (.Z(w3063), .A1(w3056), .B1(w3057), .A2(w3055), .B2(w3945) );
	vdp_aon22 g3567 (.Z(w3064), .A1(w3058), .B1(w3057), .A2(w3055), .B2(w3944) );
	vdp_aon22 g3568 (.Z(w3066), .A1(w3059), .B1(w3057), .A2(w3055), .B2(w3943) );
	vdp_aon22 g3569 (.Z(w3065), .A1(w3060), .B1(w3057), .A2(w3055), .B2(w3942) );
	vdp_aon22 g3570 (.Z(w3486), .A1(w3061), .B1(w3057), .A2(w3055), .B2(w3941) );
	vdp_aon22 g3571 (.Z(w3107), .A1(w3202), .B1(w3884), .A2(w3100), .B2(w3201) );
	vdp_aon22 g3572 (.Z(w3111), .A1(w3202), .B1(w3101), .A2(w3102), .B2(w3201) );
	vdp_aon22 g3573 (.Z(w3109), .A1(w3202), .B1(w3106), .A2(w3105), .B2(w3201) );
	vdp_aon22 g3574 (.Z(w3110), .A1(w3202), .B1(w3103), .A2(w3104), .B2(w3201) );
	vdp_aon222 g3575 (.Z(w3886), .A1(w3315), .B1(w3314), .C1(w3313), .A2(w3263), .B2(w3264), .C2(w3262) );
	vdp_aon222 g3576 (.Z(w3325), .A1(w3319), .B1(w3286), .C1(w3318), .A2(w3263), .B2(w3264), .C2(w3262) );
	vdp_aon222 g3577 (.Z(w3302), .A1(w3320), .B1(w3317), .C1(w3287), .A2(w3263), .B2(w3264), .C2(w3262) );
	vdp_aon222 g3578 (.A1(w3321), .B1(w3288), .C1(w3316), .A2(w3263), .B2(w3264), .C2(w3262), .Z(w3322) );
	vdp_and5 g3579 (.Z(w3362), .A(w3351), .B(w3358), .C(w3350), .D(w3732), .E(w3344) );
	vdp_aon22 g3580 (.Z(w3407), .A1(w3220), .B1(w3406), .A2(w3042), .B2(w3219) );
	vdp_aon22 g3581 (.Z(w3310), .A1(w3222), .B1(w3406), .A2(w3042), .B2(w3221) );
	vdp_aon22 g3582 (.Z(w3309), .A1(w3224), .B1(w3406), .A2(w3042), .B2(w3223) );
	vdp_aon22 g3583 (.Z(w3311), .A1(w3218), .B1(w3406), .A2(w3042), .B2(w4287) );
	vdp_aon22 g3584 (.Z(w3021), .A1(w3306), .B1(w3046), .A2(w3022), .B2(M5) );
	vdp_and4 g3585 (.Z(w3307), .A(w3365), .B(w3312), .C(w3353), .D(w3308) );
	vdp_comp_we g3586 (.Z(w3042), .nZ(w3406), .A(w3305) );
	vdp_comp_we g3587 (.Z(w3201), .nZ(w3202), .A(w3000) );
	vdp_comp_we g3588 (.Z(w3170), .nZ(w3169), .A(w3000) );
	vdp_comp_we g3589 (.Z(w3012), .nZ(w3015), .A(w3095) );
	vdp_comp_we g3590 (.Z(w3055), .nZ(w3057), .A(w3573) );
	vdp_comp_we g3591 (.Z(w3043), .nZ(w3346), .A(w3351) );
	vdp_not g3592 (.nZ(w3911), .A(M5) );
	vdp_dlatch_inv g3593 (.nQ(w3901), .D(w3017), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g3594 (.Z(w3181), .A(DCLK2), .B(w2928) );
	vdp_and g3595 (.Z(w3182), .A(DCLK2), .B(w2927) );
	vdp_and g3596 (.Z(w3180), .A(DCLK2), .B(w2930) );
	vdp_and g3597 (.Z(w3179), .A(DCLK2), .B(w2931) );
	vdp_and g3598 (.Z(w2990), .A(w3901), .B(DCLK2) );
	vdp_and g3599 (.Z(w2991), .A(w3900), .B(DCLK2) );
	vdp_and g3600 (.Z(w2989), .A(w3402), .B(DCLK2) );
	vdp_and g3601 (.Z(w3898), .A(w3899), .B(DCLK2) );
	vdp_and g3602 (.Z(w2975), .A(DCLK2), .B(w3902) );
	vdp_and g3603 (.Z(w3284), .A(DCLK2), .B(w3871) );
	vdp_and g3604 (.Z(w3283), .A(DCLK2), .B(w3903) );
	vdp_and g3605 (.Z(w2968), .A(DCLK2), .B(w3904) );
	vdp_and g3606 (.Z(w2999), .A(w3889), .B(HCLK2) );
	vdp_and g3607 (.Z(w3172), .A(w3137), .B(w3008) );
	vdp_and g3608 (.Z(w3216), .A(w3363), .B(HCLK2) );
	vdp_or g3609 (.Z(w3308), .A(w3911), .B(w3265) );
	vdp_and g3610 (.Z(w3023), .A(w3021), .B(DCLK2) );
	vdp_and g3611 (.Z(w3361), .A(DCLK2), .B(w3906) );
	vdp_and g3612 (.Z(w3360), .A(DCLK2), .B(w3907) );
	vdp_and g3613 (.Z(w3359), .A(DCLK2), .B(w3908) );
	vdp_and g3614 (.Z(w3171), .A(DCLK2), .B(w3905) );
	vdp_and g3615 (.Z(w3305), .A(M5), .B(w3265) );
	vdp_and g3616 (.Z(w3942), .A(VSCR), .B(HPOS[7]) );
	vdp_and g3617 (.Z(w3941), .A(VSCR), .B(HPOS[8]) );
	vdp_and g3618 (.Z(w3054), .A(DCLK2), .B(w3047) );
	vdp_and g3619 (.Z(w3943), .A(VSCR), .B(HPOS[6]) );
	vdp_and g3620 (.Z(w3053), .A(DCLK2), .B(w3893) );
	vdp_and g3621 (.Z(w3052), .A(DCLK2), .B(w3394) );
	vdp_and g3622 (.Z(w3050), .A(DCLK2), .B(w3395) );
	vdp_and g3623 (.Z(w3944), .A(VSCR), .B(HPOS[5]) );
	vdp_and g3624 (.Z(w2924), .A(DCLK2), .B(w3046) );
	vdp_and g3625 (.Z(w3945), .A(VSCR), .B(HPOS[4]) );
	vdp_aon22 g3626 (.Z(w3062), .A1(w3024), .B1(w3057), .A2(w3055), .B2(w3946) );
	vdp_and g3627 (.nZ(w3025), .A(VSCR), .B(M5) );
	vdp_or4 g3628 (.Z(w2872), .D(w3090), .C(w3091), .B(w3092), .A(w3093) );
	vdp_or g3629 (.Z(w3095), .A(w77), .B(w14) );
	vdp_or g3630 (.Z(w3351), .A(w9), .B(w75) );
	vdp_or4 g3631 (.Z(w2873), .A(w3409), .B(w3408), .C(w3392), .D(w3323) );
	vdp_not g3632 (.nZ(w3909), .A(w3268) );
	vdp_not g3633 (.nZ(w3004), .A(w3113) );
	vdp_not g3634 (.nZ(w3306), .A(M5) );
	vdp_aoi21 g3635 (.Z(w3268), .A1(w90), .A2(w3002), .B(w16) );
	vdp_aoi21 g3636 (.Z(w3113), .A1(w91), .A2(w3002), .B(w10) );
	vdp_aoi21 g3637 (.Z(w3135), .A1(w88), .A2(w3002), .B(w11) );
	vdp_nand4 g3638 (.D(w3000), .C(w3010), .Z(w3888), .A(w3883), .B(w3014) );
	vdp_nand3 g3639 (.Z(w3148), .A(w3146), .B(w3007), .C(w3147) );
	vdp_not g3640 (.nZ(w3128), .A(w3148) );
	vdp_nand3 g3641 (.Z(w3214), .A(w3147), .B(w3146), .C(w3155) );
	vdp_not g3642 (.nZ(w3118), .A(w3214) );
	vdp_not g3643 (.nZ(w3264), .A(w3260) );
	vdp_not g3644 (.nZ(w3263), .A(w3261) );
	vdp_not g3645 (.nZ(w3887), .A(w3265) );
	vdp_not g3646 (.nZ(w3262), .A(M5) );
	vdp_not g3647 (.nZ(w3914), .A(PLANE_A_PRIO) );
	vdp_not g3648 (.nZ(w3894), .A(PLANE_B_PRIO) );
	vdp_bufif0 g3649 (.Z(COL[5]), .A(w3096), .nE(w3894) );
	vdp_bufif0 g3650 (.Z(COL[6]), .A(w3176), .nE(w3894) );
	vdp_bufif0 g3651 (.Z(COL[4]), .A(w3098), .nE(w3894) );
	vdp_bufif0 g3652 (.Z(COL[3]), .A(w3099), .nE(w3894) );
	vdp_bufif0 g3653 (.Z(COL[2]), .A(w3094), .nE(w3894) );
	vdp_bufif0 g3654 (.Z(COL[1]), .A(w3108), .nE(w3894) );
	vdp_bufif0 g3655 (.Z(COL[0]), .A(w3097), .nE(w3894) );
	vdp_bufif0 g3656 (.Z(COL[5]), .A(w3300), .nE(w3914) );
	vdp_bufif0 g3657 (.Z(COL[6]), .A(w3393), .nE(w3914) );
	vdp_bufif0 g3658 (.Z(COL[4]), .A(w3299), .nE(w3914) );
	vdp_bufif0 g3659 (.Z(COL[3]), .A(w3301), .nE(w3914) );
	vdp_bufif0 g3660 (.Z(COL[2]), .A(w3266), .nE(w3914) );
	vdp_bufif0 g3661 (.Z(COL[1]), .A(w3913), .nE(w3914) );
	vdp_bufif0 g3662 (.Z(COL[0]), .A(w3324), .nE(w3914) );
	vdp_nand g3663 (.Z(w3011), .B(HCLK1), .A(w3005) );
	vdp_nand g3664 (.Z(w3017), .B(HCLK1), .A(w3004) );
	vdp_nand g3665 (.Z(w2972), .A(w3503), .B(HCLK1) );
	vdp_nand g3666 (.Z(w2923), .A(w3909), .B(HCLK1) );
	vdp_nor g3667 (.Z(w3910), .A(w3307), .B(w3362) );
	vdp_nand g3668 (.Z(w3020), .A(w3989), .B(HCLK1) );
	vdp_nand g3669 (.Z(w3261), .A(M5), .B(w3265) );
	vdp_nand g3670 (.Z(w3260), .A(M5), .B(w3887) );
	vdp_xor g3671 (.Z(w3424), .A(w3423), .B(w3422) );
	vdp_aon22 g3672 (.Z(w3422), .A1(w3420), .B1(w3498), .A2(VPOS[3]), .B2(w3421) );
	vdp_xnor g3673 (.Z(w3426), .A(w3423), .B(w3499) );
	vdp_aon22 g3674 (.Z(w3499), .A1(w3420), .B1(w3498), .A2(VPOS[2]), .B2(w3425) );
	vdp_xnor g3675 (.Z(w3428), .A(w3423), .B(w3497) );
	vdp_aon22 g3676 (.Z(w3497), .A1(w3420), .B1(w3498), .A2(VPOS[1]), .B2(w3427) );
	vdp_notif0 g3677 (.nZ(VRAMA[4]), .A(w3426), .nE(w3477) );
	vdp_notif0 g3678 (.nZ(VRAMA[3]), .A(w3428), .nE(w3477) );
	vdp_xnor g3679 (.Z(w3495), .A(w3423), .B(w3496) );
	vdp_aon22 g3680 (.Z(w3496), .A1(w3420), .B1(w3498), .A2(VPOS[0]), .B2(w3429) );
	vdp_notif0 g3681 (.nZ(VRAMA[2]), .A(w3495), .nE(w3477) );
	vdp_notif0 g3682 (.nZ(VRAMA[1]), .A(w3494), .nE(w3477) );
	vdp_notif0 g3683 (.nZ(VRAMA[0]), .A(1'b1), .nE(w3477) );
	vdp_not g3684 (.nZ(w3491), .A(w3502) );
	vdp_not g3685 (.nZ(w3477), .A(w3501) );
	vdp_comp_we g3686 (.Z(w3420), .nZ(w3498), .A(w3983) );
	vdp_comp_we g3687 (.Z(w3430), .nZ(w3493), .A(w1) );
	vdp_notif0 g3688 (.nZ(VRAMA[5]), .A(w3432), .nE(w3491) );
	vdp_aoi22 g3689 (.Z(w3432), .A1(w3424), .B1(w3431), .A2(w3430), .B2(w3493) );
	vdp_notif0 g3690 (.nZ(VRAMA[6]), .A(w3433), .nE(w3491) );
	vdp_aoi22 g3691 (.Z(w3433), .A1(w3431), .B1(w3434), .A2(w3430), .B2(w3493) );
	vdp_notif0 g3692 (.nZ(VRAMA[7]), .A(w3435), .nE(w3491) );
	vdp_aoi22 g3693 (.Z(w3435), .A1(w3434), .B1(w3436), .A2(w3430), .B2(w3493) );
	vdp_notif0 g3694 (.nZ(VRAMA[8]), .A(w3437), .nE(w3491) );
	vdp_aoi22 g3695 (.Z(w3437), .A1(w3436), .B1(w3438), .A2(w3430), .B2(w3493) );
	vdp_notif0 g3696 (.nZ(VRAMA[9]), .A(w3917), .nE(w3491) );
	vdp_aoi22 g3697 (.Z(w3917), .A1(w3438), .B1(w3440), .A2(w3430), .B2(w3493) );
	vdp_notif0 g3698 (.nZ(VRAMA[10]), .A(w3439), .nE(w3491) );
	vdp_aoi22 g3699 (.Z(w3439), .A1(w3440), .B1(w3441), .A2(w3430), .B2(w3493) );
	vdp_notif0 g3700 (.nZ(VRAMA[11]), .A(w3916), .nE(w3491) );
	vdp_aoi22 g3701 (.Z(w3916), .A1(w3441), .B1(w3443), .A2(w3430), .B2(w3493) );
	vdp_notif0 g3702 (.nZ(VRAMA[12]), .A(w3444), .nE(w3491) );
	vdp_aoi22 g3703 (.Z(w3444), .A1(w3443), .B1(w3442), .A2(w3430), .B2(w3493) );
	vdp_notif0 g3704 (.nZ(VRAMA[13]), .A(w3446), .nE(w3491) );
	vdp_aoi22 g3705 (.Z(w3446), .A1(w3442), .B1(w3445), .A2(w3430), .B2(w3493) );
	vdp_not g3706 (.nZ(w3492), .A(w3939) );
	vdp_notif0 g3707 (.nZ(VRAMA[14]), .A(w3448), .nE(w3492) );
	vdp_aoi22 g3708 (.Z(w3448), .A1(w3445), .B1(w3447), .A2(w3430), .B2(w3493) );
	vdp_notif0 g3709 (.nZ(VRAMA[15]), .A(w3450), .nE(w3492) );
	vdp_aoi22 g3710 (.Z(w3450), .A1(w3447), .B1(w3449), .A2(w3430), .B2(w3493) );
	vdp_notif0 g3711 (.nZ(VRAMA[16]), .A(w3452), .nE(w3492) );
	vdp_aoi22 g3712 (.Z(w3452), .A1(w3449), .B1(w3451), .A2(w3430), .B2(w3493) );
	vdp_notif0 g3713 (.nZ(VRAMA[5]), .A(w3455), .nE(w3490) );
	vdp_aoi22 g3714 (.Z(w3455), .A1(w3453), .B1(w3424), .A2(w3454), .B2(w3489) );
	vdp_notif0 g3715 (.nZ(VRAMA[6]), .A(w3457), .nE(w3490) );
	vdp_aoi22 g3716 (.Z(w3457), .A1(w3453), .B1(w3454), .A2(w3456), .B2(w3489) );
	vdp_notif0 g3717 (.nZ(VRAMA[7]), .A(w3458), .nE(w3490) );
	vdp_aoi22 g3718 (.Z(w3458), .A1(w3453), .B1(w3456), .A2(w3476), .B2(w3489) );
	vdp_notif0 g3719 (.nZ(VRAMA[8]), .A(w3459), .nE(w3490) );
	vdp_aoi22 g3720 (.Z(w3459), .A1(w3453), .B1(w3476), .A2(w3460), .B2(w3489) );
	vdp_notif0 g3721 (.nZ(VRAMA[9]), .A(w3461), .nE(w3490) );
	vdp_aoi22 g3722 (.Z(w3461), .A1(w3453), .B1(w3460), .A2(w3462), .B2(w3489) );
	vdp_notif0 g3723 (.nZ(VRAMA[10]), .A(w3464), .nE(w3490) );
	vdp_aoi22 g3724 (.Z(w3464), .A1(w3453), .B1(w3462), .A2(w3463), .B2(w3489) );
	vdp_notif0 g3725 (.nZ(VRAMA[11]), .A(w3466), .nE(w3488) );
	vdp_aoi22 g3726 (.Z(w3466), .A1(w3453), .B1(w3463), .A2(w3465), .B2(w3489) );
	vdp_notif0 g3727 (.nZ(VRAMA[12]), .A(w3468), .nE(w3488) );
	vdp_aoi22 g3728 (.Z(w3468), .A1(w3453), .B1(w3465), .A2(w3467), .B2(w3489) );
	vdp_notif0 g3729 (.nZ(VRAMA[14]), .A(w3471), .nE(w3488) );
	vdp_aoi22 g3730 (.Z(w3471), .A1(w3453), .B1(w3469), .A2(w3472), .B2(w3489) );
	vdp_notif0 g3731 (.nZ(VRAMA[15]), .A(w3474), .nE(w3488) );
	vdp_aoi22 g3732 (.Z(w3474), .A1(w3453), .B1(w3472), .A2(w3473), .B2(w3489) );
	vdp_notif0 g3733 (.nZ(VRAMA[16]), .A(w3475), .nE(w3488) );
	vdp_aoi22 g3734 (.Z(w3475), .A1(w3453), .B1(w3473), .A2(w3451), .B2(w3489) );
	vdp_notif0 g3735 (.nZ(VRAMA[13]), .A(w3470), .nE(w3488) );
	vdp_aoi22 g3736 (.Z(w3470), .A1(w3453), .B1(w3467), .A2(w3469), .B2(w3489) );
	vdp_not g3737 (.nZ(w3490), .A(w3419) );
	vdp_comp_we g3738 (.Z(w3489), .nZ(w3453), .A(w1) );
	vdp_aon22 g3739 (.Z(w3451), .A1(w3414), .B1(w3413), .A2(w3415), .B2(w3485) );
	vdp_not g3740 (.nZ(w3488), .A(w3419) );
	vdp_not g3741 (.nZ(w3415), .A(w3485) );
	vdp_sr_bit g3742 (.Q(w3501), .D(w3516), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3743 (.Q(w3485), .D(HPOS[3]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3744 (.Q(w3494), .D(w3552), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3745 (.Q(w3502), .D(w3991), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3746 (.Q(w3500), .D(w3982), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3747 (.Q(w3520), .D(w3981), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3748 (.Q(w3487), .D(w3980), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3749 (.Q(w3956), .D(w3957), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3750 (.Q(w3958), .D(w3956), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3751 (.Q(w3503), .D(w3958), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3752 (.Q(w3534), .D(w94), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3753 (.Q(w3513), .D(w32), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3754 (.Q(w3959), .D(w33), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3755 (.Q(w3574), .D(w3959), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3756 (.Q(w3575), .D(w3513), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3757 (.Q(w3572), .D(w3534), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3758 (.Q(w3576), .D(w3486), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3759 (.Q(w3577), .D(w3065), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3760 (.Q(w3578), .D(w3066), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3761 (.Q(w3579), .D(w3064), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3762 (.Q(w3607), .D(w3063), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3763 (.Q(w3608), .D(w3062), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3764 (.Q(w3511), .D(w3509), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3765 (.Q(w3512), .D(w3511), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3766 (.Q(w3960), .D(w3512), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_aon22 g3767 (.Z(w3525), .A1(H40), .B1(HPOS[8]), .A2(w3523), .B2(w3522) );
	vdp_aon22 g3768 (.Z(w3604), .A1(w3505), .B1(HPOS[8]), .A2(w3525), .B2(w3515) );
	vdp_aon22 g3769 (.Z(w3566), .A1(w3510), .B1(w3523), .A2(w3525), .B2(w3515) );
	vdp_or3 g3770 (.Z(w3573), .A(w3534), .B(w3513), .C(w3959) );
	vdp_or g3771 (.Z(w3526), .A(M5), .B(w3352) );
	vdp_bufif0 g3772 (.Z(VRAMA[1]), .A(w3955), .nE(w3514) );
	vdp_or g3773 (.Z(w3600), .A(w3525), .B(HPOS[4]) );
	vdp_bufif0 g3774 (.Z(VRAMA[2]), .A(w3528), .nE(w3514) );
	vdp_or g3775 (.Z(w3601), .A(w3525), .B(HPOS[5]) );
	vdp_bufif0 g3776 (.Z(VRAMA[3]), .A(w3529), .nE(w3514) );
	vdp_or g3777 (.Z(w3605), .A(w3525), .B(HPOS[6]) );
	vdp_bufif0 g3778 (.Z(VRAMA[4]), .A(w3530), .nE(w3514) );
	vdp_or g3779 (.Z(w3603), .A(w3525), .B(HPOS[7]) );
	vdp_bufif0 g3780 (.Z(VRAMA[5]), .A(w3531), .nE(w3514) );
	vdp_bufif0 g3781 (.Z(VRAMA[5]), .A(w3504), .nE(w3514) );
	vdp_not g3782 (.nZ(w3519), .A(w3412) );
	vdp_not g3783 (.nZ(w3961), .A(HPOS[3]) );
	vdp_dlatch_inv g3784 (.nQ(w3509), .D(w3508), .C(DCLK1), .nC(nDCLK1) );
	vdp_not g3785 (.nZ(w3523), .A(w3938) );
	vdp_not g3786 (.nZ(w3515), .A(w3525) );
	vdp_not g3787 (.nZ(w3522), .A(H40) );
	vdp_not g3788 (.nZ(w3514), .A(w3521) );
	vdp_bufif0 g3789 (.Z(VRAMA[0]), .A(1'b0), .nE(w3514) );
	vdp_or g3790 (.Z(w3521), .A(w3500), .B(w3520) );
	vdp_or g3791 (.Z(w3957), .A(w3518), .B(w6) );
	vdp_nand3 g3792 (.Z(w3571), .A(M5), .B(w3519), .C(HPOS[3]) );
	vdp_nand3 g3793 (.Z(w3532), .A(M5), .B(w3519), .C(w3961) );
	vdp_and g3794 (.Z(w3533), .A(DCLK2), .B(w3960) );
	vdp_and g3795 (.Z(w3507), .A(w3512), .B(DCLK2) );
	vdp_and g3796 (.Z(w3570), .A(w3511), .B(DCLK2) );
	vdp_and g3797 (.Z(w3506), .A(w3509), .B(DCLK2) );
	vdp_and g3798 (.Z(w3939), .A(M5), .B(w3502) );
	vdp_and g3799 (.Z(w3560), .A(HPOS[3]), .B(w3524) );
	vdp_and g3800 (.Z(w3980), .A(w3412), .B(w6) );
	vdp_and g3801 (.Z(w3981), .A(w3519), .B(w6) );
	vdp_and3 g3802 (.Z(w3982), .A(w3518), .B(M5), .C(w3517) );
	vdp_nor g3803 (.Z(w3524), .A(M5), .B(w3525) );
	vdp_nand g3804 (.Z(w3508), .A(w3173), .B(HCLK1) );
	vdp_oai21 g3805 (.A1(HPOS[6]), .A2(HPOS[7]), .B(HPOS[8]), .Z(w3938) );
	vdp_slatch g3806 (.Q(w3549), .D(REG_BUS[0]), .C(w3595), .nC(w3594) );
	vdp_slatch g3807 (.Q(w3545), .D(S[0]), .C(w3590), .nC(w3589) );
	vdp_slatch g3808 (.Q(w3546), .D(S[0]), .C(w3591), .nC(w3588) );
	vdp_slatch g3809 (.Q(w3547), .D(REG_BUS[1]), .C(w3595), .nC(w3594) );
	vdp_slatch g3810 (.Q(w3543), .D(S[1]), .C(w3590), .nC(w3589) );
	vdp_slatch g3811 (.Q(w3615), .D(S[1]), .C(w3591), .nC(w3588) );
	vdp_slatch g3812 (.Q(w3616), .D(REG_BUS[2]), .C(w3595), .nC(w3594) );
	vdp_slatch g3813 (.Q(w3537), .D(S[2]), .C(w3590), .nC(w3589) );
	vdp_slatch g3814 (.Q(w3617), .D(S[2]), .C(w3591), .nC(w3588) );
	vdp_slatch g3815 (.Q(w3613), .D(REG_BUS[3]), .C(w3595), .nC(w3594) );
	vdp_slatch g3816 (.Q(w3612), .D(S[3]), .C(w3590), .nC(w3589) );
	vdp_slatch g3817 (.Q(w4278), .D(S[3]), .C(w3591), .nC(w3588) );
	vdp_slatch g3818 (.Q(w3559), .D(REG_BUS[4]), .C(w3595), .nC(w3594) );
	vdp_slatch g3819 (.Q(w3611), .D(S[4]), .C(w3590), .nC(w3589) );
	vdp_slatch g3820 (.Q(w3610), .D(S[4]), .C(w3591), .nC(w3588) );
	vdp_slatch g3821 (.Q(w3609), .D(REG_BUS[5]), .C(w3595), .nC(w3594) );
	vdp_slatch g3822 (.Q(w3598), .D(S[5]), .C(w3590), .nC(w3589) );
	vdp_slatch g3823 (.Q(w3597), .D(S[5]), .C(w3591), .nC(w3588) );
	vdp_slatch g3824 (.Q(w3596), .D(REG_BUS[6]), .C(w3595), .nC(w3594) );
	vdp_slatch g3825 (.Q(w3592), .D(S[6]), .C(w3590), .nC(w3589) );
	vdp_slatch g3826 (.Q(w3593), .D(S[6]), .C(w3591), .nC(w3588) );
	vdp_slatch g3827 (.Q(w3587), .D(REG_BUS[7]), .C(w3595), .nC(w3594) );
	vdp_slatch g3828 (.Q(w3586), .D(S[7]), .C(w3590), .nC(w3589) );
	vdp_slatch g3829 (.Q(w3585), .D(S[7]), .C(w3591), .nC(w3588) );
	vdp_slatch g3830 (.Q(w3583), .D(S[0]), .C(w3569), .nC(w3580) );
	vdp_slatch g3831 (.Q(w3564), .D(S[0]), .C(w3563), .nC(w3584) );
	vdp_slatch g3832 (.Q(w3568), .D(S[1]), .C(w3563), .nC(w3584) );
	vdp_slatch g3833 (.Q(w3567), .D(S[1]), .C(w3569), .nC(w3580) );
	vdp_slatch g3834 (.Q(w3561), .D(w3587), .C(w3542), .nC(w3541) );
	vdp_slatch g3835 (.Q(w3555), .D(w3596), .C(w3542), .nC(w3541) );
	vdp_slatch g3836 (.Q(w3558), .D(w3609), .C(w3542), .nC(w3541) );
	vdp_slatch g3837 (.Q(w3619), .D(w3559), .C(w3542), .nC(w3541) );
	vdp_slatch g3838 (.Q(w3535), .D(w3613), .C(w3542), .nC(w3541) );
	vdp_slatch g3839 (.Q(w3536), .D(w3616), .C(w3542), .nC(w3541) );
	vdp_slatch g3840 (.Q(w3544), .D(w3547), .C(w3542), .nC(w3541) );
	vdp_slatch g3841 (.Q(w3548), .D(w3549), .C(w3542), .nC(w3541) );
	vdp_fa g3842 (.CI(w3935), .SUM(w3882), .B(w3566), .A(w3582) );
	vdp_fa g3843 (.CO(w3935), .CI(w3565), .SUM(w3759), .B(w3604), .A(w3934) );
	vdp_fa g3844 (.CO(w3934), .CI(w3562), .SUM(w3531), .B(w3603), .A(w3933) );
	vdp_fa g3845 (.CO(w3933), .CI(w3556), .SUM(w3530), .B(w3605), .A(w3606) );
	vdp_fa g3846 (.CO(w3606), .CI(w3557), .SUM(w3529), .B(w3601), .A(w3602) );
	vdp_fa g3847 (.CO(w3602), .CI(w3658), .SUM(w3528), .B(w3600), .A(w3599) );
	vdp_fa g3848 (.CO(w3599), .CI(w3526), .SUM(w3955), .B(w3560), .A(1'b1) );
	vdp_aon222 g3849 (.A1(w3539), .B1(w3527), .C1(w3538), .A2(w3567), .B2(w3568), .C2(1'b0), .Z(w3582) );
	vdp_aon222 g3850 (.A1(w3539), .B1(w3527), .C1(w3538), .A2(w3583), .B2(w3564), .C2(1'b0), .Z(w3565) );
	vdp_aon222 g3851 (.A1(w3539), .B1(w3527), .C1(w3538), .A2(w3585), .B2(w3586), .C2(w3561), .Z(w3562) );
	vdp_aon222 g3852 (.A1(w3539), .B1(w3527), .C1(w3538), .A2(w3593), .B2(w3592), .C2(w3555), .Z(w3556) );
	vdp_aon222 g3853 (.A1(w3539), .B1(w3527), .C1(w3538), .A2(w3597), .B2(w3598), .C2(w3558), .Z(w3557) );
	vdp_aon222 g3854 (.A1(w3539), .B1(w3527), .C1(w3538), .A2(w3610), .B2(w3611), .C2(w3619), .Z(w3658) );
	vdp_aon222 g3855 (.A1(w3539), .B1(w3527), .C1(w3538), .A2(w4278), .B2(w3612), .C2(w3535), .Z(w3352) );
	vdp_aon222 g3856 (.A1(w3539), .B1(w3527), .C1(w3538), .A2(w3617), .B2(w3537), .C2(w3536), .Z(w3051) );
	vdp_aon222 g3857 (.A1(w3539), .B1(w3527), .A2(w3615), .B2(w3543), .C2(w3544), .Z(w3349), .C1(w3538) );
	vdp_aon222 g3858 (.A1(w3539), .B1(w3527), .C1(w3538), .A2(w3546), .B2(w3545), .C2(w3548), .Z(w3347) );
	vdp_comp_strong g3859 (.Z(w3569), .nZ(w3580), .A(w3533) );
	vdp_comp_strong g3860 (.Z(w3563), .nZ(w3584), .A(w3570) );
	vdp_not g3861 (.nZ(w3527), .A(w3532) );
	vdp_not g3862 (.nZ(w3539), .A(w3571) );
	vdp_not g3863 (.nZ(w3538), .A(w3614) );
	vdp_not g3864 (.nZ(w3550), .A(w81) );
	vdp_not g3865 (.nZ(w3517), .A(w89) );
	vdp_not g3866 (.nZ(w3551), .A(w3552) );
	vdp_not g3867 (.nZ(w3518), .A(w3553) );
	vdp_not g3868 (.nZ(w3554), .A(M5) );
	vdp_comp_strong g3869 (.Z(w3590), .nZ(w3589), .A(w3506) );
	vdp_comp_strong g3870 (.Z(w3591), .nZ(w3588), .A(w3507) );
	vdp_comp_strong g3871 (.Z(w3595), .nZ(w3594), .A(w764) );
	vdp_comp_strong g3872 (.Z(w3542), .nZ(w3541), .A(w3618) );
	vdp_or g3873 (.Z(w3614), .A(w3940), .B(M5) );
	vdp_or g3874 (.Z(w3991), .A(w12), .B(w3551) );
	vdp_or g3875 (.Z(w3516), .A(w12), .B(w13) );
	vdp_or g3876 (.Z(w3618), .A(w4), .B(w88) );
	vdp_or5 g3877 (.E(w3550), .C(VPOS[6]), .D(VPOS[5]), .Z(w3940), .A(VPOS[7]), .B(VPOS[4]) );
	vdp_aoi21 g3878 (.Z(w3553), .A1(w89), .A2(w3002), .B(w7) );
	vdp_nand g3879 (.Z(w3552), .A(w13), .B(w3554) );
	vdp_slatch g3880 (.Q(w3653), .D(w4269), .C(w3622), .nC(w3623) );
	vdp_slatch g3881 (.Q(w3628), .D(w4270), .C(w3622), .nC(w3623) );
	vdp_slatch g3882 (.Q(w3629), .D(w4271), .C(w3622), .nC(w3623) );
	vdp_slatch g3883 (.Q(w3630), .D(w4268), .C(w3622), .nC(w3623) );
	vdp_slatch g3884 (.Q(w3632), .D(w4267), .C(w3622), .nC(w3623) );
	vdp_slatch g3885 (.Q(w3631), .D(w4266), .C(w3622), .nC(w3623) );
	vdp_slatch g3886 (.nQ(w3637), .D(w4274), .C(w3624), .nC(w3625) );
	vdp_slatch g3887 (.Q(w3648), .D(w4275), .C(w3624), .nC(w3625) );
	vdp_slatch g3888 (.Q(w3636), .D(w4276), .C(w3624), .nC(w3625) );
	vdp_slatch g3889 (.Q(w3635), .D(w4277), .C(w3624), .nC(w3625) );
	vdp_slatch g3890 (.Q(w3634), .D(w4273), .C(w3624), .nC(w3625) );
	vdp_slatch g3891 (.Q(w3633), .D(w4272), .C(w3624), .nC(w3625) );
	vdp_comp_strong g3892 (.Z(w3622), .nZ(w3623), .A(w3642) );
	vdp_comp_strong g3893 (.Z(w3624), .nZ(w3625), .A(w3962) );
	vdp_cgi2a g3894 (.Z(w3881), .A(w3633), .B(HPOS[4]), .C(1'b1) );
	vdp_cgi2a g3895 (.Z(w3876), .A(w3634), .B(HPOS[5]), .C(w3881) );
	vdp_cgi2a g3896 (.Z(w3875), .A(w3635), .B(HPOS[6]), .C(w3876) );
	vdp_cgi2a g3897 (.Z(w3877), .A(w3636), .B(HPOS[7]), .C(w3875) );
	vdp_cgi2a g3898 (.Z(w3638), .A(w3648), .B(HPOS[8]), .C(w3877) );
	vdp_cgi2a g3899 (.Z(w3643), .A(w3640), .B(w3628), .C(w3964) );
	vdp_cgi2a g3900 (.Z(w3964), .A(w3641), .B(w3629), .C(w3878) );
	vdp_cgi2a g3901 (.Z(w3878), .A(w3644), .B(w3630), .C(w3879) );
	vdp_cgi2a g3902 (.Z(w3879), .A(w3647), .B(w3632), .C(w3880) );
	vdp_cgi2a g3903 (.Z(w3880), .A(w3646), .B(w3631), .C(1'b0) );
	vdp_slatch g3904 (.Q(w4269), .D(REG_BUS[7]), .C(w3650), .nC(w3627) );
	vdp_slatch g3905 (.Q(w4270), .D(REG_BUS[4]), .C(w3650), .nC(w3627) );
	vdp_slatch g3906 (.Q(w4271), .D(REG_BUS[3]), .C(w3650), .nC(w3627) );
	vdp_slatch g3907 (.Q(w4268), .D(REG_BUS[2]), .C(w3650), .nC(w3627) );
	vdp_slatch g3908 (.Q(w4267), .D(REG_BUS[1]), .C(w3650), .nC(w3627) );
	vdp_slatch g3909 (.Q(w4266), .D(REG_BUS[0]), .C(w3650), .nC(w3627) );
	vdp_comp_strong g3910 (.Z(w3650), .nZ(w3627), .A(w793) );
	vdp_slatch g3911 (.Q(w4274), .D(REG_BUS[7]), .C(w3651), .nC(w3649) );
	vdp_slatch g3912 (.Q(w4275), .D(REG_BUS[4]), .C(w3651), .nC(w3649) );
	vdp_slatch g3913 (.Q(w4276), .D(REG_BUS[3]), .C(w3651), .nC(w3649) );
	vdp_slatch g3914 (.Q(w4277), .D(REG_BUS[2]), .C(w3651), .nC(w3649) );
	vdp_slatch g3915 (.Q(w4273), .D(REG_BUS[1]), .C(w3651), .nC(w3649) );
	vdp_slatch g3916 (.Q(w4272), .D(REG_BUS[0]), .C(w3651), .nC(w3649) );
	vdp_comp_strong g3917 (.Z(w3651), .nZ(w3649), .A(w794) );
	vdp_xor g3918 (.Z(w3652), .A(w3653), .B(w3643) );
	vdp_xor g3919 (.Z(w3639), .A(w3637), .B(w3638) );
	vdp_aon22 g3920 (.Z(w3640), .A1(w3645), .B1(w3656), .A2(VPOS[8]), .B2(VPOS[7]) );
	vdp_aon22 g3921 (.Z(w3641), .A1(w3645), .B1(w3656), .A2(VPOS[7]), .B2(VPOS[6]) );
	vdp_aon22 g3922 (.Z(w3644), .A1(w3645), .B1(w3656), .A2(VPOS[6]), .B2(VPOS[5]) );
	vdp_aon22 g3923 (.Z(w3647), .A1(w3645), .B1(w3656), .A2(VPOS[5]), .B2(VPOS[4]) );
	vdp_aon22 g3924 (.Z(w3646), .A1(w3645), .B1(w3656), .A2(VPOS[4]), .B2(VPOS[3]) );
	vdp_aon22 g3925 (.Z(w3663), .A1(w3645), .B1(w3656), .A2(VPOS[3]), .B2(VPOS[2]) );
	vdp_aon22 g3926 (.Z(w3662), .A1(w3645), .B1(w3656), .A2(VPOS[2]), .B2(VPOS[1]) );
	vdp_aon22 g3927 (.Z(w3661), .A1(w3645), .B1(w3656), .A2(VPOS[1]), .B2(VPOS[0]) );
	vdp_comp_we g3928 (.Z(w3645), .nZ(w3656), .A(w1) );
	vdp_not g3929 (.nZ(w3412), .A(w3963) );
	vdp_not g3930 (.nZ(w3655), .A(HPOS[3]) );
	vdp_not g3931 (.nZ(w3966), .A(w3965) );
	vdp_or g3932 (.Z(w3962), .A(w88), .B(w4) );
	vdp_or g3933 (.Z(w3642), .A(w88), .B(w3966) );
	vdp_oai21 g3934 (.Z(w3965), .A1(w5), .A2(M5), .B(w4) );
	vdp_and g3935 (.Z(w3654), .A(w3639), .B(w3657) );
	vdp_oai211 g3936 (.Z(w3963), .A1(w3655), .A2(M5), .B(w3654), .C(w3652) );
	vdp_slatch g3937 (.nQ(w3696), .D(REG_BUS[4]), .C(w3668), .nC(w3669) );
	vdp_slatch g3938 (.nQ(w3698), .D(REG_BUS[4]), .C(w3666), .nC(w3667) );
	vdp_slatch g3939 (.nQ(w3697), .D(REG_BUS[5]), .C(w3668), .nC(w3669) );
	vdp_slatch g3940 (.nQ(w3699), .D(REG_BUS[5]), .C(w3666), .nC(w3667) );
	vdp_slatch g3941 (.nQ(w3672), .D(REG_BUS[6]), .C(w3668), .nC(w3669) );
	vdp_slatch g3942 (.nQ(w3673), .D(REG_BUS[6]), .C(w3666), .nC(w3667) );
	vdp_slatch g3943 (.nQ(w4265), .D(REG_BUS[1]), .C(w3666), .nC(w3667) );
	vdp_slatch g3944 (.nQ(w3692), .D(REG_BUS[2]), .C(w3668), .nC(w3669) );
	vdp_slatch g3945 (.nQ(w3693), .D(REG_BUS[2]), .C(w3666), .nC(w3667) );
	vdp_slatch g3946 (.nQ(w3694), .D(REG_BUS[3]), .C(w3668), .nC(w3669) );
	vdp_slatch g3947 (.nQ(w3695), .D(REG_BUS[3]), .C(w3666), .nC(w3667) );
	vdp_slatch g3948 (.nQ(w3700), .D(REG_BUS[0]), .C(w3666), .nC(w3667) );
	vdp_slatch g3949 (.nQ(w3670), .D(REG_BUS[1]), .C(w3668), .nC(w3669) );
	vdp_slatch g3950 (.Q(w3414), .D(REG_BUS[0]), .C(w3659), .nC(w3660) );
	vdp_slatch g3951 (.Q(w3413), .D(REG_BUS[4]), .C(w3659), .nC(w3660) );
	vdp_not g3952 (.nZ(w3968), .A(w3670) );
	vdp_aoi22 g3953 (.Z(w3689), .A1(HPOS[8]), .B1(w3646), .A2(w3665), .B2(w3664) );
	vdp_aoi22 g3954 (.Z(w3690), .A1(w3646), .B1(w3647), .A2(w3665), .B2(w3664) );
	vdp_aoi22 g3955 (.Z(w3677), .A1(w3647), .B1(w3644), .A2(w3665), .B2(w3664) );
	vdp_aoi22 g3956 (.Z(w3702), .A1(w3641), .B1(w3640), .A2(w3665), .B2(w3664) );
	vdp_aoi22 g3957 (.Z(w3691), .A1(w3644), .B1(w3641), .A2(w3665), .B2(w3664) );
	vdp_comp_strong g3958 (.Z(w3659), .nZ(w3660), .A(w765) );
	vdp_comp_strong g3959 (.Z(w3668), .nZ(w3669), .A(w791) );
	vdp_comp_strong g3960 (.Z(w3666), .nZ(w3667), .A(w1421) );
	vdp_aoi22 g3961 (.Z(w3701), .A1(w3640), .B1(w3664), .A2(w3665), .B2(w3968) );
	vdp_nand g3962 (.Z(w3703), .A(w3640), .B(HSCR) );
	vdp_nand g3963 (.Z(w3676), .A(w3641), .B(HSCR) );
	vdp_nand g3964 (.Z(w3704), .A(w3647), .B(HSCR) );
	vdp_nand g3965 (.Z(w3678), .A(w3644), .B(HSCR) );
	vdp_nand g3966 (.Z(w3688), .A(w3646), .B(HSCR) );
	vdp_nand g3967 (.Z(w3967), .A(w3663), .B(LSCR) );
	vdp_nand g3968 (.Z(w3992), .A(w3662), .B(LSCR) );
	vdp_nand g3969 (.Z(w3684), .A(w3661), .B(LSCR) );
	vdp_nand g3970 (.Z(w3657), .A(HPOS[7]), .B(HPOS[8]) );
	vdp_comp_we g3971 (.Z(w3665), .nZ(w3664), .A(H40) );
	vdp_notif0 g3972 (.nZ(VRAMA[16]), .A(w3673), .nE(w3671) );
	vdp_notif0 g3973 (.nZ(VRAMA[16]), .A(w3672), .nE(w3675) );
	vdp_notif0 g3974 (.nZ(VRAMA[15]), .A(w3699), .nE(w3671) );
	vdp_notif0 g3975 (.nZ(VRAMA[15]), .A(w3697), .nE(w3675) );
	vdp_notif0 g3976 (.nZ(VRAMA[14]), .A(w3698), .nE(w3671) );
	vdp_notif0 g3977 (.nZ(VRAMA[14]), .A(w3696), .nE(w3675) );
	vdp_notif0 g3978 (.nZ(VRAMA[13]), .A(w3695), .nE(w3671) );
	vdp_notif0 g3979 (.nZ(VRAMA[13]), .A(w3694), .nE(w3675) );
	vdp_notif0 g3980 (.nZ(VRAMA[12]), .A(w3693), .nE(w3671) );
	vdp_notif0 g3981 (.nZ(VRAMA[12]), .A(w3692), .nE(w3675) );
	vdp_notif0 g3982 (.nZ(VRAMA[11]), .A(w4265), .nE(w3671) );
	vdp_notif0 g3983 (.nZ(VRAMA[11]), .A(w3701), .nE(w3675) );
	vdp_notif0 g3984 (.nZ(VRAMA[10]), .A(w3700), .nE(w3671) );
	vdp_notif0 g3985 (.nZ(VRAMA[10]), .A(w3702), .nE(w3675) );
	vdp_notif0 g3986 (.nZ(VRAMA[9]), .A(w3703), .nE(w3674) );
	vdp_notif0 g3987 (.nZ(VRAMA[9]), .A(w3691), .nE(w3675) );
	vdp_notif0 g3988 (.nZ(VRAMA[6]), .A(w3704), .nE(w3674) );
	vdp_notif0 g3989 (.nZ(VRAMA[6]), .A(w3689), .nE(w3679) );
	vdp_notif0 g3990 (.nZ(VRAMA[5]), .A(w3688), .nE(w3674) );
	vdp_notif0 g3991 (.nZ(VRAMA[5]), .A(w3687), .nE(w3679) );
	vdp_notif0 g3992 (.nZ(VRAMA[4]), .A(w3967), .nE(w3674) );
	vdp_notif0 g3993 (.nZ(VRAMA[4]), .A(w3686), .nE(w3679) );
	vdp_notif0 g3994 (.nZ(VRAMA[3]), .A(w3992), .nE(w3674) );
	vdp_notif0 g3995 (.nZ(VRAMA[3]), .A(w3685), .nE(w3679) );
	vdp_notif0 g3996 (.nZ(VRAMA[2]), .A(w3684), .nE(w3674) );
	vdp_notif0 g3997 (.nZ(VRAMA[2]), .A(w3683), .nE(w3679) );
	vdp_notif0 g3998 (.nZ(VRAMA[1]), .A(1'b1), .nE(w3674) );
	vdp_notif0 g3999 (.nZ(VRAMA[1]), .A(1'b1), .nE(w3679) );
	vdp_notif0 g4000 (.nZ(VRAMA[0]), .A(w3681), .nE(w3674) );
	vdp_notif0 g4001 (.nZ(VRAMA[0]), .A(w3681), .nE(w3679) );
	vdp_notif0 g4002 (.nZ(VRAMA[8]), .A(w3676), .nE(w3674) );
	vdp_notif0 g4003 (.nZ(VRAMA[8]), .A(w3677), .nE(w3679) );
	vdp_notif0 g4004 (.nZ(VRAMA[7]), .A(w3678), .nE(w3674) );
	vdp_notif0 g4005 (.nZ(VRAMA[7]), .A(w3690), .nE(w3679) );
	vdp_not g4006 (.nZ(w3681), .A(1'b0) );
	vdp_not g4007 (.nZ(w3683), .A(HPOS[4]) );
	vdp_not g4008 (.nZ(w3685), .A(HPOS[5]) );
	vdp_not g4009 (.nZ(w3686), .A(HPOS[6]) );
	vdp_not g4010 (.nZ(w3687), .A(HPOS[7]) );
	vdp_not g4011 (.nZ(w3674), .A(w3172) );
	vdp_not g4012 (.nZ(w3671), .A(w3172) );
	vdp_not g4013 (.nZ(w3679), .A(w3487) );
	vdp_not g4014 (.nZ(w3675), .A(w3487) );
	vdp_not g4015 (.nZ(w3711), .A(w3874) );
	vdp_comp_strong g4016 (.Z(w3705), .nZ(w3706), .A(w790) );
	vdp_comp_we g4017 (.Z(w3710), .nZ(w3709), .A(w3500) );
	vdp_comp_strong g4018 (.Z(w3708), .nZ(w3707), .A(w792) );
	vdp_slatch g4019 (.Q(w3731), .D(REG_BUS[6]), .C(w3705), .nC(w3706) );
	vdp_slatch g4020 (.Q(w3977), .D(REG_BUS[3]), .C(w3708), .nC(w3707) );
	vdp_slatch g4021 (.Q(w3730), .D(REG_BUS[5]), .C(w3705), .nC(w3706) );
	vdp_slatch g4022 (.Q(w3728), .D(REG_BUS[2]), .C(w3708), .nC(w3707) );
	vdp_slatch g4023 (.Q(w3714), .D(REG_BUS[4]), .C(w3705), .nC(w3706) );
	vdp_slatch g4024 (.Q(w4279), .D(REG_BUS[1]), .C(w3708), .nC(w3707) );
	vdp_slatch g4025 (.Q(w3717), .D(REG_BUS[3]), .C(w3705), .nC(w3706) );
	vdp_slatch g4026 (.Q(w3978), .D(REG_BUS[0]), .C(w3708), .nC(w3707) );
	vdp_slatch g4027 (.Q(w3725), .D(REG_BUS[1]), .C(w3705), .nC(w3706) );
	vdp_slatch g4028 (.Q(w3722), .D(REG_BUS[2]), .C(w3705), .nC(w3706) );
	vdp_bufif0 g4029 (.Z(VRAMA[11]), .A(w3724), .nE(w3713) );
	vdp_bufif0 g4030 (.Z(VRAMA[10]), .A(w3718), .nE(w3713) );
	vdp_bufif0 g4031 (.Z(VRAMA[13]), .A(w3726), .nE(w3713) );
	vdp_bufif0 g4032 (.Z(VRAMA[9]), .A(w3716), .nE(w3713) );
	vdp_bufif0 g4033 (.Z(VRAMA[8]), .A(w3715), .nE(w3713) );
	vdp_bufif0 g4034 (.Z(VRAMA[14]), .A(w3727), .nE(w3711) );
	vdp_bufif0 g4035 (.Z(VRAMA[7]), .A(w3712), .nE(w3713) );
	vdp_bufif0 g4036 (.Z(VRAMA[15]), .A(w3937), .nE(w3711) );
	vdp_bufif0 g4037 (.Z(VRAMA[16]), .A(w3729), .nE(w3711) );
	vdp_aon22 g4038 (.Z(w3729), .A1(w3709), .B1(w3710), .A2(w3731), .B2(w3977) );
	vdp_aon22 g4039 (.Z(w3937), .A1(w3709), .B1(w3710), .A2(w3730), .B2(w3728) );
	vdp_aon22 g4040 (.Z(w3727), .A1(w3709), .B1(w3710), .A2(w3714), .B2(w4279) );
	vdp_aon22 g4041 (.Z(w3726), .A1(w3709), .B1(w3710), .A2(w3717), .B2(w3978) );
	vdp_aon22 g4042 (.Z(w3724), .A1(w3720), .B1(w3723), .A2(w3725), .B2(w3721) );
	vdp_aon22 g4043 (.Z(w3719), .A1(w3720), .B1(w3733), .A2(w3722), .B2(w3721) );
	vdp_bufif0 g4044 (.Z(VRAMA[12]), .A(w3719), .nE(w3713) );
	vdp_not g4045 (.nZ(w3713), .A(w3521) );
	vdp_and g4046 (.Z(w3874), .A(w3521), .B(M5) );
	vdp_comp_we g4047 (.Z(w3721), .nZ(w3720), .A(M5) );
	vdp_fa g4048 (.CO(w3748), .CI(w3924), .SUM(w3768), .B(VPOS[6]), .A(w3923) );
	vdp_fa g4049 (.CO(w3923), .CI(w3926), .SUM(w3749), .B(VPOS[5]), .A(w3925) );
	vdp_fa g4050 (.CO(w3925), .CI(w3928), .SUM(w3750), .B(VPOS[4]), .A(w3927) );
	vdp_fa g4051 (.CO(w3927), .CI(w3816), .SUM(w3421), .B(VPOS[3]), .A(w3929) );
	vdp_fa g4052 (.CO(w3929), .CI(w3931), .SUM(w3425), .B(VPOS[2]), .A(w3930) );
	vdp_fa g4053 (.CO(w3930), .CI(w3869), .SUM(w3427), .B(VPOS[1]), .A(w3932) );
	vdp_fa g4054 (.CO(w3932), .CI(w3829), .SUM(w3429), .B(VPOS[0]), .A(1'b0) );
	vdp_fa g4055 (.CO(w3767), .CI(w3922), .SUM(w3765), .B(VPOS[7]), .A(w3748) );
	vdp_fa g4056 (.CO(w3747), .CI(w3802), .SUM(w3776), .B(VPOS[8]), .A(w3767) );
	vdp_fa g4057 (.CO(w3775), .CI(w3803), .SUM(w3742), .B(1'b0), .A(w3747) );
	vdp_fa g4058 (.CI(w3787), .SUM(w3743), .B(1'b0), .A(w3775) );
	vdp_aon22 g4059 (.Z(w3787), .A1(w3785), .B1(w3786), .A2(w3746), .B2(w3745) );
	vdp_aon22 g4060 (.Z(w3803), .A1(w3872), .B1(w3790), .A2(w3746), .B2(w3745) );
	vdp_aon22 g4061 (.Z(w3802), .A1(w3791), .B1(w3792), .A2(w3746), .B2(w3745) );
	vdp_aon22 g4062 (.Z(w3922), .A1(w3794), .B1(w3795), .A2(w3746), .B2(w3745) );
	vdp_aon22 g4063 (.Z(w3924), .A1(w3801), .B1(w3798), .A2(w3746), .B2(w3745) );
	vdp_aon22 g4064 (.Z(w3926), .A1(w3806), .B1(w3805), .A2(w3746), .B2(w3745) );
	vdp_aon22 g4065 (.Z(w3928), .A1(w3810), .B1(w3811), .A2(w3746), .B2(w3745) );
	vdp_aon22 g4066 (.Z(w3816), .A1(w3815), .B1(w3814), .A2(w3746), .B2(w3745) );
	vdp_aon22 g4067 (.Z(w3931), .A1(w3817), .B1(w3818), .A2(w3746), .B2(w3745) );
	vdp_aon22 g4068 (.Z(w3869), .A1(w3821), .B1(w3873), .A2(w3746), .B2(w3745) );
	vdp_aon22 g4069 (.Z(w3829), .A1(w3823), .B1(w3822), .A2(w3746), .B2(w3745) );
	vdp_comp_we g4070 (.Z(w3746), .nZ(w3745), .A(w3754) );
	vdp_comp_strong g4071 (.Z(w3756), .nZ(w3751), .A(w779) );
	vdp_sr_bit g4072 (.Q(w3777), .D(RD_DATA[1]), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4073 (.Q(w3752), .D(RD_DATA[2]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4074 (.Q(w3826), .D(w3777), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4075 (.Q(w3840), .D(w3752), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4076 (.Q(w3825), .D(HPOS[3]), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4077 (.Q(w3505), .D(REG_BUS[0]), .C(w3756), .nC(w3751) );
	vdp_slatch g4078 (.Q(w3510), .D(REG_BUS[1]), .C(w3756), .nC(w3751) );
	vdp_slatch g4079 (.Q(w3772), .D(REG_BUS[5]), .C(w3756), .nC(w3751) );
	vdp_slatch g4080 (.Q(w3771), .D(REG_BUS[4]), .C(w3756), .nC(w3751) );
	vdp_slatch g4081 (.Q(w3823), .D(w3827), .C(w3778), .nC(w3782) );
	vdp_slatch g4082 (.Q(w3988), .D(w3828), .C(w3784), .nC(w3779) );
	vdp_slatch g4083 (.Q(w3821), .D(w3820), .C(w3778), .nC(w3782) );
	vdp_slatch g4084 (.Q(w3987), .D(w3819), .C(w3784), .nC(w3779) );
	vdp_slatch g4085 (.Q(w3817), .D(w3842), .C(w3778), .nC(w3782) );
	vdp_slatch g4086 (.Q(w3986), .D(w3813), .C(w3784), .nC(w3779) );
	vdp_slatch g4087 (.Q(w3815), .D(w3812), .C(w3778), .nC(w3782) );
	vdp_slatch g4088 (.Q(w3985), .D(w3809), .C(w3784), .nC(w3779) );
	vdp_slatch g4089 (.Q(w3810), .D(w3808), .C(w3778), .nC(w3782) );
	vdp_slatch g4090 (.Q(w3984), .D(w3807), .C(w3784), .nC(w3779) );
	vdp_slatch g4091 (.Q(w3806), .D(w3800), .C(w3778), .nC(w3782) );
	vdp_slatch g4092 (.Q(w3995), .D(w3799), .C(w3784), .nC(w3779) );
	vdp_slatch g4093 (.Q(w3801), .D(w3796), .C(w3778), .nC(w3782) );
	vdp_slatch g4094 (.Q(w3996), .D(w3797), .C(w3784), .nC(w3779) );
	vdp_slatch g4095 (.Q(w3794), .D(w3793), .C(w3778), .nC(w3782) );
	vdp_slatch g4096 (.Q(w3792), .D(w3804), .C(w3784), .nC(w3779) );
	vdp_slatch g4097 (.Q(w3791), .D(w3847), .C(w3778), .nC(w3782) );
	vdp_slatch g4098 (.Q(w3790), .D(w3789), .C(w3784), .nC(w3779) );
	vdp_slatch g4099 (.Q(w3872), .D(w3788), .C(w3778), .nC(w3782) );
	vdp_slatch g4100 (.Q(w3786), .D(w3936), .C(w3784), .nC(w3779) );
	vdp_slatch g4101 (.Q(w3785), .D(w3783), .C(w3778), .nC(w3782) );
	vdp_slatch g4102 (.Q(w3971), .D(REG_BUS[0]), .C(w3831), .nC(w3830) );
	vdp_aon22 g4103 (.Z(w3824), .A1(w3827), .B1(w3839), .A2(w3841), .B2(w3971) );
	vdp_slatch g4104 (.Q(w3843), .D(REG_BUS[1]), .C(w3831), .nC(w3830) );
	vdp_aon22 g4105 (.Z(w3828), .A1(w3820), .B1(w3839), .A2(w3841), .B2(w3843) );
	vdp_slatch g4106 (.Q(w3970), .D(REG_BUS[2]), .C(w3831), .nC(w3830) );
	vdp_aon22 g4107 (.Z(w3819), .A1(w3842), .B1(w3839), .A2(w3841), .B2(w3970) );
	vdp_slatch g4108 (.Q(w3844), .D(REG_BUS[3]), .C(w3831), .nC(w3830) );
	vdp_aon22 g4109 (.Z(w3813), .A1(w3812), .B1(w3839), .A2(w3841), .B2(w3844) );
	vdp_slatch g4110 (.Q(w3845), .D(REG_BUS[4]), .C(w3831), .nC(w3830) );
	vdp_aon22 g4111 (.Z(w3809), .A1(w3808), .B1(w3839), .A2(w3841), .B2(w3845) );
	vdp_slatch g4112 (.Q(w3870), .D(REG_BUS[5]), .C(w3831), .nC(w3830) );
	vdp_aon22 g4113 (.Z(w3807), .A1(w3800), .B1(w3839), .A2(w3841), .B2(w3870) );
	vdp_slatch g4114 (.Q(w3969), .D(REG_BUS[6]), .C(w3831), .nC(w3830) );
	vdp_aon22 g4115 (.Z(w3799), .A1(w3796), .B1(w3839), .A2(w3841), .B2(w3969) );
	vdp_slatch g4116 (.Q(w3846), .D(REG_BUS[7]), .C(w3831), .nC(w3830) );
	vdp_aon22 g4117 (.Z(w3797), .A1(w3793), .B1(w3839), .A2(w3841), .B2(w3846) );
	vdp_aon22 g4118 (.Z(w3804), .A1(w3847), .B1(w3839), .A2(w3841), .B2(1'b0) );
	vdp_aon22 g4119 (.Z(w3789), .A1(w3788), .B1(w3839), .A2(w3841), .B2(1'b0) );
	vdp_aon22 g4120 (.Z(w3936), .A1(w3783), .B1(w3839), .A2(w3841), .B2(1'b0) );
	vdp_notif0 g4121 (.nZ(RD_DATA[2]), .A(w3862), .nE(w3835) );
	vdp_slatch g4122 (.nQ(w3862), .D(w3783), .C(w3834), .nC(w3833) );
	vdp_notif0 g4123 (.nZ(RD_DATA[1]), .A(w3848), .nE(w3835) );
	vdp_slatch g4124 (.nQ(w3848), .D(w3788), .C(w3834), .nC(w3833) );
	vdp_notif0 g4125 (.nZ(RD_DATA[0]), .A(w3994), .nE(w3835) );
	vdp_slatch g4126 (.nQ(w3994), .D(w3847), .C(w3834), .nC(w3833) );
	vdp_notif0 g4127 (.nZ(AD_DATA[7]), .A(w4285), .nE(w3835) );
	vdp_slatch g4128 (.nQ(w4285), .D(w3793), .C(w3834), .nC(w3833) );
	vdp_notif0 g4129 (.nZ(AD_DATA[6]), .A(w3849), .nE(w3835) );
	vdp_slatch g4130 (.nQ(w3849), .D(w3796), .C(w3834), .nC(w3833) );
	vdp_notif0 g4131 (.nZ(AD_DATA[5]), .A(w3850), .nE(w3835) );
	vdp_slatch g4132 (.nQ(w3850), .D(w3800), .C(w3834), .nC(w3833) );
	vdp_notif0 g4133 (.nZ(AD_DATA[4]), .A(w3851), .nE(w3835) );
	vdp_slatch g4134 (.nQ(w3851), .D(w3808), .C(w3834), .nC(w3833) );
	vdp_notif0 g4135 (.nZ(AD_DATA[3]), .A(w3860), .nE(w3835) );
	vdp_slatch g4136 (.nQ(w3860), .D(w3812), .C(w3834), .nC(w3833) );
	vdp_notif0 g4137 (.nZ(AD_DATA[2]), .A(w3858), .nE(w3835) );
	vdp_slatch g4138 (.nQ(w3858), .D(w3842), .C(w3834), .nC(w3833) );
	vdp_notif0 g4139 (.nZ(AD_DATA[1]), .A(w3853), .nE(w3835) );
	vdp_slatch g4140 (.nQ(w3853), .D(w3820), .C(w3834), .nC(w3833) );
	vdp_notif0 g4141 (.nZ(AD_DATA[0]), .A(w3857), .nE(w3835) );
	vdp_slatch g4142 (.nQ(w3857), .D(w3827), .C(w3834), .nC(w3833) );
	vdp_sr_bit g4143 (.Q(w3856), .D(w3572), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4144 (.Q(w3863), .D(w3867), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4145 (.Q(w3867), .D(RD_DATA[0]), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4146 (.Q(w3993), .D(w3824), .C(w3784), .nC(w3779) );
	vdp_comp_strong g4147 (.Z(w3784), .nZ(w3779), .A(w3838) );
	vdp_comp_strong g4148 (.Z(w3778), .nZ(w3782), .A(w3836) );
	vdp_comp_strong g4149 (.Z(w3831), .nZ(w3830), .A(w763) );
	vdp_sr_bit g4150 (.Q(w3780), .D(w3974), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_comp_strong g4151 (.Z(w3834), .nZ(w3833), .A(w3855) );
	vdp_not g4152 (.nZ(w3835), .A(w3856) );
	vdp_and g4153 (.Z(w3855), .A(w3572), .B(HCLK1) );
	vdp_and g4154 (.Z(w3795), .A(w3996), .B(w3780) );
	vdp_and g4155 (.Z(w3798), .A(w3995), .B(w3780) );
	vdp_and g4156 (.Z(w3805), .A(w3984), .B(w3780) );
	vdp_and g4157 (.Z(w3811), .A(w3985), .B(w3780) );
	vdp_and g4158 (.Z(w3814), .A(w3986), .B(w3780) );
	vdp_and g4159 (.Z(w3818), .A(w3987), .B(w3780) );
	vdp_and g4160 (.Z(w3873), .A(w3988), .B(w3780) );
	vdp_and g4161 (.Z(w3822), .A(w3993), .B(w3780) );
	vdp_not g4162 (.nZ(w3973), .A(w3972) );
	vdp_not g4163 (.nZ(w3836), .A(w3837) );
	vdp_not g4164 (.nZ(w3754), .A(w3753) );
	vdp_not g4165 (.nZ(w3758), .A(w3505) );
	vdp_not g4166 (.nZ(w3757), .A(w3510) );
	vdp_not g4167 (.nZ(w3735), .A(w3975) );
	vdp_not g4168 (.nZ(w3734), .A(w3976) );
	vdp_not g4169 (.nZ(w3736), .A(w3979) );
	vdp_not g4170 (.nZ(w3921), .A(M5) );
	vdp_not g4171 (.nZ(w3774), .A(w3920) );
	vdp_aon22 g4172 (.Z(w3762), .A1(w3741), .B1(w3749), .A2(w3768), .B2(w3744) );
	vdp_aon22 g4173 (.Z(w3766), .A1(w3741), .B1(w3768), .A2(w3765), .B2(w3744) );
	vdp_ha g4174 (.CO(w3770), .SUM(w3740), .B(w3769), .A(w3766) );
	vdp_aon222 g4175 (.A1(w3736), .B1(w3734), .C1(w3735), .A2(w3764), .B2(w3763), .C2(w3740), .Z(w3716) );
	vdp_aon22 g4176 (.Z(w3919), .A1(w3741), .B1(w3765), .A2(w3776), .B2(w3744) );
	vdp_ha g4177 (.SUM(w3739), .B(w3770), .A(w3919) );
	vdp_aon222 g4178 (.A1(w3736), .B1(w3734), .C1(w3735), .A2(w3763), .B2(w3740), .C2(w3739), .Z(w3718) );
	vdp_ha g4179 (.CO(w3769), .SUM(w3763), .B(w3762), .A(w3773) );
	vdp_aon222 g4180 (.A1(w3736), .B1(w3734), .C1(w3735), .A2(w3760), .B2(w3764), .C2(w3763), .Z(w3715) );
	vdp_aon22 g4181 (.Z(w3764), .A1(w3741), .B1(w3750), .A2(w3749), .B2(w3744) );
	vdp_aon222 g4182 (.A1(w3736), .B1(w3734), .C1(w3735), .A2(w3882), .B2(w3760), .C2(w3764), .Z(w3712) );
	vdp_aon222 g4183 (.A1(w3736), .B1(w3734), .C1(w3735), .A2(w3759), .B2(w3759), .C2(w3760), .Z(w3504) );
	vdp_aon22 g4184 (.Z(w3760), .A1(w3741), .B1(w3421), .A2(w3750), .B2(w3744) );
	vdp_comp_we g4185 (.Z(w3841), .nZ(w3839), .A(M5) );
	vdp_comp_we g4186 (.Z(w3741), .nZ(w3744), .A(w1) );
	vdp_and g4187 (.Z(w3773), .A(w3774), .B(w3921) );
	vdp_aon222 g4188 (.A1(w3736), .B1(w3734), .C1(w3735), .A2(w3740), .B2(w3739), .C2(w3737), .Z(w3723) );
	vdp_aon222 g4189 (.A1(w3736), .B1(w3734), .C1(w3735), .A2(w3739), .B2(w3737), .C2(w3918), .Z(w3733) );
	vdp_aon22 g4190 (.Z(w3738), .A1(w3741), .B1(w3742), .A2(w3743), .B2(w3744) );
	vdp_aon22 g4191 (.Z(w3761), .A1(w3741), .B1(w3776), .A2(w3742), .B2(w3744) );
	vdp_and g4192 (.Z(w3737), .B(w3761), .A(w3771) );
	vdp_and g4193 (.Z(w3918), .B(w3738), .A(w3772) );
	vdp_oai21 g4194 (.Z(w3753), .A1(VSCR), .A2(w3825), .B(M5) );
	vdp_aoi21 g4195 (.Z(w3837), .A1(HCLK1), .A2(w15), .B(w88) );
	vdp_oai211 g4196 (.Z(w3972), .A1(HCLK1), .A2(w4), .B(w5), .C(M5) );
	vdp_or g4197 (.Z(w3838), .A(w88), .B(w3973) );
	vdp_nand3 g4198 (.Z(w3974), .A(w80), .B(HPOS[6]), .C(HPOS[7]) );
	vdp_nand g4199 (.Z(w3979), .A(w3510), .B(w3505) );
	vdp_nand g4200 (.Z(w3976), .A(w3505), .B(w3757) );
	vdp_nand g4201 (.Z(w3975), .A(w3757), .B(w3758) );
	vdp_aoi31 g4202 (.Z(w3920), .B3(w3919), .B2(w3766), .B1(w3762), .A(w3761) );
	vdp_slatch g4203 (.Q(w3454), .D(S[0]), .C(w3416), .nC(w3045) );
	vdp_slatch g4204 (.Q(w3456), .D(S[1]), .C(w3416), .nC(w3045) );
	vdp_slatch g4205 (.Q(w3476), .D(S[2]), .C(w3416), .nC(w3045) );
	vdp_slatch g4206 (.Q(w3460), .D(S[3]), .C(w3416), .nC(w3045) );
	vdp_slatch g4207 (.Q(w3462), .D(S[4]), .C(w3416), .nC(w3045) );
	vdp_slatch g4208 (.Q(w3463), .D(S[5]), .C(w3416), .nC(w3045) );
	vdp_slatch g4209 (.Q(w3465), .D(S[6]), .C(w3416), .nC(w3045) );
	vdp_slatch g4210 (.Q(w3467), .D(S[7]), .C(w3416), .nC(w3045) );
	vdp_slatch g4211 (.Q(w3469), .D(S[0]), .C(w3411), .nC(w3410) );
	vdp_slatch g4212 (.Q(w3472), .D(S[1]), .C(w3411), .nC(w3410) );
	vdp_slatch g4213 (.Q(w3473), .D(S[2]), .C(w3411), .nC(w3410) );
	vdp_slatch g4214 (.Q(w2992), .D(S[3]), .C(w3411), .nC(w3410) );
	vdp_slatch g4215 (.Q(w3480), .D(S[4]), .C(w3411), .nC(w3410) );
	vdp_slatch g4216 (.Q(w2969), .D(S[5]), .C(w3411), .nC(w3410) );
	vdp_slatch g4217 (.Q(w2971), .D(S[6]), .C(w3411), .nC(w3410) );
	vdp_slatch g4218 (.Q(w2997), .D(S[7]), .C(w3411), .nC(w3410) );
	vdp_comp_strong g4219 (.Z(w3411), .nZ(w3410), .A(w3179) );
	vdp_comp_strong g4220 (.Z(w3416), .nZ(w3045), .A(w3180) );
	vdp_comp_strong g4221 (.Z(w3417), .nZ(w3478), .A(w3181) );
	vdp_slatch g4222 (.Q(w3954), .D(S[7]), .C(w3417), .nC(w3478) );
	vdp_slatch g4223 (.Q(w3953), .D(S[6]), .C(w3417), .nC(w3478) );
	vdp_slatch g4224 (.Q(w3952), .D(S[5]), .C(w3417), .nC(w3478) );
	vdp_slatch g4225 (.Q(w3483), .D(S[4]), .C(w3417), .nC(w3478) );
	vdp_slatch g4226 (.Q(w3951), .D(S[3]), .C(w3417), .nC(w3478) );
	vdp_slatch g4227 (.Q(w3449), .D(S[2]), .C(w3417), .nC(w3478) );
	vdp_slatch g4228 (.Q(w3447), .D(S[1]), .C(w3417), .nC(w3478) );
	vdp_slatch g4229 (.Q(w3445), .D(S[0]), .C(w3417), .nC(w3478) );
	vdp_slatch g4230 (.Q(w3442), .D(S[7]), .C(w3418), .nC(w3479) );
	vdp_slatch g4231 (.Q(w3443), .D(S[6]), .C(w3418), .nC(w3479) );
	vdp_slatch g4232 (.Q(w3441), .D(S[5]), .C(w3418), .nC(w3479) );
	vdp_slatch g4233 (.Q(w3440), .D(S[4]), .C(w3418), .nC(w3479) );
	vdp_slatch g4234 (.Q(w3438), .D(S[3]), .C(w3418), .nC(w3479) );
	vdp_slatch g4235 (.Q(w3436), .D(S[2]), .C(w3418), .nC(w3479) );
	vdp_slatch g4236 (.Q(w3434), .D(S[1]), .C(w3418), .nC(w3479) );
	vdp_slatch g4237 (.Q(w3431), .D(S[0]), .C(w3418), .nC(w3479) );
	vdp_sr_bit g4238 (.Q(w3983), .D(w3412), .C1(HCLK2), .C2(HCLK1), .nC2(nHCLK1), .nC1(nHCLK2) );
	vdp_sr_bit g4239 (.Q(w3419), .D(w3950), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and g4240 (.Z(w3950), .A(w13), .B(M5) );
	vdp_not g4241 (.nZ(w3949), .A(w3419) );
	vdp_aon22 g4242 (.Z(w2996), .A1(w3954), .B1(w3483), .A2(w3482), .B2(w3912) );
	vdp_aon22 g4243 (.Z(w2993), .A1(w3953), .B1(1'b0), .A2(w3482), .B2(w3912) );
	vdp_aon22 g4244 (.Z(w3481), .A1(w3483), .B1(w3449), .A2(w3482), .B2(w3912) );
	vdp_aon22 g4245 (.Z(w2967), .A1(w3951), .B1(w3447), .A2(w3482), .B2(w3912) );
	vdp_aon22 g4246 (.Z(w2970), .A1(w3952), .B1(w3951), .A2(w3482), .B2(w3912) );
	vdp_comp_strong g4247 (.Z(w3418), .nZ(w3479), .A(w3182) );
	vdp_comp_we g4248 (.Z(w3482), .nZ(w3912), .A(M5) );
	vdp_aon22 g4249 (.Z(w3423), .A1(w3480), .B1(w3481), .A2(w3419), .B2(w3949) );
	vdp_sr_bit g4250 (.Q(w3864), .D(FIFOo[0]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4251 (.Q(w3868), .D(FIFOo[1]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4252 (.Q(w3866), .D(FIFOo[2]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4253 (.Q(w3865), .D(FIFOo[3]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4254 (.Q(w3854), .D(FIFOo[4]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4255 (.Q(w3852), .D(FIFOo[5]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4256 (.Q(w3859), .D(FIFOo[6]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4257 (.Q(w3861), .D(FIFOo[7]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_aon22 g4258 (.Z(w1343), .B1(w4327), .A1(w1373), .B2(w4345), .A2(w40) );
	vdp_not g4259 (.nZ(w4345), .A(w40) );
	vdp_not g4260 (.nZ(w4317), .A(w4306) );
	vdp_not g4261 (.nZ(w4316), .A(w4317) );
	vdp_not g4262 (.nZ(w4315), .A(w4316) );
	vdp_not g4263 (.nZ(w4314), .A(w4315) );
	vdp_and g4264 (.Z(w4327), .B(w4318), .A(w4322) );
	vdp_not g4265 (.nZ(w4318), .A(w4321) );
	vdp_not g4266 (.nZ(w4321), .A(w4320) );
	vdp_not g4267 (.nZ(w4320), .A(w4319) );
	vdp_not g4268 (.nZ(w4319), .A(w4322) );
	vdp_or g4269 (.Z(w4322), .B(w4304), .A(w4303) );
	vdp_dff g4270 (.Q(w4304), .R(w4293), .D(w4303), .C(w4302) );
	vdp_not g4271 (.nZ(w4302), .A(w4323) );
	vdp_nor g4272 (.Z(w4301), .B(w4324), .A(w4303) );
	vdp_dff g4273 (.Q(w4303), .R(w4293), .D(w4324), .C(w4323) );
	vdp_dff g4274 (.Q(w4324), .R(w4293), .D(w4301), .C(w4323) );
	vdp_not g4275 (.nZ(w4323), .A(w4312) );
	vdp_not g4276 (.nZ(w4299), .A(w4312) );
	vdp_dff g4277 (.Q(w4296), .R(w4293), .D(w4325), .C(w4295) );
	vdp_dff g4278 (.Q(w4325), .R(w4293), .D(w4294), .C(w4292) );
	vdp_not g4279 (.nZ(w4292), .A(w4333) );
	vdp_dff g4280 (.Q(w4294), .R(w4293), .D(w4313), .C(w4292) );
	vdp_not g4281 (.nZ(w4295), .A(w4292) );
	vdp_nor g4282 (.Z(w4352), .B(w4328), .A(w4329) );
	vdp_nor g4283 (.Z(w4330), .B(w4328), .A(H40) );
	vdp_not g4284 (.nZ(w4329), .A(H40) );
	vdp_not g4285 (.nZ(w4307), .A(PAL) );
	vdp_aoi222 g4286 (.Z(w4300), .B1(w4332), .A1(w4331), .B2(w4352), .A2(w4328), .C1(w4299), .C2(w4330) );
	vdp_not g4287 (.nZ(EDCLK_O), .A(w4300) );
	vdp_or g4288 (.Z(w4326), .B(w4296), .A(w4325) );
	vdp_nor g4289 (.Z(w4313), .B(w4294), .A(w4325) );
	vdp_not g4290 (.nZ(w4289), .A(w4351) );
	vdp_nand g4291 (.Z(w4308), .B(w4289), .A(w4288) );
	vdp_sr_bit g4292 (.Q(w4351), .D(w4288), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_not g4293 (.nZ(w4350), .A(w4336) );
	vdp_not g4294 (.nZ(w1119), .A(w4349) );
	vdp_not g4295 (.nZ(SYSRES), .A(w4350) );
	vdp_comp_dff g4296 (.Q(w4288), .D(w4336), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_not g4297 (.nZ(w4346), .A(w4347) );
	vdp_not g4298 (.nZ(w4293), .A(w4348) );
	vdp_not g4299 (.nZ(w4335), .A(w4334) );
	vdp_nand g4300 (.Z(w4348), .B(w4335), .A(w4291) );
	vdp_not g4301 (.nZ(w4333), .A(w4337) );
	vdp_nand g4302 (.Z(w4340), .B(w4339), .A(w4338) );
	vdp_not g4303 (.nZ(w4312), .A(w4297) );
	vdp_nand g4304 (.Z(w4343), .B(w4342), .A(w4341) );
	vdp_not g4305 (.nZ(w4306), .A(w4311) );
	vdp_not g4306 (.nZ(RES), .A(w4308) );
	vdp_dff g4307 (.Q(w4291), .R(1'b0), .D(w4336), .C(w4309) );
	vdp_dff g4308 (.Q(w4334), .R(1'b0), .D(w4291), .C(w4309) );
	vdp_dff g4309 (.Q(w4347), .R(w4293), .D(w4337), .C(w4309) );
	vdp_dff g4310 (.Q(w4337), .R(w4293), .D(w4346), .C(w4309) );
	vdp_dff g4311 (.Q(w4338), .R(w4293), .D(w4297), .C(w4309) );
	vdp_dff g4312 (.Q(w4339), .R(w4293), .D(w4338), .C(w4309) );
	vdp_dff g4313 (.Q(w4297), .R(w4293), .D(w4340), .C(w4309) );
	vdp_dff g4314 (.Q(w4341), .R(w4293), .D(w4311), .C(w4309) );
	vdp_dff g4315 (.Q(w4342), .R(w4293), .D(w4341), .C(w4309) );
	vdp_dff g4316 (.Q(w4344), .R(w4293), .D(w4343), .C(w4309) );
	vdp_dff g4317 (.Q(w4311), .R(w4293), .D(w4344), .C(w4309) );
	vdp_not g4318 (.nZ(w4332), .A(w4333) );
	vdp_nand g4319 (.Z(w4336), .B(w1374), .A(w4349) );
	vdp_not g4320 (.nZ(M68K_CPU_CLOCK), .A(w4305) );
	vdp_or g4321 (.Z(w4328), .B(w40), .A(RS0) );
	vdp_aon22 g4322 (.Z(w4298), .B1(w4326), .A1(w4327), .B2(PAL), .A2(w4307) );
	vdp_or g4323 (.Z(w4305), .B(w4314), .A(w4306) );
	vdp_comp_we g4324 (.A(w2545), .nZ(nHCLK2), .Z(HCLK2) );
	vdp_comp_we g4325 (.A(w2544), .nZ(nHCLK1), .Z(HCLK1) );
	vdp_comp_we g4326 (.A(w4359), .nZ(nDCLK2), .Z(DCLK2) );
	vdp_comp_we g4327 (.A(EDCLK_O), .nZ(nDCLK1), .Z(DCLK1) );
	vdp_not g4328 (.nZ(w4359), .A(EDCLK_O) );
	vdp_sr_bit g4329 (.Q(w4453), .D(w4452), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4330 (.Q(w4471), .D(w4448), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4331 (.Q(w4448), .D(w4432), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4332 (.Q(w4432), .D(w4425), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4333 (.Q(w4428), .D(w6284), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4334 (.Q(w6284), .D(w6285), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4335 (.Q(w6285), .D(w6287), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4336 (.Q(w6287), .D(w6286), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4337 (.Q(w6286), .D(w6288), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4338 (.Q(w6288), .D(w6289), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4339 (.Q(w6289), .D(w6291), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4340 (.Q(w6291), .D(w6290), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4341 (.Q(w6290), .D(w6163), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4342 (.Q(w6163), .D(w4374), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4343 (.Q(w4410), .D(w4411), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4344 (.Q(w4411), .D(w23), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4345 (.Q(w4667), .D(w6292), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4346 (.Q(w4379), .D(w4701), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4347 (.Q(w4378), .D(w6280), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4348 (.Q(w6027), .D(w4455), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4349 (.Q(w4454), .D(w6293), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4350 (.Q(w4456), .D(w4446), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4351 (.Q(w6282), .D(w4), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4352 (.Q(w4398), .D(w4418), .nC(w4421), .C(w4422) );
	vdp_slatch g4353 (.Q(w4403), .D(w4419), .nC(w4421), .C(w4422) );
	vdp_slatch g4354 (.Q(w4390), .D(w4420), .nC(w4421), .C(w4422) );
	vdp_slatch g4355 (.Q(w4382), .D(w4426), .nC(w4421), .C(w4422) );
	vdp_slatch g4356 (.Q(w4381), .D(w4417), .nC(w4421), .C(w4422) );
	vdp_slatch g4357 (.Q(w4380), .D(w4416), .nC(w4421), .C(w4422) );
	vdp_slatch g4358 (.Q(w4430), .D(w4415), .nC(w4421), .C(w4422) );
	vdp_slatch g4359 (.Q(w4383), .D(w4413), .nC(w4421), .C(w4422) );
	vdp_slatch g4360 (.Q(w4386), .D(w4414), .nC(w4421), .C(w4422) );
	vdp_slatch g4361 (.Q(w4387), .D(w4412), .nC(w4421), .C(w4422) );
	vdp_comp_str g4362 (.nZ(w4421), .A(w4427), .Z(w4422) );
	vdp_sr_bit g4363 (.Q(w4449), .D(w4472), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4364 (.Q(w6013), .D(w35), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_xor g4365 (.Z(w4396), .B(w4388), .A(w4399) );
	vdp_xor g4366 (.Z(w4391), .B(w4389), .A(w4397) );
	vdp_xor g4367 (.Z(w4393), .B(w4376), .A(w4390) );
	vdp_xor g4368 (.Z(w6114), .B(w4376), .A(w4382) );
	vdp_xor g4369 (.Z(w6115), .B(w4376), .A(w4381) );
	vdp_xor g4370 (.Z(w6110), .B(w4376), .A(w4380) );
	vdp_aon22 g4371 (.Z(w6111), .B2(w4404), .B1(w4398), .A1(w4396), .A2(w4392) );
	vdp_aon22 g4372 (.Z(w6112), .B2(w4404), .B1(w4396), .A1(w4391), .A2(w4392) );
	vdp_aon22 g4373 (.Z(w6113), .B2(w4404), .B1(w4391), .A1(w4393), .A2(w4392) );
	vdp_aon22 g4374 (.Z(w4394), .B2(w4385), .B1(w4390), .A1(w4403), .A2(w4395) );
	vdp_aon22 g4375 (.Z(w4400), .B2(w4385), .B1(w4403), .A1(w4398), .A2(w4395) );
	vdp_aon22 g4376 (.Z(w4464), .B2(w4457), .B1(w4460), .A1(w4461), .A2(w69) );
	vdp_aon22 g4377 (.Z(w4465), .B2(w4459), .B1(w4460), .A1(w4461), .A2(w68) );
	vdp_aon22 g4378 (.Z(w4466), .B2(w4458), .B1(w4460), .A1(w4461), .A2(w67) );
	vdp_aon22 g4379 (.Z(w4467), .B2(w4462), .B1(w4460), .A1(w4461), .A2(w66) );
	vdp_aon22 g4380 (.Z(w4468), .B2(w4463), .B1(w4460), .A1(w4461), .A2(w65) );
	vdp_not g4381 (.nZ(w4433), .A(w4374) );
	vdp_not g4382 (.nZ(w4407), .A(w4437) );
	vdp_not g4383 (.nZ(w4436), .A(w108) );
	vdp_not g4384 (.nZ(w4442), .A(w4440) );
	vdp_not g4385 (.nZ(w4429), .A(M5) );
	vdp_not g4386 (.nZ(w4470), .A(w70) );
	vdp_not g4387 (.nZ(w4469), .A(w71) );
	vdp_not g4388 (.nZ(w4444), .A(1'b0) );
	vdp_not g4389 (.nZ(w4445), .A(M5) );
	vdp_not g4390 (.nZ(w4373), .A(w4374) );
	vdp_not g4391 (.nZ(w4377), .A(w4408) );
	vdp_not g4392 (.nZ(w4384), .A(w4387) );
	vdp_not g4393 (.nZ(w4389), .A(w4424) );
	vdp_and g4394 (.Z(w4425), .B(w4433), .A(w4434) );
	vdp_and g4395 (.Z(w4438), .B(w4436), .A(w4448) );
	vdp_or g4396 (.Z(w4435), .B(w4438), .A(w4451) );
	vdp_or g4397 (.Z(w4431), .B(w4474), .A(w4438) );
	vdp_and g4398 (.Z(w4450), .B(w4443), .A(1'b0) );
	vdp_and g4399 (.Z(w4473), .B(w4443), .A(w4444) );
	vdp_or g4400 (.Z(w4472), .B(w35), .A(w34) );
	vdp_and g4401 (.Z(SPRITE_OVF), .B(w6425), .A(w4) );
	vdp_and g4402 (.Z(w6280), .B(w4373), .A(w4375) );
	vdp_or g4403 (.Z(w4423), .B(w4379), .A(w4378) );
	vdp_and g4404 (.Z(w4388), .B(w4383), .A(w4376) );
	vdp_comp_we g4405 (.nZ(w4385), .A(w1), .Z(w4395) );
	vdp_comp_we g4406 (.nZ(w4404), .A(w1), .Z(w4392) );
	vdp_comp_we g4407 (.nZ(w4460), .A(w108), .Z(w4461) );
	vdp_not g4408 (.nZ(w4475), .A(w4452) );
	vdp_rs_ff g4409 (.Q(w6281), .R(w6282), .S(w4423) );
	vdp_rs_ff g4410 (.Q(w6425), .R(w6282), .S(w4378) );
	vdp_ha g4411 (.SUM(w4399), .B(w4400), .A(w4401) );
	vdp_ha g4412 (.SUM(w4397), .B(w4394), .A(w4402), .CO(w4401) );
	vdp_not g4413 (.nZ(w4409), .A(w4372) );
	vdp_and g4414 (.Z(w6279), .B(w4374), .A(w4375) );
	vdp_and3 g4415 (.Z(w4402), .B(w4383), .A(w4376), .C(w4384) );
	vdp_and3 g4416 (.Z(w4455), .B(w4453), .A(M5), .C(w4475) );
	vdp_and3 g4417 (.Z(w6293), .B(w4458), .A(w4457), .C(w4456) );
	vdp_and3 g4418 (.Z(w4474), .B(w71), .A(w4470), .C(w107) );
	vdp_and3 g4419 (.Z(w6283), .B(w70), .A(w4469), .C(w107) );
	vdp_and3 g4420 (.Z(w4451), .B(w4470), .A(w4469), .C(w107) );
	vdp_or3 g4421 (.Z(w4439), .B(w6283), .A(w4438), .C(w4442) );
	vdp_and3 g4422 (.Z(w4427), .B(HCLK1), .A(w4410), .C(DCLK1) );
	vdp_or3 g4423 (.Z(w4443), .B(w4446), .A(w4471), .C(w4445) );
	vdp_oai21 g4424 (.Z(w4424), .B(w4376), .A1(w4383), .A2(w4387) );
	vdp_nor g4425 (.Z(w4372), .B(w6279), .A(w4411) );
	vdp_nor g4426 (.Z(w6292), .B(w4377), .A(w6281) );
	vdp_nand g4427 (.Z(w4447), .B(w4429), .A(w4428) );
	vdp_nand g4428 (.Z(w4406), .B(w4470), .A(w4469) );
	vdp_nand g4429 (.Z(w4437), .B(w70), .A(w4469) );
	vdp_nand g4430 (.Z(w4405), .B(w71), .A(w4470) );
	vdp_nor g4431 (.Z(w4452), .B(w4454), .A(w4370) );
	vdp_cnt_bit_rev g4432 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4457), .CI(w4479), .B(w4449), .A(w4450) );
	vdp_cnt_bit_rev g4433 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4459), .CI(w4478), .B(w4449), .A(w4450), .CO(w4479) );
	vdp_cnt_bit_rev g4434 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4458), .CI(w4477), .B(w4449), .A(w4450), .CO(w4478) );
	vdp_cnt_bit_rev g4435 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4462), .CI(w4476), .B(w4449), .A(w4450), .CO(w4477) );
	vdp_cnt_bit_rev g4436 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4463), .CI(w4473), .B(w4449), .A(w4450), .CO(w4476) );
	vdp_cnt_bit_load g4437 (.Q(w4486), .D(w4526), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4488), .CI(w6327), .L(w4527), .nL(w4492) );
	vdp_cnt_bit_load g4438 (.Q(w4489), .D(w4531), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4488), .CI(w6326), .L(w4527), .nL(w4492), .CO(w6327) );
	vdp_cnt_bit_load g4439 (.Q(w4491), .D(w4532), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4488), .CI(w6325), .L(w4527), .nL(w4492), .CO(w6326) );
	vdp_cnt_bit_load g4440 (.Q(w4493), .D(w4556), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4488), .CI(w6324), .L(w4527), .nL(w4492), .CO(w6325) );
	vdp_cnt_bit_load g4441 (.Q(w4497), .D(w4557), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4488), .CI(w6323), .L(w4527), .nL(w4492), .CO(w6324) );
	vdp_cnt_bit_load g4442 (.Q(w4494), .D(w4558), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4488), .CI(w6322), .L(w4527), .nL(w4492), .CO(w6323) );
	vdp_cnt_bit_load g4443 (.Q(w4490), .D(w4559), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4488), .CI(w4487), .L(w4527), .nL(w4492), .CO(w6322) );
	vdp_fa g4444 (.SUM(w4634), .CO(w6337), .CI(1'b1), .A(w4689), .B(w4637) );
	vdp_fa g4445 (.SUM(w4636), .CO(w6338), .CI(w6337), .A(w4688), .B(w4641) );
	vdp_fa g4446 (.SUM(w4642), .CO(w6339), .CI(w6338), .A(w4687), .B(w4645) );
	vdp_fa g4447 (.SUM(w4644), .CO(w6340), .CI(w6339), .A(w4686), .B(w4647) );
	vdp_fa g4448 (.SUM(w4649), .CO(w6341), .CI(w6340), .A(w4685), .B(w4651) );
	vdp_fa g4449 (.SUM(w4655), .CO(w6342), .CI(w6341), .A(w4684), .B(w4680) );
	vdp_fa g4450 (.SUM(w4658), .CO(w6343), .CI(w6342), .A(w4682), .B(w4657) );
	vdp_fa g4451 (.SUM(w4662), .CO(w6344), .CI(w6343), .A(w4694), .B(w4661) );
	vdp_fa g4452 (.SUM(w4664), .CO(w6345), .CI(w6344), .A(w4695), .B(w4663) );
	vdp_fa g4453 (.SUM(w4678), .CI(w6345), .A(w4699), .B(w4677) );
	vdp_fa g4454 (.SUM(w4689), .CO(w6328), .CI(1'b0), .A(VPOS[0]), .B(w4690) );
	vdp_fa g4455 (.SUM(w4688), .CO(w6329), .CI(w6328), .A(VPOS[1]), .B(w1) );
	vdp_fa g4456 (.SUM(w4687), .CO(w6330), .CI(w6329), .A(VPOS[2]), .B(1'b0) );
	vdp_fa g4457 (.SUM(w4686), .CO(w6331), .CI(w6330), .A(VPOS[3]), .B(1'b0) );
	vdp_fa g4458 (.SUM(w4685), .CO(w6332), .CI(w6331), .A(VPOS[4]), .B(1'b0) );
	vdp_fa g4459 (.SUM(w4684), .CO(w6333), .CI(w6332), .A(VPOS[5]), .B(1'b0) );
	vdp_fa g4460 (.SUM(w4682), .CO(w6334), .CI(w6333), .A(VPOS[6]), .B(1'b0) );
	vdp_fa g4461 (.SUM(w4694), .CO(w6335), .CI(w6334), .A(VPOS[7]), .B(w4690) );
	vdp_fa g4462 (.SUM(w4695), .CO(w6336), .CI(w6335), .A(VPOS[8]), .B(w1) );
	vdp_fa g4463 (.SUM(w4699), .CI(w6336), .A(VPOS[9]), .B(1'b0) );
	vdp_slatch g4464 (.nC(w4582), .C(w4581), .Q(w4627), .D(S[0]) );
	vdp_dlatch_inv g4465 (.nQ(w4626), .D(w4595), .nC(nHCLK2), .C(HCLK2) );
	vdp_slatch g4466 (.nC(w4567), .C(w4566), .Q(w4595), .D(w4584) );
	vdp_slatch g4467 (.nC(w4582), .C(w4581), .Q(w4624), .D(S[1]) );
	vdp_slatch g4468 (.nC(w4567), .C(w4566), .Q(w6367), .D(w4586) );
	vdp_slatch g4469 (.nC(w4582), .C(w4581), .Q(w4622), .D(S[2]) );
	vdp_slatch g4470 (.nC(w4567), .C(w4566), .Q(w6368), .D(w4577) );
	vdp_slatch g4471 (.nC(w4582), .C(w4581), .Q(w4620), .D(S[3]) );
	vdp_slatch g4472 (.nC(w4567), .C(w4566), .Q(w6369), .D(w4573) );
	vdp_slatch g4473 (.nC(w4582), .C(w4581), .Q(w4617), .D(S[4]) );
	vdp_slatch g4474 (.nC(w4567), .C(w4566), .Q(w6370), .D(w4569) );
	vdp_slatch g4475 (.nC(w4582), .C(w4581), .Q(w4616), .D(S[5]) );
	vdp_slatch g4476 (.nC(w4567), .C(w4566), .Q(w6371), .D(w4565) );
	vdp_slatch g4477 (.nC(w4582), .C(w4581), .Q(w4613), .D(S[6]) );
	vdp_slatch g4478 (.nC(w4567), .C(w4566), .Q(w6372), .D(w6314) );
	vdp_slatch g4479 (.nC(w4582), .C(w4581), .Q(w6373), .D(S[7]) );
	vdp_slatch g4480 (.nC(w4567), .C(w4566), .Q(w6374), .D(w4597) );
	vdp_slatch g4481 (.nC(w4567), .C(w4566), .Q(w4598), .D(w4599) );
	vdp_slatch g4482 (.nC(w4567), .C(w4566), .Q(w6375), .D(w4601) );
	vdp_dlatch_inv g4483 (.nQ(w4623), .D(w6367), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4484 (.nQ(w4621), .D(w6368), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4485 (.nQ(w4619), .D(w6369), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4486 (.nQ(w4618), .D(w6370), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4487 (.nQ(w4615), .D(w6371), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4488 (.nQ(w4612), .D(w6372), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4489 (.nQ(w4611), .D(w6374), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4490 (.nQ(w4610), .D(w4598), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4491 (.nQ(w4600), .D(w6375), .nC(nHCLK2), .C(HCLK2) );
	vdp_sr_bit g4492 (.Q(w4552), .D(w4483), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4493 (.Z(w4408), .B2(w4548), .B1(w4554), .A1(M5), .A2(w4553) );
	vdp_sr_bit g4494 (.Q(w4483), .D(w4549), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4495 (.Q(w4549), .D(w4550), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4496 (.Q(w4550), .D(w4528), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4497 (.Q(w4589), .D(w4591), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4498 (.Q(w4580), .D(w4594), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4499 (.Q(w4576), .D(w4587), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4500 (.Q(w4572), .D(w4588), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4501 (.Q(w4568), .D(w4570), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4502 (.Q(w4564), .D(w4562), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4503 (.Q(w4596), .D(w4563), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4504 (.Q(w6376), .D(w4561), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4505 (.Q(w4510), .D(w4560), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4506 (.Q(w4517), .D(w4555), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4507 (.Q(w4551), .D(w4484), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4508 (.Q(w4484), .D(w4506), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4509 (.Q(w4736), .D(w116), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4510 (.Q(w4738), .D(VRAMA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4511 (.Q(w4506), .D(w8), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4512 (.Q(w4739), .D(w6321), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4513 (.Q(w6321), .D(w4736), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4514 (.Q(w6365), .D(w4722), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4515 (.Q(w6363), .D(w4725), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4516 (.Q(w6361), .D(w4741), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4517 (.Q(w6359), .D(w4702), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4518 (.Q(w6357), .D(w4526), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4519 (.Q(w6355), .D(w4531), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4520 (.Q(w6353), .D(w4532), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4521 (.Q(w6351), .D(w4556), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4522 (.Q(w6349), .D(w4557), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4523 (.Q(w6347), .D(w4558), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4524 (.Q(w4720), .D(w4559), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4525 (.Q(w4712), .D(w6346), .nC(w4711), .C(w4703) );
	vdp_dlatch_inv g4526 (.nQ(w6346), .D(w4720), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4527 (.Q(w4713), .D(w6348), .nC(w4711), .C(w4703) );
	vdp_dlatch_inv g4528 (.nQ(w6348), .D(w6347), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4529 (.Q(w4714), .D(w6350), .nC(w4711), .C(w4703) );
	vdp_dlatch_inv g4530 (.nQ(w6350), .D(w6349), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4531 (.Q(w4715), .D(w6352), .nC(w4711), .C(w4703) );
	vdp_dlatch_inv g4532 (.nQ(w6352), .D(w6351), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4533 (.Q(w4716), .D(w6354), .nC(w4711), .C(w4703) );
	vdp_dlatch_inv g4534 (.nQ(w6354), .D(w6353), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4535 (.Q(w6320), .D(w6356), .nC(w4711), .C(w4703) );
	vdp_dlatch_inv g4536 (.nQ(w6356), .D(w6355), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4537 (.Q(w4717), .D(w6358), .nC(w4711), .C(w4703) );
	vdp_dlatch_inv g4538 (.nQ(w6358), .D(w6357), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4539 (.Q(w4707), .D(w6360), .nC(w4711), .C(w4703) );
	vdp_dlatch_inv g4540 (.nQ(w6360), .D(w6359), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4541 (.Q(w4710), .D(w6362), .nC(w4711), .C(w4703) );
	vdp_dlatch_inv g4542 (.nQ(w6362), .D(w6361), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4543 (.Q(w4708), .D(w6364), .nC(w4711), .C(w4703) );
	vdp_dlatch_inv g4544 (.nQ(w6364), .D(w6363), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4545 (.Q(w4709), .D(w6366), .nC(w4711), .C(w4703) );
	vdp_dlatch_inv g4546 (.nQ(w6366), .D(w6365), .nC(nHCLK1), .C(HCLK1) );
	vdp_aon22 g4547 (.Z(w6181), .B2(w4536), .B1(w4486), .A1(w4485), .A2(w6161) );
	vdp_aon22 g4548 (.Z(w6182), .B2(w4536), .B1(w4489), .A1(w4485), .A2(w4541) );
	vdp_aon22 g4549 (.Z(w6183), .B2(w4536), .B1(w4491), .A1(w4485), .A2(w4540) );
	vdp_aon22 g4550 (.Z(w6184), .B2(w4536), .B1(w4493), .A1(w4485), .A2(w4539) );
	vdp_aon22 g4551 (.Z(w6185), .B2(w4536), .B1(w4497), .A1(w4485), .A2(w4538) );
	vdp_aon22 g4552 (.Z(w6187), .B2(w4536), .B1(w4494), .A1(w4485), .A2(w4537) );
	vdp_aon22 g4553 (.Z(w6186), .B2(w4536), .B1(w4490), .A1(w4485), .A2(w4535) );
	vdp_aon22 g4554 (.Z(w4752), .B2(w4499), .B1(w3), .A1(w4495), .A2(w4490) );
	vdp_aon22 g4555 (.Z(w4648), .B2(w4608), .B1(w4617), .A1(w4618), .A2(w4632) );
	vdp_2x_sr_bit g4556 (.Q(w4547), .D(w4490), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4557 (.Z(w6162), .B2(w4499), .B1(w4547), .A1(w4495), .A2(w4494) );
	vdp_2x_sr_bit g4558 (.Q(w4496), .D(w4494), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4559 (.Z(w4805), .B2(w4499), .B1(w4496), .A1(w4495), .A2(w4497) );
	vdp_2x_sr_bit g4560 (.Q(w4534), .D(w4497), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4561 (.Z(w4811), .B2(w4499), .B1(w4534), .A1(w4495), .A2(w4493) );
	vdp_2x_sr_bit g4562 (.Q(w4498), .D(w4493), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4563 (.Z(w4860), .B2(w4499), .B1(w4498), .A1(w4495), .A2(w4491) );
	vdp_2x_sr_bit g4564 (.Q(w4501), .D(w4491), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4565 (.Z(w4911), .B2(w4499), .B1(w4501), .A1(w4495), .A2(w4489) );
	vdp_aon22 g4566 (.Z(w4925), .B2(w4499), .B1(1'b1), .A1(w4495), .A2(w4486) );
	vdp_aon22 g4567 (.Z(w4584), .B2(w4509), .B1(w4585), .A1(w4512), .A2(w4583) );
	vdp_dlatch_inv g4568 (.nQ(w4583), .D(w4589), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4569 (.nZ(w4585), .A(S[0]) );
	vdp_aon22 g4570 (.Z(w4586), .B2(w4509), .B1(w4579), .A1(w4512), .A2(w4578) );
	vdp_dlatch_inv g4571 (.nQ(w4578), .D(w4580), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4572 (.nZ(w4579), .A(S[1]) );
	vdp_aon22 g4573 (.Z(w4577), .B2(w4509), .B1(w4575), .A1(w4512), .A2(w4574) );
	vdp_dlatch_inv g4574 (.nQ(w4574), .D(w4576), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4575 (.nZ(w4575), .A(S[2]) );
	vdp_aon22 g4576 (.Z(w4573), .B2(w4509), .B1(w4533), .A1(w4512), .A2(w4571) );
	vdp_dlatch_inv g4577 (.nQ(w4571), .D(w4572), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4578 (.nZ(w4533), .A(S[3]) );
	vdp_aon22 g4579 (.Z(w4569), .B2(w4509), .B1(w4529), .A1(w4512), .A2(w4530) );
	vdp_dlatch_inv g4580 (.nQ(w4530), .D(w4568), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4581 (.nZ(w4529), .A(S[4]) );
	vdp_aon22 g4582 (.Z(w4565), .B2(w4509), .B1(w4525), .A1(w4512), .A2(w4524) );
	vdp_dlatch_inv g4583 (.nQ(w4524), .D(w4564), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4584 (.nZ(w4525), .A(S[5]) );
	vdp_aon22 g4585 (.Z(w6314), .B2(w4509), .B1(w4520), .A1(w4512), .A2(w4519) );
	vdp_dlatch_inv g4586 (.nQ(w4519), .D(w4596), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4587 (.nZ(w4520), .A(S[6]) );
	vdp_aon22 g4588 (.Z(w4597), .B2(w4509), .B1(w4513), .A1(w4512), .A2(w4511) );
	vdp_dlatch_inv g4589 (.nQ(w4511), .D(w6376), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4590 (.nZ(w4513), .A(S[7]) );
	vdp_aon22 g4591 (.Z(w4599), .B2(w4509), .B1(w4747), .A1(w4512), .A2(1'b1) );
	vdp_dlatch_inv g4592 (.nQ(w4747), .D(w4510), .nC(nHCLK1), .C(HCLK1) );
	vdp_aon22 g4593 (.Z(w4601), .B2(w4509), .B1(1'b1), .A1(w4512), .A2(w4518) );
	vdp_dlatch_inv g4594 (.nQ(w4518), .D(w4517), .nC(nHCLK1), .C(HCLK1) );
	vdp_sr_bit g4595 (.Q(w4488), .D(w6310), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4596 (.Q(w4500), .D(w28), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4597 (.Q(w4521), .D(w4500), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4598 (.Q(w4505), .D(w5), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4599 (.Q(w4515), .D(w4505), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4600 (.Q(w4528), .D(w6309), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_not g4601 (.nZ(w4523), .A(w4522) );
	vdp_not g4602 (.nZ(w4516), .A(M5) );
	vdp_not g4603 (.nZ(w6310), .A(w4514) );
	vdp_not g4604 (.nZ(w4504), .A(w4515) );
	vdp_not g4605 (.nZ(w6309), .A(w4507) );
	vdp_not g4606 (.nZ(w4502), .A(w4487) );
	vdp_aon22 g4607 (.Z(w4607), .B2(w4603), .B1(w4420), .A1(w4602), .A2(w4419) );
	vdp_aon22 g4608 (.Z(w4606), .B2(w4603), .B1(w4419), .A1(w4602), .A2(w4418) );
	vdp_aon22 g4609 (.Z(w4605), .B2(w4603), .B1(w4418), .A1(w4602), .A2(1'b0) );
	vdp_slatch g4610 (.nQ(w6385), .D(w4735), .nC(w4719), .C(w4724) );
	vdp_aon22 g4611 (.Z(w4735), .B2(w4718), .B1(w4591), .A1(w4723), .A2(w4559) );
	vdp_notif0 g4612 (.A(w6385), .nZ(AD_DATA[0]), .nE(w4729) );
	vdp_slatch g4613 (.nQ(w6384), .D(w4734), .nC(w4719), .C(w4724) );
	vdp_aon22 g4614 (.Z(w4734), .B2(w4718), .B1(w4594), .A1(w4723), .A2(w4558) );
	vdp_notif0 g4615 (.A(w6384), .nZ(AD_DATA[1]), .nE(w4729) );
	vdp_slatch g4616 (.nQ(w6383), .D(w4733), .nC(w4719), .C(w4724) );
	vdp_aon22 g4617 (.Z(w4733), .B2(w4718), .B1(w4587), .A1(w4723), .A2(w4557) );
	vdp_notif0 g4618 (.A(w6383), .nZ(AD_DATA[2]), .nE(w4729) );
	vdp_slatch g4619 (.nQ(w6382), .D(w6318), .nC(w4719), .C(w4724) );
	vdp_aon22 g4620 (.Z(w6318), .B2(w4718), .B1(w4588), .A1(w4723), .A2(w4556) );
	vdp_notif0 g4621 (.A(w6382), .nZ(AD_DATA[3]), .nE(w4729) );
	vdp_slatch g4622 (.nQ(w6381), .D(w6317), .nC(w4719), .C(w4724) );
	vdp_aon22 g4623 (.Z(w6317), .B2(w4718), .B1(w4570), .A1(w4723), .A2(w4532) );
	vdp_notif0 g4624 (.A(w6381), .nZ(AD_DATA[4]), .nE(w4729) );
	vdp_slatch g4625 (.nQ(w6380), .D(w6316), .nC(w4719), .C(w4724) );
	vdp_aon22 g4626 (.Z(w6316), .B2(w4718), .B1(w4562), .A1(w4723), .A2(w4531) );
	vdp_notif0 g4627 (.A(w6380), .nZ(AD_DATA[5]), .nE(w4729) );
	vdp_slatch g4628 (.nQ(w6379), .D(w4732), .nC(w4719), .C(w4724) );
	vdp_aon22 g4629 (.Z(w4732), .B2(w4718), .B1(w4563), .A1(w4723), .A2(w4526) );
	vdp_notif0 g4630 (.A(w6379), .nZ(AD_DATA[6]), .nE(w4729) );
	vdp_slatch g4631 (.nQ(w6378), .D(w4740), .nC(w4719), .C(w4724) );
	vdp_aon22 g4632 (.Z(w4740), .B2(w4718), .B1(w4561), .A1(w4723), .A2(w4702) );
	vdp_notif0 g4633 (.A(w6378), .nZ(AD_DATA[7]), .nE(w4729) );
	vdp_slatch g4634 (.nQ(w4731), .D(w4730), .nC(w4719), .C(w4724) );
	vdp_aon22 g4635 (.Z(w4730), .B2(w4718), .B1(w4560), .A1(w4723), .A2(w4741) );
	vdp_notif0 g4636 (.A(w4731), .nZ(RD_DATA[0]), .nE(w4729) );
	vdp_slatch g4637 (.nQ(w4728), .D(w4727), .nC(w4719), .C(w4724) );
	vdp_aon22 g4638 (.Z(w4727), .B2(w4718), .B1(w4555), .A1(w4723), .A2(w4725) );
	vdp_notif0 g4639 (.A(w4728), .nZ(RD_DATA[1]), .nE(w4729) );
	vdp_slatch g4640 (.nQ(w4726), .D(w4721), .nC(w4719), .C(w4724) );
	vdp_aon22 g4641 (.Z(w4721), .B2(w4718), .B1(1'b0), .A1(w4723), .A2(w4722) );
	vdp_notif0 g4642 (.A(w4726), .nZ(RD_DATA[2]), .nE(w4729) );
	vdp_not g4643 (.nZ(w4729), .A(w4739) );
	vdp_sr_bit g4644 (.Q(w4413), .D(w6389), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4645 (.Q(w4414), .D(w4697), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4646 (.Q(w4693), .D(w4691), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_dlatch_inv g4647 (.nQ(w4692), .D(w4593), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4648 (.nQ(w4691), .D(w4631), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g4649 (.nQ(w4637), .D(w4633), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4650 (.nQ(w6315), .D(w4634), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4651 (.nQ(w4641), .D(w4635), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4652 (.nQ(w4639), .D(w4636), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4653 (.nQ(w4645), .D(w4640), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4654 (.nQ(w4643), .D(w4642), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4655 (.nQ(w4647), .D(w4646), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4656 (.nQ(w4656), .D(w4644), .nC(nHCLK2), .C(HCLK2) );
	vdp_aon22 g4657 (.Z(w4646), .B2(w4608), .B1(w4620), .A1(w4619), .A2(w4632) );
	vdp_aon22 g4658 (.Z(w4640), .B2(w4608), .B1(w4622), .A1(w4621), .A2(w4632) );
	vdp_aon22 g4659 (.Z(w4635), .B2(w4608), .B1(w4624), .A1(w4623), .A2(w4632) );
	vdp_aon22 g4660 (.Z(w4633), .B2(w4608), .B1(w4627), .A1(w4626), .A2(w4632) );
	vdp_not g4661 (.nZ(w4630), .A(w4593) );
	vdp_not g4662 (.nZ(w4416), .A(w6315) );
	vdp_not g4663 (.nZ(w4417), .A(w4639) );
	vdp_not g4664 (.nZ(w4426), .A(w4643) );
	vdp_not g4665 (.nZ(w4420), .A(w4656) );
	vdp_not g4666 (.nZ(w4652), .A(w4648) );
	vdp_not g4667 (.nZ(w4419), .A(w4650) );
	vdp_dlatch_inv g4668 (.nQ(w4651), .D(w4648), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4669 (.nQ(w4650), .D(w4649), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g4670 (.nZ(w4418), .A(w4659) );
	vdp_dlatch_inv g4671 (.nQ(w4680), .D(w4614), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4672 (.nQ(w4659), .D(w4655), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g4673 (.nZ(w4660), .A(w4681) );
	vdp_dlatch_inv g4674 (.nQ(w4657), .D(w4681), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4675 (.nQ(w4670), .D(w4658), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g4676 (.nZ(w4654), .A(w4665) );
	vdp_dlatch_inv g4677 (.nQ(w4661), .D(w4665), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4678 (.nQ(w4671), .D(w4662), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4679 (.nQ(w4663), .D(w4653), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4680 (.nQ(w4668), .D(w4664), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4681 (.nQ(w4677), .D(w4666), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4682 (.nQ(w4679), .D(w4678), .nC(nHCLK2), .C(HCLK2) );
	vdp_sr_bit g4683 (.Q(w4412), .D(w6377), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4684 (.Z(w4666), .B2(w4608), .B1(1'b0), .A1(w4600), .A2(w4632) );
	vdp_aon22 g4685 (.Z(w4653), .B2(w4608), .B1(1'b0), .A1(w4610), .A2(w4632) );
	vdp_aon22 g4686 (.Z(w6377), .B2(w4706), .B1(M5), .A1(w117), .A2(w4743) );
	vdp_not g4687 (.nZ(w4696), .A(w1) );
	vdp_not g4688 (.nZ(w4746), .A(w4709) );
	vdp_not g4689 (.nZ(w4697), .A(w4708) );
	vdp_not g4690 (.nZ(w4744), .A(w4710) );
	vdp_not g4691 (.nZ(w4706), .A(w4707) );
	vdp_not g4692 (.nZ(w4743), .A(M5) );
	vdp_not g4693 (.nZ(w4701), .A(w4704) );
	vdp_not g4694 (.nZ(w4698), .A(w4412) );
	vdp_not g4695 (.nZ(w6386), .A(w4413) );
	vdp_not g4696 (.nZ(w4745), .A(M5) );
	vdp_not g4697 (.nZ(w4669), .A(w1) );
	vdp_not g4698 (.nZ(w4673), .A(w4605) );
	vdp_bufif0 g4699 (.A(1'b0), .Z(VRAMA[0]), .nE(w4502) );
	vdp_bufif0 g4700 (.A(w4490), .Z(VRAMA[1]), .nE(w4502) );
	vdp_bufif0 g4701 (.A(w4494), .Z(VRAMA[2]), .nE(w4502) );
	vdp_bufif0 g4702 (.A(w4497), .Z(VRAMA[3]), .nE(w4502) );
	vdp_bufif0 g4703 (.A(w4493), .Z(VRAMA[4]), .nE(w4502) );
	vdp_bufif0 g4704 (.A(w4491), .Z(VRAMA[5]), .nE(w4502) );
	vdp_bufif0 g4705 (.A(1'b0), .Z(VRAMA[6]), .nE(w4502) );
	vdp_bufif0 g4706 (.A(1'b0), .Z(VRAMA[7]), .nE(w4502) );
	vdp_aon22 g4707 (.Z(w4665), .B2(w4608), .B1(w6373), .A1(w4611), .A2(w4632) );
	vdp_aon22 g4708 (.Z(w4681), .B2(w4608), .B1(w4613), .A1(w4612), .A2(w4632) );
	vdp_aon22 g4709 (.Z(w4614), .B2(w4608), .B1(w4616), .A1(w4615), .A2(w4632) );
	vdp_comp_str g4710 (.A(w4629), .nZ(w4567), .Z(w4566) );
	vdp_and g4711 (.Z(w4592), .B(w4552), .A(w4548) );
	vdp_comp_we g4712 (.A(w4592), .nZ(w4632), .Z(w4608) );
	vdp_comp_str g4713 (.A(w4625), .nZ(w4582), .Z(w4581) );
	vdp_not g4714 (.nZ(w4548), .A(M5) );
	vdp_comp_str g4715 (.A(w4700), .nZ(w4711), .Z(w4703) );
	vdp_comp_str g4716 (.A(w4737), .nZ(w4719), .Z(w4724) );
	vdp_comp_we g4717 (.A(M5), .nZ(w4509), .Z(w4512) );
	vdp_comp_we g4718 (.A(w4543), .nZ(w4536), .Z(w4485) );
	vdp_comp_we g4719 (.A(w4523), .nZ(w4492), .Z(w4527) );
	vdp_comp_we g4720 (.A(M5), .nZ(w4499), .Z(w4495) );
	vdp_comp_we g4721 (.A(w1), .nZ(w4603), .Z(w4602) );
	vdp_comp_we g4722 (.nZ(w4718), .A(w4738), .Z(w4723) );
	vdp_and g4723 (.Z(w4629), .B(w4691), .A(DCLK2) );
	vdp_and g4724 (.Z(w4625), .B(w4693), .A(DCLK2) );
	vdp_and g4725 (.Z(w4690), .B(M5), .A(w4696) );
	vdp_and g4726 (.Z(w6389), .B(w4744), .A(M5) );
	vdp_and g4727 (.Z(w6388), .B(w4698), .A(w4413) );
	vdp_and g4728 (.Z(w4737), .B(w4736), .A(HCLK1) );
	vdp_or g4729 (.Z(w4672), .B(w4669), .A(w4679) );
	vdp_or g4730 (.Z(w6390), .B(w4745), .A(w4668) );
	vdp_and g4731 (.Z(w4487), .B(w4516), .A(w4500) );
	vdp_and g4732 (.Z(w4544), .B(w4481), .A(w4546) );
	vdp_and g4733 (.Z(w6178), .B(w4546), .A(w4482) );
	vdp_and g4734 (.Z(w6179), .B(w4480), .A(w4482) );
	vdp_and g4735 (.Z(w6180), .B(w4481), .A(w4480) );
	vdp_and g4736 (.Z(w6154), .B(H40), .A(VRAMA[9]) );
	vdp_or g4737 (.Z(w4554), .B(w4483), .A(w4552) );
	vdp_or g4738 (.Z(w4553), .B(w4483), .A(w4549) );
	vdp_not g4739 (.nZ(w4480), .A(w4546) );
	vdp_oai21 g4740 (.Z(w4507), .B(w28), .A1(w29), .A2(w5) );
	vdp_oai21 g4741 (.Z(w4704), .B(w4408), .A1(w4628), .A2(w4705) );
	vdp_aoi22 g4742 (.Z(w4593), .B2(w4548), .B1(w4549), .A1(M5), .A2(w4590) );
	vdp_or3 g4743 (.Z(w4590), .B(w4549), .A(w4550), .C(w4551) );
	vdp_and3 g4744 (.Z(w4700), .B(DCLK1), .A(HCLK2), .C(w4692) );
	vdp_oai21 g4745 (.Z(w4522), .B(M5), .A1(w4500), .A2(w4521) );
	vdp_2a3oi g4746 (.Z(w4514), .B(w4505), .A1(w4504), .A2(w4), .C(SYSRES) );
	vdp_or8 g4747 (.Z(w4705), .B(w4717), .A(M5), .C(w6320), .D(w4716), .F(w4714), .E(w4715), .G(w4713), .H(w4712) );
	vdp_and9 g4748 (.Z(w4375), .B(w4674), .A(w4676), .C(w4675), .D(w4673), .F(w4671), .E(w4672), .G(w4670), .H(w4667), .I(w6390) );
	vdp_nor12 g4749 (.Z(w4628), .B(w4614), .A(1'b0), .C(w4654), .D(M5), .F(w4666), .E(w4653), .G(w4660), .H(w4652), .J(w4635), .I(w4640), .K(w4633), .L(w4646) );
	vdp_or4 g4750 (.Z(w4543), .B(w4482), .A(w4481), .C(w4542), .D(w4484) );
	vdp_nand g4751 (.Z(w4631), .B(w4630), .A(HCLK1) );
	vdp_nand g4752 (.Z(w4676), .B(w4607), .A(w6387) );
	vdp_nand g4753 (.Z(w4675), .B(w4606), .A(w6386) );
	vdp_nor g4754 (.Z(w6387), .B(w4412), .A(w4413) );
	vdp_nand3 g4755 (.Z(w4674), .B(w4606), .A(w6388), .C(w4607) );
	vdp_sr_bit g4756 (.Q(w4415), .D(w4746), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4757 (.Q(w4754), .D(w26), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4758 (.Q(w4434), .D(w6311), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4759 (.Q(w4753), .D(w6295), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4760 (.Q(w6295), .D(w6296), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4761 (.Q(w6296), .D(w4752), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4762 (.Z(w4757), .B2(w4753), .B1(w5105), .A1(DB[4]), .A2(w5106) );
	vdp_notif0 g4763 (.A(HPOS[1]), .nZ(VRAMA[1]), .nE(w4968) );
	vdp_aon22 g4764 (.Z(w6311), .B2(w4751), .B1(w4754), .A1(M5), .A2(w26) );
	vdp_not g4765 (.nZ(w4751), .A(M5) );
	vdp_lfsr_bit g4766 (.Q(w4758), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6562), .A1(w4757), .A2(w6563) );
	vdp_lfsr_bit g4767 (.Q(w4761), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6560), .A1(w4758), .A2(w6561) );
	vdp_lfsr_bit g4768 (.Q(w4763), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6558), .A1(w4761), .A2(w6559) );
	vdp_lfsr_bit g4769 (.Q(w4764), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6556), .A1(w4763), .A2(w6557) );
	vdp_lfsr_bit g4770 (.Q(w4768), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6554), .A1(w4764), .A2(w6555) );
	vdp_lfsr_bit g4771 (.Q(w4766), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6552), .A1(w4768), .A2(w6553) );
	vdp_lfsr_bit g4772 (.Q(w4770), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6550), .A1(w4766), .A2(w6551) );
	vdp_lfsr_bit g4773 (.Q(w4750), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6549), .A1(w4770), .A2(w6548) );
	vdp_lfsr_bit g4774 (.Q(w4774), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4948), .A1(w4750), .A2(w6547) );
	vdp_lfsr_bit g4775 (.Q(w4776), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5109), .A1(w4774), .A2(w5110) );
	vdp_lfsr_bit g4776 (.Q(w4780), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4994), .A1(w4776), .A2(w4995) );
	vdp_lfsr_bit g4777 (.Q(w4777), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4991), .A1(w4780), .A2(w4992) );
	vdp_lfsr_bit g4778 (.Q(w4779), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4989), .A1(w4777), .A2(w4990) );
	vdp_lfsr_bit g4779 (.Q(w4783), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6545), .A1(w4779), .A2(w6544) );
	vdp_lfsr_bit g4780 (.Q(w4784), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4986), .A1(w4783), .A2(w4987) );
	vdp_lfsr_bit g4781 (.Q(w4788), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6542), .A1(w4784), .A2(w6543) );
	vdp_lfsr_bit g4782 (.Q(w4787), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6546), .A1(w4788), .A2(w6616) );
	vdp_lfsr_bit g4783 (.Q(w4792), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4983), .A1(w4787), .A2(w4984) );
	vdp_lfsr_bit g4784 (.Q(w4794), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4982), .A1(w4792), .A2(w4981) );
	vdp_lfsr_bit g4785 (.Q(w4749), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4979), .A1(w4794), .A2(w4980) );
	vdp_bufif0 g4786 (.A(w4750), .Z(VRAMA[1]), .nE(w6313) );
	vdp_bufif0 g4787 (.A(1'b0), .Z(VRAMA[1]), .nE(w5002) );
	vdp_notif0 g4788 (.A(w4749), .nZ(DB[4]), .nE(w5111) );
	vdp_sr_bit g4789 (.Q(w4799), .D(w6298), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4790 (.Q(w6298), .D(w6297), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4791 (.Q(w6297), .D(w6162), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4792 (.Z(w4756), .B2(w4799), .B1(w5105), .A1(DB[5]), .A2(w5106) );
	vdp_notif0 g4793 (.A(w4807), .nZ(VRAMA[2]), .nE(w4968) );
	vdp_lfsr_bit g4794 (.Q(w4759), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6562), .A1(w4756), .A2(w6563) );
	vdp_lfsr_bit g4795 (.Q(w4760), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6560), .A1(w4759), .A2(w6561) );
	vdp_lfsr_bit g4796 (.Q(w4762), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6558), .A1(w4760), .A2(w6559) );
	vdp_lfsr_bit g4797 (.Q(w4765), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6556), .A1(w4762), .A2(w6557) );
	vdp_lfsr_bit g4798 (.Q(w4769), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6554), .A1(w4765), .A2(w6555) );
	vdp_lfsr_bit g4799 (.Q(w4767), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6552), .A1(w4769), .A2(w6553) );
	vdp_lfsr_bit g4800 (.Q(w4771), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6550), .A1(w4767), .A2(w6551) );
	vdp_lfsr_bit g4801 (.Q(w4772), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6549), .A1(w4771), .A2(w6548) );
	vdp_lfsr_bit g4802 (.Q(w4775), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4948), .A1(w4772), .A2(w6547) );
	vdp_lfsr_bit g4803 (.Q(w4773), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5109), .A1(w4775), .A2(w5110) );
	vdp_lfsr_bit g4804 (.Q(w4781), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4994), .A1(w4773), .A2(w4995) );
	vdp_lfsr_bit g4805 (.Q(w4778), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4991), .A1(w4781), .A2(w4992) );
	vdp_lfsr_bit g4806 (.Q(w4782), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4989), .A1(w4778), .A2(w4990) );
	vdp_lfsr_bit g4807 (.Q(w4786), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6545), .A1(w4782), .A2(w6544) );
	vdp_lfsr_bit g4808 (.Q(w4785), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4986), .A1(w4786), .A2(w4987) );
	vdp_lfsr_bit g4809 (.Q(w4789), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6542), .A1(w4785), .A2(w6543) );
	vdp_lfsr_bit g4810 (.Q(w4790), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6546), .A1(w4789), .A2(w6616) );
	vdp_lfsr_bit g4811 (.Q(w4791), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4983), .A1(w4790), .A2(w4984) );
	vdp_lfsr_bit g4812 (.Q(w4795), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4982), .A1(w4791), .A2(w4981) );
	vdp_lfsr_bit g4813 (.Q(w4797), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4979), .A1(w4795), .A2(w4980) );
	vdp_bufif0 g4814 (.A(w4772), .Z(VRAMA[2]), .nE(w6313) );
	vdp_bufif0 g4815 (.A(1'b1), .Z(VRAMA[2]), .nE(w5002) );
	vdp_notif0 g4816 (.A(w4797), .nZ(DB[5]), .nE(w5111) );
	vdp_aon22 g4817 (.Z(w4796), .B2(w4788), .B1(w4976), .A1(w4975), .A2(w4749) );
	vdp_dlatch_inv g4818 (.nQ(w4808), .D(w4801), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g4819 (.nQ(w4803), .D(w4755), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g4820 (.Z(w4802), .B(w4803), .A(DCLK2) );
	vdp_nand g4821 (.Z(w4801), .B(HCLK1), .A(w4434) );
	vdp_nand g4822 (.Z(w4755), .B(HCLK1), .A(w26) );
	vdp_sr_bit g4823 (.Q(w4800), .D(w6300), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4824 (.Q(w6300), .D(w6299), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4825 (.Q(w6299), .D(w4805), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4826 (.Z(w4816), .B2(w4800), .B1(w5105), .A1(DB[6]), .A2(w5106) );
	vdp_notif0 g4827 (.A(w4814), .nZ(VRAMA[3]), .nE(w4968) );
	vdp_lfsr_bit g4828 (.Q(w4818), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6562), .A1(w4816), .A2(w6563) );
	vdp_lfsr_bit g4829 (.Q(w4819), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6560), .A1(w4818), .A2(w6561) );
	vdp_lfsr_bit g4830 (.Q(w4822), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6558), .A1(w4819), .A2(w6559) );
	vdp_lfsr_bit g4831 (.Q(w4823), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6556), .A1(w4822), .A2(w6557) );
	vdp_lfsr_bit g4832 (.Q(w4828), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6554), .A1(w4823), .A2(w6555) );
	vdp_lfsr_bit g4833 (.Q(w4827), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6552), .A1(w4828), .A2(w6553) );
	vdp_lfsr_bit g4834 (.Q(w4830), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6550), .A1(w4827), .A2(w6551) );
	vdp_lfsr_bit g4835 (.Q(w4832), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6549), .A1(w4830), .A2(w6548) );
	vdp_lfsr_bit g4836 (.Q(w4834), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4948), .A1(w4832), .A2(w6547) );
	vdp_lfsr_bit g4837 (.Q(w4836), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5109), .A1(w4834), .A2(w5110) );
	vdp_lfsr_bit g4838 (.Q(w4838), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4994), .A1(w4836), .A2(w4995) );
	vdp_lfsr_bit g4839 (.Q(w4840), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4991), .A1(w4838), .A2(w4992) );
	vdp_lfsr_bit g4840 (.Q(w4842), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4989), .A1(w4840), .A2(w4990) );
	vdp_lfsr_bit g4841 (.Q(w4845), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6545), .A1(w4842), .A2(w6544) );
	vdp_lfsr_bit g4842 (.Q(w4846), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4986), .A1(w4845), .A2(w4987) );
	vdp_lfsr_bit g4843 (.Q(w4847), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6542), .A1(w4846), .A2(w6543) );
	vdp_lfsr_bit g4844 (.Q(w4852), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6546), .A1(w4847), .A2(w6616) );
	vdp_lfsr_bit g4845 (.Q(w4851), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4983), .A1(w4852), .A2(w4984) );
	vdp_lfsr_bit g4846 (.Q(w4854), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4982), .A1(w4851), .A2(w4981) );
	vdp_lfsr_bit g4847 (.Q(w4798), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4979), .A1(w4854), .A2(w4980) );
	vdp_bufif0 g4848 (.A(w4832), .Z(VRAMA[3]), .nE(w6313) );
	vdp_bufif0 g4849 (.A(w4796), .Z(VRAMA[3]), .nE(w5002) );
	vdp_notif0 g4850 (.A(w4798), .nZ(DB[6]), .nE(w5111) );
	vdp_aon22 g4851 (.Z(w4855), .B2(w4789), .B1(w4976), .A1(w4975), .A2(w4797) );
	vdp_sr_bit g4852 (.Q(w4810), .D(w4808), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g4853 (.Q(w4804), .D(w4803), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_and g4854 (.Z(w4806), .B(w4808), .A(DCLK2) );
	vdp_and g4855 (.Z(w4812), .B(DCLK2), .A(w4810) );
	vdp_and g4856 (.Z(w4809), .B(w4804), .A(DCLK2) );
	vdp_sr_bit g4857 (.Q(w4867), .D(w6301), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4858 (.Q(w6301), .D(w6302), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4859 (.Q(w6302), .D(w4811), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4860 (.Z(w4815), .B2(w4867), .B1(w5105), .A1(DB[7]), .A2(w5106) );
	vdp_notif0 g4861 (.A(w4865), .nZ(VRAMA[4]), .nE(w4968) );
	vdp_lfsr_bit g4862 (.Q(w4817), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6562), .A1(w4815), .A2(w6563) );
	vdp_lfsr_bit g4863 (.Q(w4820), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6560), .A1(w4817), .A2(w6561) );
	vdp_lfsr_bit g4864 (.Q(w4821), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6558), .A1(w4820), .A2(w6559) );
	vdp_lfsr_bit g4865 (.Q(w4824), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6556), .A1(w4821), .A2(w6557) );
	vdp_lfsr_bit g4866 (.Q(w4825), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6554), .A1(w4824), .A2(w6555) );
	vdp_lfsr_bit g4867 (.Q(w4826), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6552), .A1(w4825), .A2(w6553) );
	vdp_lfsr_bit g4868 (.Q(w4829), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6550), .A1(w4826), .A2(w6551) );
	vdp_lfsr_bit g4869 (.Q(w4831), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6549), .A1(w4829), .A2(w6548) );
	vdp_lfsr_bit g4870 (.Q(w4833), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4948), .A1(w4831), .A2(w6547) );
	vdp_lfsr_bit g4871 (.Q(w4835), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5109), .A1(w4833), .A2(w5110) );
	vdp_lfsr_bit g4872 (.Q(w4837), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4994), .A1(w4835), .A2(w4995) );
	vdp_lfsr_bit g4873 (.Q(w4839), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4991), .A1(w4837), .A2(w4992) );
	vdp_lfsr_bit g4874 (.Q(w4841), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4989), .A1(w4839), .A2(w4990) );
	vdp_lfsr_bit g4875 (.Q(w4844), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6545), .A1(w4841), .A2(w6544) );
	vdp_lfsr_bit g4876 (.Q(w4843), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4986), .A1(w4844), .A2(w4987) );
	vdp_lfsr_bit g4877 (.Q(w4848), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6542), .A1(w4843), .A2(w6543) );
	vdp_lfsr_bit g4878 (.Q(w4849), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6546), .A1(w4848), .A2(w6616) );
	vdp_lfsr_bit g4879 (.Q(w4850), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4983), .A1(w4849), .A2(w4984) );
	vdp_lfsr_bit g4880 (.Q(w4853), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4982), .A1(w4850), .A2(w4981) );
	vdp_lfsr_bit g4881 (.Q(w4869), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4979), .A1(w4853), .A2(w4980) );
	vdp_bufif0 g4882 (.A(w4831), .Z(VRAMA[4]), .nE(w6313) );
	vdp_bufif0 g4883 (.A(w4855), .Z(VRAMA[4]), .nE(w5002) );
	vdp_notif0 g4884 (.A(w4869), .nZ(DB[7]), .nE(w5111) );
	vdp_aon22 g4885 (.Z(w4870), .B2(w4847), .B1(w4976), .A1(w4975), .A2(w4798) );
	vdp_aon22 g4886 (.Z(w4864), .B2(w4857), .B1(w117), .A1(w4813), .A2(w4863) );
	vdp_not g4887 (.nZ(w4813), .A(w117) );
	vdp_comp_str g4888 (.nZ(w4858), .A(w4809), .Z(w4859) );
	vdp_comp_str g4889 (.nZ(w4862), .A(w4812), .Z(w4861) );
	vdp_sr_bit g4890 (.Q(w4866), .D(w6304), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4891 (.Q(w6304), .D(w6303), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4892 (.Q(w6303), .D(w4860), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4893 (.Z(w4910), .B2(w4866), .B1(w5105), .A1(DB[8]), .A2(w5106) );
	vdp_notif0 g4894 (.A(w4864), .nZ(VRAMA[5]), .nE(w4968) );
	vdp_lfsr_bit g4895 (.Q(w4908), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6562), .A1(w4910), .A2(w6563) );
	vdp_lfsr_bit g4896 (.Q(w4905), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6560), .A1(w4908), .A2(w6561) );
	vdp_lfsr_bit g4897 (.Q(w4904), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6558), .A1(w4905), .A2(w6559) );
	vdp_lfsr_bit g4898 (.Q(w4901), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6556), .A1(w4904), .A2(w6557) );
	vdp_lfsr_bit g4899 (.Q(w4900), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6554), .A1(w4901), .A2(w6555) );
	vdp_lfsr_bit g4900 (.Q(w4897), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6552), .A1(w4900), .A2(w6553) );
	vdp_lfsr_bit g4901 (.Q(w4896), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6550), .A1(w4897), .A2(w6551) );
	vdp_lfsr_bit g4902 (.Q(w4874), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6549), .A1(w4896), .A2(w6548) );
	vdp_lfsr_bit g4903 (.Q(w4893), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4948), .A1(w4874), .A2(w6547) );
	vdp_lfsr_bit g4904 (.Q(w4868), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5109), .A1(w4893), .A2(w5110) );
	vdp_lfsr_bit g4905 (.Q(w4890), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4994), .A1(w4868), .A2(w4995) );
	vdp_lfsr_bit g4906 (.Q(w4889), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4991), .A1(w4890), .A2(w4992) );
	vdp_lfsr_bit g4907 (.Q(w4886), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4989), .A1(w4889), .A2(w4990) );
	vdp_lfsr_bit g4908 (.Q(w4884), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6545), .A1(w4886), .A2(w6544) );
	vdp_lfsr_bit g4909 (.Q(w4883), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4986), .A1(w4884), .A2(w4987) );
	vdp_lfsr_bit g4910 (.Q(w4872), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6542), .A1(w4883), .A2(w6543) );
	vdp_lfsr_bit g4911 (.Q(w4879), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6546), .A1(w4872), .A2(w6616) );
	vdp_lfsr_bit g4912 (.Q(w4877), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4983), .A1(w4879), .A2(w4984) );
	vdp_lfsr_bit g4913 (.Q(w4875), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4982), .A1(w4877), .A2(w4981) );
	vdp_lfsr_bit g4914 (.Q(w4892), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4979), .A1(w4875), .A2(w4980) );
	vdp_bufif0 g4915 (.A(w4874), .Z(VRAMA[5]), .nE(w6313) );
	vdp_bufif0 g4916 (.A(w4870), .Z(VRAMA[5]), .nE(w5002) );
	vdp_notif0 g4917 (.A(w4892), .nZ(DB[8]), .nE(w5111) );
	vdp_aon22 g4918 (.Z(w4871), .B2(w4848), .B1(w4976), .A1(w4975), .A2(w4869) );
	vdp_slatch g4919 (.D(S[0]), .nC(w4862), .C(w4861), .Q(w4915) );
	vdp_slatch g4920 (.D(S[0]), .nC(w4858), .C(w4859), .Q(w4856) );
	vdp_aoi22 g4921 (.Z(w4863), .B2(w4914), .B1(w4915), .A1(w4913), .A2(w4856) );
	vdp_sr_bit g4922 (.Q(w4922), .D(w6306), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4923 (.Q(w6306), .D(w6305), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4924 (.Q(w6305), .D(w4911), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4925 (.Z(w4909), .B2(w4922), .B1(w5105), .A1(DB[9]), .A2(w5106) );
	vdp_notif0 g4926 (.A(w4912), .nZ(VRAMA[6]), .nE(w4968) );
	vdp_lfsr_bit g4927 (.Q(w4907), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6562), .A1(w4909), .A2(w6563) );
	vdp_lfsr_bit g4928 (.Q(w4906), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6560), .A1(w4907), .A2(w6561) );
	vdp_lfsr_bit g4929 (.Q(w4903), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6558), .A1(w4906), .A2(w6559) );
	vdp_lfsr_bit g4930 (.Q(w4902), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6556), .A1(w4903), .A2(w6557) );
	vdp_lfsr_bit g4931 (.Q(w4899), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6554), .A1(w4902), .A2(w6555) );
	vdp_lfsr_bit g4932 (.Q(w4898), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6552), .A1(w4899), .A2(w6553) );
	vdp_lfsr_bit g4933 (.Q(w4895), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6550), .A1(w4898), .A2(w6551) );
	vdp_lfsr_bit g4934 (.Q(w4873), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6549), .A1(w4895), .A2(w6548) );
	vdp_lfsr_bit g4935 (.Q(w4894), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4948), .A1(w4873), .A2(w6547) );
	vdp_lfsr_bit g4936 (.Q(w4920), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5109), .A1(w4894), .A2(w5110) );
	vdp_lfsr_bit g4937 (.Q(w4891), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4994), .A1(w4920), .A2(w4995) );
	vdp_lfsr_bit g4938 (.Q(w4888), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4991), .A1(w4891), .A2(w4992) );
	vdp_lfsr_bit g4939 (.Q(w4887), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4989), .A1(w4888), .A2(w4990) );
	vdp_lfsr_bit g4940 (.Q(w4885), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6545), .A1(w4887), .A2(w6544) );
	vdp_lfsr_bit g4941 (.Q(w4882), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4986), .A1(w4885), .A2(w4987) );
	vdp_lfsr_bit g4942 (.Q(w4881), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6542), .A1(w4882), .A2(w6543) );
	vdp_lfsr_bit g4943 (.Q(w4880), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6546), .A1(w4881), .A2(w6616) );
	vdp_lfsr_bit g4944 (.Q(w4878), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4983), .A1(w4880), .A2(w4984) );
	vdp_lfsr_bit g4945 (.Q(w4876), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4982), .A1(w4878), .A2(w4981) );
	vdp_lfsr_bit g4946 (.Q(w4917), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4979), .A1(w4876), .A2(w4980) );
	vdp_bufif0 g4947 (.A(w4873), .Z(VRAMA[6]), .nE(w6313) );
	vdp_bufif0 g4948 (.A(w4871), .Z(VRAMA[6]), .nE(w5002) );
	vdp_notif0 g4949 (.A(w4917), .nZ(DB[9]), .nE(w5111) );
	vdp_aon22 g4950 (.Z(w4919), .B2(w4872), .B1(w4976), .A1(w4975), .A2(w4892) );
	vdp_aoi22 g4951 (.Z(w4912), .B2(w4914), .B1(w4924), .A1(w4913), .A2(w4916) );
	vdp_slatch g4952 (.D(S[1]), .nC(w4862), .C(w4861), .Q(w4924) );
	vdp_slatch g4953 (.D(S[1]), .nC(w4858), .C(w4859), .Q(w4916) );
	vdp_sr_bit g4954 (.Q(w4921), .D(w6308), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4955 (.Q(w6308), .D(w6307), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4956 (.Q(w6307), .D(w4925), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4957 (.Z(w4967), .B2(w4921), .B1(w5105), .A1(DB[10]), .A2(w5106) );
	vdp_notif0 g4958 (.A(w4970), .nZ(VRAMA[7]), .nE(w4971) );
	vdp_lfsr_bit g4959 (.Q(w4966), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6562), .A1(w4967), .A2(w6563) );
	vdp_lfsr_bit g4960 (.Q(w4961), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6560), .A1(w4966), .A2(w6561) );
	vdp_lfsr_bit g4961 (.Q(w4962), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6558), .A1(w4961), .A2(w6559) );
	vdp_lfsr_bit g4962 (.Q(w4956), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6556), .A1(w4962), .A2(w6557) );
	vdp_lfsr_bit g4963 (.Q(w4957), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6554), .A1(w4956), .A2(w6555) );
	vdp_lfsr_bit g4964 (.Q(w4954), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6552), .A1(w4957), .A2(w6553) );
	vdp_lfsr_bit g4965 (.Q(w4952), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6550), .A1(w4954), .A2(w6551) );
	vdp_lfsr_bit g4966 (.Q(w4918), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6549), .A1(w4952), .A2(w6548) );
	vdp_lfsr_bit g4967 (.Q(w4949), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4948), .A1(w4918), .A2(w6547) );
	vdp_lfsr_bit g4968 (.Q(w4944), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5109), .A1(w4949), .A2(w5110) );
	vdp_lfsr_bit g4969 (.Q(w4946), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4994), .A1(w4944), .A2(w4995) );
	vdp_lfsr_bit g4970 (.Q(w4943), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4991), .A1(w4946), .A2(w4992) );
	vdp_lfsr_bit g4971 (.Q(w4942), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4989), .A1(w4943), .A2(w4990) );
	vdp_lfsr_bit g4972 (.Q(w4939), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6545), .A1(w4942), .A2(w6544) );
	vdp_lfsr_bit g4973 (.Q(w4937), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4986), .A1(w4939), .A2(w4987) );
	vdp_lfsr_bit g4974 (.Q(w4935), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6542), .A1(w4937), .A2(w6543) );
	vdp_lfsr_bit g4975 (.Q(w4933), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6546), .A1(w4935), .A2(w6616) );
	vdp_lfsr_bit g4976 (.Q(w4931), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4983), .A1(w4933), .A2(w4984) );
	vdp_lfsr_bit g4977 (.Q(w4929), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4982), .A1(w4931), .A2(w4981) );
	vdp_lfsr_bit g4978 (.Q(w4927), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4979), .A1(w4929), .A2(w4980) );
	vdp_bufif0 g4979 (.A(w4918), .Z(VRAMA[7]), .nE(w6313) );
	vdp_bufif0 g4980 (.A(w4919), .Z(VRAMA[7]), .nE(w5002) );
	vdp_notif0 g4981 (.A(w4927), .nZ(DB[10]), .nE(w5111) );
	vdp_aon22 g4982 (.Z(w4926), .B2(w4881), .B1(w4976), .A1(w4975), .A2(w4917) );
	vdp_aoi22 g4983 (.Z(w4970), .B2(w4914), .B1(w4972), .A1(w4913), .A2(w4923) );
	vdp_slatch g4984 (.D(S[2]), .nC(w4862), .C(w4861), .Q(w4972) );
	vdp_slatch g4985 (.D(S[2]), .nC(w4858), .C(w4859), .Q(w4923) );
	vdp_sr_bit g4986 (.Q(w4997), .D(w27), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4987 (.Q(w4996), .D(w21), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4988 (.Z(w4964), .B2(w4411), .B1(w5105), .A1(DB[11]), .A2(w5106) );
	vdp_notif0 g4989 (.A(w4969), .nZ(VRAMA[8]), .nE(w4971) );
	vdp_lfsr_bit g4990 (.Q(w4965), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6562), .A1(w4964), .A2(w6563) );
	vdp_lfsr_bit g4991 (.Q(w4960), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6560), .A1(w4965), .A2(w6561) );
	vdp_lfsr_bit g4992 (.Q(w4963), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6558), .A1(w4960), .A2(w6559) );
	vdp_lfsr_bit g4993 (.Q(w4959), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6556), .A1(w4963), .A2(w6557) );
	vdp_lfsr_bit g4994 (.Q(w4958), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6554), .A1(w4959), .A2(w6555) );
	vdp_lfsr_bit g4995 (.Q(w4955), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6552), .A1(w4958), .A2(w6553) );
	vdp_lfsr_bit g4996 (.Q(w4953), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6550), .A1(w4955), .A2(w6551) );
	vdp_lfsr_bit g4997 (.Q(w4951), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6549), .A1(w4953), .A2(w6548) );
	vdp_lfsr_bit g4998 (.Q(w4950), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4948), .A1(w4951), .A2(w6547) );
	vdp_lfsr_bit g4999 (.Q(w4947), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5109), .A1(w4950), .A2(w5110) );
	vdp_lfsr_bit g5000 (.Q(w4945), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4994), .A1(w4947), .A2(w4995) );
	vdp_lfsr_bit g5001 (.Q(w4941), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4991), .A1(w4945), .A2(w4992) );
	vdp_lfsr_bit g5002 (.Q(w4940), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4989), .A1(w4941), .A2(w4990) );
	vdp_lfsr_bit g5003 (.Q(w4938), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6545), .A1(w4940), .A2(w6544) );
	vdp_lfsr_bit g5004 (.Q(w4936), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4986), .A1(w4938), .A2(w4987) );
	vdp_lfsr_bit g5005 (.Q(w4934), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6542), .A1(w4936), .A2(w6543) );
	vdp_lfsr_bit g5006 (.Q(w4932), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6546), .A1(w4934), .A2(w6616) );
	vdp_lfsr_bit g5007 (.Q(w4930), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4983), .A1(w4932), .A2(w4984) );
	vdp_lfsr_bit g5008 (.Q(w4928), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4982), .A1(w4930), .A2(w4981) );
	vdp_lfsr_bit g5009 (.Q(w4993), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4979), .A1(w4928), .A2(w4980) );
	vdp_bufif0 g5010 (.A(1'b0), .Z(VRAMA[0]), .nE(w6313) );
	vdp_bufif0 g5011 (.A(w4926), .Z(VRAMA[8]), .nE(w5002) );
	vdp_notif0 g5012 (.A(w4993), .nZ(DB[11]), .nE(w5111) );
	vdp_aon22 g5013 (.Z(w5003), .B2(w4977), .B1(w4976), .A1(w4975), .A2(w4927) );
	vdp_aoi22 g5014 (.Z(w4969), .B2(w4914), .B1(w4973), .A1(w4913), .A2(w4974) );
	vdp_slatch g5015 (.D(S[3]), .nC(w4862), .C(w4861), .Q(w4973) );
	vdp_slatch g5016 (.D(S[3]), .nC(w4858), .C(w4859), .Q(w4974) );
	vdp_bufif0 g5017 (.A(1'b0), .Z(VRAMA[0]), .nE(w5002) );
	vdp_bufif0 g5018 (.A(w5005), .Z(VRAMA[8]), .nE(w5009) );
	vdp_aon22 g5019 (.Z(w5032), .B2(w4420), .B1(w5105), .A1(DB[3]), .A2(w5106) );
	vdp_lfsr_bit g5020 (.Q(w5030), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6562), .A1(w5032), .A2(w6563) );
	vdp_lfsr_bit g5021 (.Q(w5028), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6560), .A1(w5030), .A2(w6561) );
	vdp_lfsr_bit g5022 (.Q(w5026), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6558), .A1(w5028), .A2(w6559) );
	vdp_lfsr_bit g5023 (.Q(w5024), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6556), .A1(w5026), .A2(w6557) );
	vdp_lfsr_bit g5024 (.Q(w5021), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6554), .A1(w5024), .A2(w6555) );
	vdp_lfsr_bit g5025 (.Q(w5020), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6552), .A1(w5021), .A2(w6553) );
	vdp_lfsr_bit g5026 (.Q(w5018), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6550), .A1(w5020), .A2(w6551) );
	vdp_lfsr_bit g5027 (.Q(w5016), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6549), .A1(w5018), .A2(w6548) );
	vdp_lfsr_bit g5028 (.Q(w5001), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4948), .A1(w5016), .A2(w6547) );
	vdp_lfsr_bit g5029 (.Q(w4999), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5109), .A1(w5001), .A2(w5110) );
	vdp_notif0 g5030 (.A(w4999), .nZ(DB[3]), .nE(w5111) );
	vdp_not g5031 (.nZ(w4988), .A(M5) );
	vdp_not g5032 (.nZ(w4998), .A(H40) );
	vdp_notif0 g5033 (.A(1'b1), .nZ(VRAMA[0]), .nE(w4968) );
	vdp_aoi22 g5034 (.Z(w4857), .B2(w5036), .B1(w5001), .A1(w4913), .A2(w4999) );
	vdp_not g5035 (.nZ(w5034), .A(M5) );
	vdp_or g5036 (.Z(w5035), .B(w4997), .A(w4996) );
	vdp_sr_bit g5037 (.Q(w5006), .D(w8), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5038 (.Q(w5012), .D(w28), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_comp_we g5039 (.nZ(w4979), .A(w5004), .Z(w4980) );
	vdp_comp_we g5040 (.nZ(w4982), .A(w5004), .Z(w4981) );
	vdp_comp_we g5041 (.nZ(w4983), .A(w5004), .Z(w4984) );
	vdp_comp_we g5042 (.nZ(w6546), .A(w5004), .Z(w6616) );
	vdp_comp_we g5043 (.nZ(w6542), .A(w5004), .Z(w6543) );
	vdp_comp_we g5044 (.nZ(w4976), .A(H40), .Z(w4975) );
	vdp_comp_we g5045 (.nZ(w4986), .A(w5004), .Z(w4987) );
	vdp_comp_we g5046 (.nZ(w6545), .A(w5004), .Z(w6544) );
	vdp_comp_we g5047 (.nZ(w4989), .A(w5004), .Z(w4990) );
	vdp_comp_we g5048 (.nZ(w4991), .A(w5004), .Z(w4992) );
	vdp_comp_we g5049 (.nZ(w4994), .A(w5004), .Z(w4995) );
	vdp_comp_we g5050 (.nZ(w4914), .A(w4996), .Z(w4913) );
	vdp_not g5051 (.nZ(w4971), .A(w5000) );
	vdp_not g5052 (.nZ(w4968), .A(w5000) );
	vdp_not g5053 (.nZ(w5002), .A(w5008) );
	vdp_not g5054 (.nZ(w6313), .A(w4985) );
	vdp_and g5055 (.Z(w4985), .B(w5006), .A(w4988) );
	vdp_oai21 g5056 (.Z(w5011), .B(w4988), .A1(w5012), .A2(w5006) );
	vdp_aon333 g5057 (.Z(w4374), .B1(M5), .A1(1'b1), .C1(M5), .A2(w4988), .A3(w4951), .B2(w4934), .B3(w4998), .C2(H40), .C3(w4993) );
	vdp_aon22 g5058 (.Z(w5031), .B2(w4426), .B1(w5105), .A1(DB[2]), .A2(w5106) );
	vdp_lfsr_bit g5059 (.Q(w5029), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6562), .A1(w5031), .A2(w6563) );
	vdp_lfsr_bit g5060 (.Q(w5027), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6560), .A1(w5029), .A2(w6561) );
	vdp_lfsr_bit g5061 (.Q(w5025), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6558), .A1(w5027), .A2(w6559) );
	vdp_lfsr_bit g5062 (.Q(w5023), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6556), .A1(w5025), .A2(w6557) );
	vdp_lfsr_bit g5063 (.Q(w5022), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6554), .A1(w5023), .A2(w6555) );
	vdp_lfsr_bit g5064 (.Q(w5019), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6552), .A1(w5022), .A2(w6553) );
	vdp_lfsr_bit g5065 (.Q(w5017), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6550), .A1(w5019), .A2(w6551) );
	vdp_lfsr_bit g5066 (.Q(w5015), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6549), .A1(w5017), .A2(w6548) );
	vdp_lfsr_bit g5067 (.Q(w5014), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4948), .A1(w5015), .A2(w6547) );
	vdp_lfsr_bit g5068 (.Q(w5013), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5109), .A1(w5014), .A2(w5110) );
	vdp_notif0 g5069 (.A(w5013), .nZ(DB[2]), .nE(w5111) );
	vdp_aoi22 g5070 (.Z(w4865), .B2(w5036), .B1(w5014), .A1(w4913), .A2(w5013) );
	vdp_aoi22 g5071 (.Z(w5048), .B2(w5036), .B1(w5049), .A1(w4913), .A2(w4376) );
	vdp_notif0 g5072 (.A(w5048), .nZ(VRAMA[9]), .nE(w4971) );
	vdp_slatch g5074 (.D(S[4]), .nC(w4859), .C(w4858), .Q(w4376) );
	vdp_and g5075 (.Z(w5000), .B(w5034), .A(w5035) );
	vdp_slatch g5076 (.D(REG_BUS[0]), .nC(w5108), .C(w5107), .Q(w4977) );
	vdp_slatch g5077 (.D(REG_BUS[7]), .nC(w5108), .C(w5107), .Q(w5007) );
	vdp_bufif0 g5078 (.A(w5003), .Z(VRAMA[9]), .nE(w5038) );
	vdp_bufif0 g5079 (.A(w5007), .Z(VRAMA[16]), .nE(w5038) );
	vdp_and g5080 (.Z(w5008), .B(w5006), .A(M5) );
	vdp_not g5081 (.nZ(w5038), .A(w5008) );
	vdp_not g5082 (.nZ(w5009), .A(w5010) );
	vdp_not g5083 (.nZ(w5010), .A(w5011) );
	vdp_xor g5084 (.Z(w5037), .B(w5007), .A(VRAMA[16]) );
	vdp_xor g5085 (.Z(w5041), .B(w5043), .A(w5042) );
	vdp_and3 g5086 (.Z(w6160), .B(w5047), .A(w5044), .C(M5) );
	vdp_nor g5087 (.Z(w5043), .B(H40), .A(w4977) );
	vdp_nor g5088 (.Z(w5042), .B(H40), .A(VRAMA[9]) );
	vdp_aon22 g5089 (.Z(w5067), .B2(w4417), .B1(w5105), .A1(DB[1]), .A2(w5106) );
	vdp_lfsr_bit g5090 (.Q(w5066), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6562), .A1(w5067), .A2(w6563) );
	vdp_lfsr_bit g5091 (.Q(w5065), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6560), .A1(w5066), .A2(w6561) );
	vdp_lfsr_bit g5092 (.Q(w5064), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6558), .A1(w5065), .A2(w6559) );
	vdp_lfsr_bit g5093 (.Q(w5063), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6556), .A1(w5064), .A2(w6557) );
	vdp_lfsr_bit g5094 (.Q(w5062), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6554), .A1(w5063), .A2(w6555) );
	vdp_lfsr_bit g5095 (.Q(w5061), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6552), .A1(w5062), .A2(w6553) );
	vdp_lfsr_bit g5096 (.Q(w5060), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6550), .A1(w5061), .A2(w6551) );
	vdp_lfsr_bit g5097 (.Q(w5059), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6549), .A1(w5060), .A2(w6548) );
	vdp_lfsr_bit g5098 (.Q(w5046), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w4948), .A1(w5059), .A2(w6547) );
	vdp_lfsr_bit g5099 (.Q(w5057), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5109), .A1(w5046), .A2(w5110) );
	vdp_notif0 g5100 (.A(w5057), .nZ(DB[1]), .nE(w5111) );
	vdp_slatch g5101 (.D(REG_BUS[1]), .nC(w5108), .C(w5107), .Q(w5005) );
	vdp_slatch g5102 (.D(REG_BUS[6]), .nC(w5108), .C(w5107), .Q(w5056) );
	vdp_xor g5103 (.Z(w5040), .B(w5056), .A(VRAMA[15]) );
	vdp_xor g5104 (.Z(w5039), .B(w5005), .A(VRAMA[10]) );
	vdp_aon22 g5105 (.Z(w5076), .B2(w4416), .B1(w5105), .A1(DB[0]), .A2(w5106) );
	vdp_lfsr_bit g5106 (.Q(w5077), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6562), .A1(w5076), .A2(w6563) );
	vdp_lfsr_bit g5107 (.Q(w5078), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6560), .A1(w5077), .A2(w6561) );
	vdp_lfsr_bit g5108 (.Q(w5079), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6558), .A1(w5078), .A2(w6559) );
	vdp_lfsr_bit g5109 (.Q(w5081), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6556), .A1(w5079), .A2(w6557) );
	vdp_lfsr_bit g5110 (.Q(w5080), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6554), .A1(w5081), .A2(w6555) );
	vdp_lfsr_bit g5111 (.Q(w5083), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6552), .A1(w5080), .A2(w6553) );
	vdp_lfsr_bit g5112 (.Q(w5082), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6550), .A1(w5083), .A2(w6551) );
	vdp_lfsr_bit g5113 (.Q(w5084), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6549), .A1(w5082), .A2(w6548) );
	vdp_lfsr_bit g5114 (.Q(w5058), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w4948), .A1(w5084), .A2(w6547) );
	vdp_lfsr_bit g5115 (.Q(w6312), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5109), .A1(w5058), .A2(w5110) );
	vdp_notif0 g5116 (.A(w6312), .nZ(DB[0]), .nE(w5111) );
	vdp_slatch g5117 (.D(REG_BUS[2]), .nC(w5108), .C(w5107), .Q(w5055) );
	vdp_slatch g5118 (.D(REG_BUS[5]), .nC(w5108), .C(w5107), .Q(w5099) );
	vdp_xor g5119 (.Z(w5052), .B(w5099), .A(VRAMA[14]) );
	vdp_xor g5120 (.Z(w5051), .B(w5055), .A(VRAMA[11]) );
	vdp_slatch g5121 (.D(S[5]), .nC(w4861), .C(w4862), .Q(w5070) );
	vdp_slatch g5122 (.D(S[5]), .nC(w4859), .C(w4858), .Q(w5050) );
	vdp_slatch g5123 (.D(S[6]), .nC(w4861), .C(w4862), .Q(w5071) );
	vdp_slatch g5124 (.D(S[6]), .nC(w4859), .C(w4858), .Q(w5069) );
	vdp_slatch g5125 (.D(S[7]), .nC(w4861), .C(w4862), .Q(w5104) );
	vdp_slatch g5126 (.D(S[7]), .nC(w4859), .C(w4858), .Q(w5036) );
	vdp_slatch g5127 (.D(REG_BUS[2]), .nC(w5074), .C(w5075), .Q(w5072) );
	vdp_slatch g5128 (.D(REG_BUS[5]), .nC(w5074), .C(w5075), .Q(w5068) );
	vdp_bufif0 g5129 (.A(w5055), .Z(VRAMA[9]), .nE(w5009) );
	vdp_bufif0 g5130 (.A(w5005), .Z(VRAMA[10]), .nE(w5038) );
	vdp_bufif0 g5131 (.A(w5093), .Z(VRAMA[10]), .nE(w5009) );
	vdp_bufif0 g5132 (.A(w5056), .Z(VRAMA[13]), .nE(w5009) );
	vdp_bufif0 g5133 (.A(w5099), .Z(VRAMA[14]), .nE(w5038) );
	vdp_bufif0 g5134 (.A(w5055), .Z(VRAMA[11]), .nE(w5038) );
	vdp_bufif0 g5135 (.A(w5092), .Z(VRAMA[13]), .nE(w5038) );
	vdp_bufif0 g5136 (.A(w5093), .Z(VRAMA[12]), .nE(w5038) );
	vdp_bufif0 g5137 (.A(w5092), .Z(VRAMA[11]), .nE(w5009) );
	vdp_bufif0 g5138 (.A(w5099), .Z(VRAMA[12]), .nE(w5009) );
	vdp_bufif0 g5139 (.A(w5056), .Z(VRAMA[15]), .nE(w5038) );
	vdp_slatch g5140 (.D(REG_BUS[3]), .nC(w5108), .C(w5107), .Q(w5093) );
	vdp_slatch g5141 (.D(REG_BUS[4]), .nC(w5108), .C(w5107), .Q(w5092) );
	vdp_xor g5142 (.Z(w5054), .B(w5092), .A(VRAMA[13]) );
	vdp_xor g5143 (.Z(w5053), .B(w5093), .A(VRAMA[12]) );
	vdp_dlatch_inv g5144 (.nQ(w5091), .D(w5096), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5145 (.nQ(w5090), .D(w5097), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5146 (.nQ(w5089), .D(w6418), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5147 (.nQ(w5088), .D(w6420), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5148 (.nQ(w5087), .D(w5098), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5149 (.nQ(w5086), .D(w5095), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5150 (.nQ(w5085), .D(w6419), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5151 (.nQ(w6155), .D(w5094), .nC(nDCLK1), .C(DCLK1) );
	vdp_comp_we g5152 (.nZ(w5109), .A(w5004), .Z(w5110) );
	vdp_comp_we g5153 (.nZ(w4948), .A(w5004), .Z(w6547) );
	vdp_comp_we g5154 (.nZ(w6549), .A(w5004), .Z(w6548) );
	vdp_comp_we g5155 (.nZ(w6550), .A(w5004), .Z(w6551) );
	vdp_comp_we g5156 (.nZ(w6552), .A(w5004), .Z(w6553) );
	vdp_comp_we g5157 (.nZ(w6554), .A(w5004), .Z(w6555) );
	vdp_comp_we g5158 (.nZ(w6556), .A(w5004), .Z(w6557) );
	vdp_comp_we g5159 (.nZ(w6558), .A(w5004), .Z(w6559) );
	vdp_comp_we g5160 (.nZ(w6560), .A(w5004), .Z(w6561) );
	vdp_comp_we g5161 (.nZ(w6562), .A(w5004), .Z(w6563) );
	vdp_comp_we g5162 (.nZ(w5105), .A(w106), .Z(w5106) );
	vdp_notif0 g5163 (.A(w5045), .nZ(VRAMA[10]), .nE(w4971) );
	vdp_notif0 g5164 (.A(w5073), .nZ(VRAMA[13]), .nE(w4971) );
	vdp_notif0 g5165 (.A(w5103), .nZ(VRAMA[11]), .nE(w4971) );
	vdp_notif0 g5166 (.A(w5102), .nZ(VRAMA[12]), .nE(w4971) );
	vdp_not g5167 (.nZ(w5047), .A(VRAMA[2]) );
	vdp_not g5168 (.nZ(w5073), .A(w5072) );
	vdp_not g5169 (.nZ(w5101), .A(w104) );
	vdp_aoi22 g5170 (.Z(w4814), .B2(w5036), .B1(w5046), .A1(w4913), .A2(w5057) );
	vdp_aoi22 g5171 (.Z(w5045), .B2(w5036), .B1(w5070), .A1(w4913), .A2(w5050) );
	vdp_aoi22 g5172 (.Z(w4807), .B2(w5036), .B1(w5058), .A1(w4913), .A2(w6312) );
	vdp_aoi22 g5173 (.Z(w5103), .B2(w5036), .B1(w5071), .A1(w4913), .A2(w5069) );
	vdp_aoi22 g5174 (.Z(w5102), .B2(w5036), .B1(w5104), .A1(w4913), .A2(w5036) );
	vdp_and g5175 (.Z(w5100), .B(w5101), .A(w4409) );
	vdp_nor8 g5176 (.Z(w5044), .B(w5053), .A(w5054), .C(w5052), .D(w5051), .F(w5041), .E(w5037), .G(w5039), .H(w5040) );
	vdp_not g5177 (.nZ(w5111), .A(w105) );
	vdp_comp_str g5178 (.nZ(w5108), .A(w156), .Z(w5107) );
	vdp_comp_str g5179 (.nZ(w5075), .A(w157), .Z(w5074) );
	vdp_or3 g5180 (.Z(w5004), .B(w106), .A(w105), .C(w5100) );
	vdp_not g5181 (.nZ(S[7]), .A(w5091) );
	vdp_not g5182 (.nZ(S[6]), .A(w5090) );
	vdp_not g5183 (.nZ(S[5]), .A(w5089) );
	vdp_not g5184 (.nZ(S[4]), .A(w5088) );
	vdp_not g5185 (.nZ(S[3]), .A(w5087) );
	vdp_not g5186 (.nZ(S[2]), .A(w5086) );
	vdp_not g5187 (.nZ(S[1]), .A(w5085) );
	vdp_not g5188 (.nZ(S[0]), .A(w6155) );
	vdp_aon21_sr g5189 (.Q(w5179), .A1(w5178), .A2(w6225), .B(w6226), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5190 (.Q(w6226), .A1(w5173), .A2(w6225), .B(w6564), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5191 (.Q(w6564), .A1(w5174), .A2(w6225), .B(w6565), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5192 (.Q(w6565), .A1(w5123), .A2(w6225), .B(w6566), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5193 (.Q(w6566), .A1(w5172), .A2(w6225), .B(w6567), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5194 (.Q(w6567), .A1(w5171), .A2(w6225), .B(w6568), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5195 (.Q(w6568), .A1(w5170), .A2(w6225), .B(w6569), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5196 (.Q(w6569), .A1(w5169), .A2(w6225), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5197 (.Q(w6570), .A1(w5159), .A2(w6227), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5198 (.Q(w6571), .A1(w5153), .A2(w6227), .B(w6570), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5199 (.Q(w6572), .A1(w5155), .A2(w6227), .B(w6571), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5200 (.Q(w6573), .A1(w5152), .A2(w6227), .B(w6572), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5201 (.Q(w6574), .A1(w5122), .A2(w6227), .B(w6573), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5202 (.Q(w6575), .A1(w5150), .A2(w6227), .B(w6574), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5203 (.Q(w6576), .A1(w5151), .A2(w6227), .B(w6575), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5204 (.Q(w5143), .A1(w5149), .A2(w6227), .B(w6576), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5205 (.Q(w5285), .A1(w5140), .A2(w6224), .B(w6577), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5206 (.Q(w6577), .A1(w5138), .A2(w6224), .B(w6578), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5207 (.Q(w6578), .A1(w5141), .A2(w6224), .B(w6579), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5208 (.Q(w6579), .A1(w5136), .A2(w6224), .B(w6580), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5209 (.Q(w6580), .A1(w5114), .A2(w6224), .B(w6581), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5210 (.Q(w6581), .A1(w5135), .A2(w6224), .B(w6582), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5211 (.Q(w6582), .A1(w5137), .A2(w6224), .B(w6583), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5212 (.Q(w6583), .A1(w5132), .A2(w6224), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5213 (.Q(w6585), .A1(w5184), .A2(w6223), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5214 (.Q(w6586), .A1(w5183), .A2(w6223), .B(w6585), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5215 (.Q(w6587), .A1(w5508), .A2(w6223), .B(w6586), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5216 (.Q(w6588), .A1(w5191), .A2(w6223), .B(w6587), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5217 (.Q(w6589), .A1(w5189), .A2(w6223), .B(w6588), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5218 (.Q(w6590), .A1(w5195), .A2(w6223), .B(w6589), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5219 (.Q(w6591), .A1(w5188), .A2(w6223), .B(w6590), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5220 (.Q(w5112), .A1(w5121), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .A2(w6223), .B(w6591) );
	vdp_not g5221 (.nZ(w6224), .A(nSRLOAD) );
	vdp_not g5222 (.nZ(w6223), .A(nSRLOAD) );
	vdp_not g5223 (.nZ(w6227), .A(nSRLOAD) );
	vdp_not g5224 (.nZ(w6225), .A(nSRLOAD) );
	vdp_or4 g5225 (.Z(w5177), .B(w5166), .A(w6156), .D(w5167), .C(w5165) );
	vdp_or4 g5226 (.Z(w5147), .B(w5163), .A(w5156), .D(w5161), .C(w5162) );
	vdp_or4 g5227 (.Z(w5180), .B(w5120), .A(w5121), .D(w5504), .C(w5119) );
	vdp_or4 g5228 (.Z(w5146), .B(w5118), .A(w5501), .D(w5188), .C(w5117) );
	vdp_or4 g5229 (.Z(w5142), .B(w5116), .A(w5500), .D(w5195), .C(w5115) );
	vdp_or4 g5230 (.Z(w5185), .B(w5125), .A(w5126), .D(w6157), .C(w5124) );
	vdp_or4 g5231 (.Z(w5131), .B(w5129), .A(w5130), .D(w5113), .C(w5128) );
	vdp_slatch g5232 (.Q(w5167), .D(w5232), .nC(w5157), .C(w5158) );
	vdp_comp_str g5233 (.nZ(w5157), .A(w5204), .Z(w5158) );
	vdp_slatch g5234 (.Q(w5165), .D(w5230), .nC(w5157), .C(w5158) );
	vdp_slatch g5235 (.Q(w5166), .D(w5229), .nC(w5157), .C(w5158) );
	vdp_slatch g5236 (.Q(w6156), .D(w5228), .nC(w5157), .C(w5158) );
	vdp_slatch g5237 (.Q(w5161), .D(w5227), .nC(w5157), .C(w5158) );
	vdp_slatch g5238 (.Q(w5162), .D(w5226), .nC(w5157), .C(w5158) );
	vdp_slatch g5239 (.Q(w5163), .D(w5224), .nC(w5157), .C(w5158) );
	vdp_slatch g5240 (.Q(w5156), .D(w5220), .nC(w5157), .C(w5158) );
	vdp_slatch g5241 (.Q(w5113), .D(w6220), .nC(w5127), .C(w5187) );
	vdp_slatch g5242 (.Q(w5128), .D(w6221), .nC(w5127), .C(w5187) );
	vdp_slatch g5243 (.Q(w5129), .D(w6222), .nC(w5127), .C(w5187) );
	vdp_slatch g5244 (.Q(w5130), .D(w5210), .nC(w5127), .C(w5187) );
	vdp_slatch g5245 (.Q(w6157), .D(w5208), .nC(w5127), .C(w5187) );
	vdp_slatch g5246 (.Q(w5124), .D(w5207), .nC(w5127), .C(w5187) );
	vdp_slatch g5247 (.Q(w5125), .D(w5206), .nC(w5127), .C(w5187) );
	vdp_slatch g5248 (.Q(w5126), .D(w5203), .nC(w5127), .C(w5187) );
	vdp_aon22 g5249 (.Z(w5240), .B2(w5133), .B1(w5193), .A1(w5185), .A2(w5145) );
	vdp_comp_we g5250 (.nZ(w5133), .A(w5192), .Z(w5145) );
	vdp_notif0 g5251 (.A(w5186), .nZ(DB[11]), .nE(w5202) );
	vdp_notif0 g5252 (.A(w5190), .nZ(DB[3]), .nE(w5202) );
	vdp_notif0 g5253 (.A(w5134), .nZ(DB[10]), .nE(w5202) );
	vdp_notif0 g5254 (.A(w5139), .nZ(DB[2]), .nE(w5202) );
	vdp_notif0 g5255 (.A(w5154), .nZ(DB[1]), .nE(w5202) );
	vdp_notif0 g5256 (.A(w5196), .nZ(DB[9]), .nE(w5202) );
	vdp_notif0 g5257 (.A(w5175), .nZ(DB[8]), .nE(w5202) );
	vdp_notif0 g5258 (.A(w5176), .nZ(DB[0]), .nE(w5202) );
	vdp_not g5259 (.nZ(w5181), .A(w5180) );
	vdp_aon22 g5260 (.Z(w5213), .B2(w5133), .B1(w5144), .A1(w5131), .A2(w5145) );
	vdp_aon22 g5261 (.Z(w5218), .B2(w5133), .B1(w5148), .A1(w5147), .A2(w5145) );
	vdp_aon22 g5262 (.Z(w5235), .B2(w5133), .B1(w5181), .A1(w5177), .A2(w5145) );
	vdp_comp_str g5263 (.nZ(w5127), .A(w5204), .Z(w5187) );
	vdp_not g5264 (.nZ(w5193), .A(w5194) );
	vdp_not g5265 (.nZ(w5144), .A(w5142) );
	vdp_not g5266 (.nZ(w5148), .A(w5146) );
	vdp_and3 g5267 (.Z(w6205), .B(w5216), .A(w5147), .C(w5146) );
	vdp_and3 g5268 (.Z(w5222), .B(w5236), .A(w5177), .C(w5180) );
	vdp_and3 g5269 (.Z(w5238), .B(w5214), .A(w5131), .C(w5142) );
	vdp_and3 g5270 (.Z(w5567), .B(w5185), .A(w5197), .C(w5194) );
	vdp_aon2222 g5271 (.Z(w5190), .B2(w5191), .B1(w5200), .A1(w5201), .A2(w5183), .D2(w5121), .D1(w5198), .C1(w5199), .C2(w5195) );
	vdp_aon2222 g5272 (.Z(w5186), .B2(w5508), .B1(w5200), .A1(w5201), .A2(w5184), .D2(w5188), .D1(w5198), .C1(w5199), .C2(w5189) );
	vdp_aon2222 g5273 (.Z(w5134), .B2(w5135), .B1(w5200), .A1(w5201), .A2(w5132), .D2(w5138), .D1(w5198), .C1(w5199), .C2(w5136) );
	vdp_aon2222 g5274 (.Z(w5139), .B2(w5114), .B1(w5200), .A1(w5201), .A2(w5137), .D2(w5140), .D1(w5198), .C1(w5199), .C2(w5141) );
	vdp_aon2222 g5275 (.Z(w5154), .B2(w5152), .B1(w5200), .A1(w5201), .A2(w5153), .D2(w5149), .D1(w5198), .C1(w5199), .C2(w5150) );
	vdp_aon2222 g5276 (.Z(w5196), .B2(w5155), .B1(w5200), .A1(w5201), .A2(w5159), .D2(w5151), .D1(w5198), .C1(w5199), .C2(w5122) );
	vdp_aon2222 g5277 (.Z(w5175), .B2(w5171), .B1(w5200), .A1(w5201), .A2(w5169), .D2(w5173), .D1(w5198), .C1(w5199), .C2(w5123) );
	vdp_aon2222 g5278 (.Z(w5176), .B2(w5172), .B1(w5200), .A1(w5201), .A2(w5170), .D2(w5178), .D1(w5198), .C1(w5199), .C2(w5174) );
	vdp_slatch g5279 (.Q(w5232), .D(w5252), .nC(w5251), .C(w5231) );
	vdp_comp_str g5280 (.nZ(w5251), .A(w5250), .Z(w5231) );
	vdp_slatch g5281 (.Q(w5230), .D(w5256), .nC(w5251), .C(w5231) );
	vdp_slatch g5282 (.Q(w5229), .D(w5257), .nC(w5251), .C(w5231) );
	vdp_slatch g5283 (.Q(w5228), .D(w5260), .nC(w5251), .C(w5231) );
	vdp_slatch g5284 (.Q(w5227), .D(w5265), .nC(w5266), .C(w5225) );
	vdp_comp_str g5285 (.nZ(w5266), .A(w5261), .Z(w5225) );
	vdp_slatch g5286 (.Q(w5226), .D(w5268), .nC(w5266), .C(w5225) );
	vdp_slatch g5287 (.Q(w5224), .D(w5269), .nC(w5266), .C(w5225) );
	vdp_slatch g5288 (.Q(w5220), .D(w5271), .nC(w5266), .C(w5225) );
	vdp_sr_bit g5289 (.Q(w5273), .D(w5143), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5290 (.nQ(w5219), .D(w5275), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5291 (.nQ(w5277), .D(w5217), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5292 (.nQ(w5215), .D(w5284), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5293 (.nQ(w5290), .D(w6198), .nC(nDCLK2), .C(DCLK2) );
	vdp_slatch g5294 (.Q(w5210), .D(w5252), .nC(w5292), .C(w5212) );
	vdp_slatch g5295 (.Q(w6220), .D(w5256), .nC(w5292), .C(w5212) );
	vdp_slatch g5296 (.Q(w6221), .D(w5257), .nC(w5292), .C(w5212) );
	vdp_slatch g5297 (.Q(w6222), .D(w5260), .nC(w5292), .C(w5212) );
	vdp_comp_str g5298 (.nZ(w5292), .A(w5291), .Z(w5212) );
	vdp_slatch g5299 (.Q(w5208), .D(w5265), .nC(w5303), .C(w5205) );
	vdp_slatch g5300 (.Q(w5207), .D(w5268), .nC(w5303), .C(w5205) );
	vdp_slatch g5301 (.Q(w5206), .D(w5269), .nC(w5303), .C(w5205) );
	vdp_slatch g5302 (.Q(w5203), .D(w5271), .nC(w5303), .C(w5205) );
	vdp_comp_str g5303 (.nZ(w5303), .A(w5308), .Z(w5205) );
	vdp_dlatch_inv g5304 (.nQ(w5301), .D(w5300), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5305 (.nQ(w5304), .D(w6197), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5306 (.nQ(w5239), .D(w5307), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5307 (.Z(w5306), .B(w5239), .A(w5243) );
	vdp_xor g5308 (.Z(w6216), .B(w5215), .A(w5243) );
	vdp_xor g5309 (.Z(w5274), .B(w5219), .A(w5243) );
	vdp_xor g5310 (.Z(w6165), .B(w6164), .A(w5243) );
	vdp_sr_bit g5311 (.Q(w6219), .D(w5179), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5312 (.nQ(w6164), .D(w5241), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5313 (.nQ(w6166), .D(w5234), .nC(nDCLK2), .C(DCLK2) );
	vdp_and g5314 (.Z(w5236), .B(w6165), .A(w5244) );
	vdp_and g5315 (.Z(w5237), .B(w6166), .A(DCLK1) );
	vdp_and g5316 (.Z(w5221), .B(w5277), .A(DCLK1) );
	vdp_and g5317 (.Z(w5216), .B(w5274), .A(w5244) );
	vdp_and g5318 (.Z(w5198), .B(w5279), .A(w5278) );
	vdp_and g5319 (.Z(w5199), .B(w71), .A(w5279) );
	vdp_and g5320 (.Z(w5200), .B(w72), .A(w5278) );
	vdp_and g5321 (.Z(w5201), .B(w71), .A(w72) );
	vdp_and g5322 (.Z(w5214), .B(w6216), .A(w5244) );
	vdp_and g5323 (.Z(w5233), .B(w5290), .A(DCLK1) );
	vdp_and g5324 (.Z(w5223), .B(w5304), .A(DCLK1) );
	vdp_and g5325 (.Z(w5197), .B(w5306), .A(w5244) );
	vdp_sr_bit g5326 (.Q(w5282), .D(w5285), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5327 (.Q(w5293), .D(w5263), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_not g5328 (.nZ(w5204), .A(w5211) );
	vdp_not g5329 (.nZ(w5209), .A(w111) );
	vdp_not g5330 (.nZ(w5278), .A(w71) );
	vdp_not g5331 (.nZ(w5279), .A(w72) );
	vdp_aoi21 g5332 (.Z(w5234), .B(w5247), .A1(w5235), .A2(w5236) );
	vdp_aoi21 g5333 (.Z(w5217), .B(w5247), .A1(w5218), .A2(w5216) );
	vdp_aoi21 g5334 (.Z(w6198), .B(w5289), .A1(w5213), .A2(w5214) );
	vdp_oai21 g5335 (.Z(w5211), .B(DCLK2), .A1(w5294), .A2(w5293) );
	vdp_aoi21 g5336 (.Z(w6197), .B(w5289), .A1(w5197), .A2(w5240) );
	vdp_not g5337 (.nZ(w5202), .A(w112) );
	vdp_nand g5338 (.Z(w5263), .B(w5301), .A(w5209) );
	vdp_sr_bit g5339 (.Q(w5254), .D(w5310), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5340 (.Q(w5259), .D(w6167), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5341 (.Q(w5270), .D(w6218), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5342 (.Q(w5255), .D(w5272), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5343 (.Q(w5276), .D(w2610), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5344 (.Q(w5280), .D(w5281), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5345 (.Q(w6209), .D(w5297), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5346 (.Q(w5297), .D(w5309), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5347 (.Q(w5311), .D(w5112), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g5348 (.Z(w5309), .B2(w5112), .B1(w5315), .A1(w5314), .A2(w5311) );
	vdp_aon22 g5349 (.Z(w5281), .B2(w5285), .B1(w5315), .A1(w5314), .A2(w5282) );
	vdp_aon22 g5350 (.Z(w5272), .B2(w5143), .B1(w5315), .A1(w5314), .A2(w5273) );
	vdp_aon22 g5351 (.Z(w5310), .B2(w5179), .B1(w5315), .A1(w5314), .A2(w6219) );
	vdp_not g5352 (.nZ(w5253), .A(w5307) );
	vdp_not g5353 (.nZ(w5245), .A(w72) );
	vdp_not g5354 (.nZ(w5250), .A(w5327) );
	vdp_not g5355 (.nZ(w5258), .A(M5) );
	vdp_not g5356 (.nZ(w5261), .A(w5262) );
	vdp_not g5357 (.nZ(w5248), .A(w5319) );
	vdp_not g5358 (.nZ(w5242), .A(w5317) );
	vdp_not g5359 (.nZ(w5291), .A(w5288) );
	vdp_not g5360 (.nZ(w5308), .A(w5296) );
	vdp_not g5361 (.nZ(w5302), .A(w5297) );
	vdp_comp_we g5362 (.nZ(w5315), .A(M5), .Z(w5314) );
	vdp_and g5363 (.Z(w2728), .B(w5255), .A(w5254) );
	vdp_or g5364 (.Z(w6167), .B(w5254), .A(w5258) );
	vdp_or g5365 (.Z(w5264), .B(w5267), .A(w5263) );
	vdp_and g5366 (.Z(w6218), .B(w5255), .A(M5) );
	vdp_and g5367 (.Z(w2610), .B(w5280), .A(M5) );
	vdp_or g5368 (.Z(w5305), .B(w5263), .A(w5295) );
	vdp_not g5369 (.nZ(w5326), .A(SPR_PRIO) );
	vdp_bufif0 g5370 (.A(w6209), .Z(COL[0]), .nE(w5326) );
	vdp_oai21 g5371 (.Z(w5288), .B(DCLK2), .A1(w5264), .A2(w5287) );
	vdp_bufif0 g5372 (.A(w5276), .Z(COL[6]), .nE(w5326) );
	vdp_bufif0 g5373 (.A(w5270), .Z(COL[5]), .nE(w5326) );
	vdp_bufif0 g5374 (.A(w5259), .Z(COL[4]), .nE(w5326) );
	vdp_oai21 g5375 (.Z(w5262), .B(DCLK2), .A1(w5264), .A2(w5249) );
	vdp_oai21 g5376 (.Z(w5327), .B(DCLK2), .A1(w5321), .A2(w5249) );
	vdp_and3 g5377 (.Z(w5249), .B(w5325), .A(w5248), .C(w5324) );
	vdp_and3 g5378 (.Z(w5267), .B(w5325), .A(w5248), .C(w5312) );
	vdp_and3 g5379 (.Z(w5287), .B(w5324), .A(w5313), .C(w5248) );
	vdp_and3 g5380 (.Z(w5295), .B(w5312), .A(w5313), .C(w5248) );
	vdp_or4 g5381 (.Z(w2609), .B(w5316), .A(w5299), .D(w5297), .C(w5298) );
	vdp_and4 g5382 (.Z(w2668), .B(w5298), .A(w5316), .D(w5302), .C(w5299) );
	vdp_and4 g5383 (.Z(w2667), .B(w5298), .A(w5316), .D(w5297), .C(w5299) );
	vdp_oai21 g5384 (.Z(w5296), .B(DCLK2), .A1(w5287), .A2(w5305) );
	vdp_nand3 g5385 (.Z(w5241), .B(w5242), .A(w5253), .C(w5323) );
	vdp_nand3 g5386 (.Z(w5246), .B(w5322), .A(w102), .C(w5245) );
	vdp_nand3 g5387 (.Z(w5286), .B(w71), .A(w102), .C(w5245) );
	vdp_nand g5388 (.Z(w5289), .B(w5286), .A(w5320) );
	vdp_nand g5389 (.Z(w5283), .B(w5318), .A(w5317) );
	vdp_nand g5390 (.Z(w5284), .B(w5253), .A(w5283) );
	vdp_nand g5391 (.Z(w5275), .B(w5242), .A(w5253) );
	vdp_nand g5392 (.Z(w5247), .B(w5246), .A(w5320) );
	vdp_sr_bit g5393 (.Q(w6170), .D(w6169), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5394 (.Q(w6171), .D(w6170), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5395 (.Q(w5391), .D(w6171), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5396 (.Q(w5398), .D(w5391), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5397 (.Q(w5300), .D(w6172), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5398 (.Q(w6217), .D(w5399), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5399 (.Q(w5492), .D(w6228), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5400 (.Q(w5382), .D(w6168), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_dlatch_inv g5401 (.nQ(w5349), .D(w5341), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5402 (.nQ(w5354), .D(w5340), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5403 (.nQ(w5360), .D(w5339), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5404 (.nQ(w5365), .D(w5338), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5405 (.nQ(w5366), .D(w5337), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5406 (.nQ(w5369), .D(w5336), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5407 (.nQ(w5370), .D(w5335), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5408 (.nQ(w5373), .D(w5333), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5409 (.nQ(w5395), .D(w5396), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5410 (.nQ(w5393), .D(w5378), .nC(nDCLK1), .C(DCLK1) );
	vdp_cnt_bit_load g5411 (.Q(w5396), .D(w5397), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1), .R(1'b0), .CI(w6230), .L(w5330), .nL(w5375) );
	vdp_cnt_bit_load g5412 (.Q(w5378), .D(w5377), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1), .R(1'b0), .CI(w5331), .L(w5330), .nL(w5375), .CO(w6230) );
	vdp_aon22 g5413 (.Z(w5265), .B2(w5332), .B1(DB[11]), .A1(w5373), .A2(w5350) );
	vdp_aon22 g5414 (.Z(w5333), .B2(w5334), .B1(w5362), .A1(w5361), .A2(w5353) );
	vdp_aon22 g5415 (.Z(w5268), .B2(w5332), .B1(DB[12]), .A1(w5370), .A2(w5350) );
	vdp_aon22 g5416 (.Z(w5335), .B2(w5334), .B1(w5358), .A1(w5359), .A2(w5353) );
	vdp_aon22 g5417 (.Z(w5269), .B2(w5332), .B1(DB[13]), .A1(w5369), .A2(w5350) );
	vdp_aon22 g5418 (.Z(w5336), .B2(w5334), .B1(w5351), .A1(w5352), .A2(w5353) );
	vdp_aon22 g5419 (.Z(w5271), .B2(w5332), .B1(DB[14]), .A1(w5366), .A2(w5350) );
	vdp_aon22 g5420 (.Z(w5337), .B2(w5334), .B1(w5342), .A1(w5343), .A2(w5353) );
	vdp_aon22 g5421 (.Z(w5252), .B2(w5332), .B1(DB[3]), .A1(w5365), .A2(w5350) );
	vdp_aon22 g5422 (.Z(w5338), .B2(w5334), .B1(w5361), .A1(w5362), .A2(w5353) );
	vdp_aon22 g5423 (.Z(w5256), .B2(w5332), .B1(DB[4]), .A1(w5360), .A2(w5350) );
	vdp_aon22 g5424 (.Z(w5339), .B2(w5334), .B1(w5359), .A1(w5358), .A2(w5353) );
	vdp_aon22 g5425 (.Z(w5257), .B2(w5332), .B1(DB[5]), .A1(w5354), .A2(w5350) );
	vdp_aon22 g5426 (.Z(w5340), .B2(w5334), .B1(w5352), .A1(w5351), .A2(w5353) );
	vdp_aon22 g5427 (.Z(w5260), .B2(w5332), .B1(DB[6]), .A1(w5349), .A2(w5350) );
	vdp_aon22 g5428 (.Z(w5341), .B2(w5334), .B1(w5343), .A1(w5342), .A2(w5353) );
	vdp_slatch g5429 (.Q(w6168), .D(w5385), .nC(w5329), .C(w5386) );
	vdp_dlatch_inv g5430 (.nQ(w5383), .D(w5382), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5431 (.nQ(w5399), .D(w25), .nC(nHCLK1), .C(HCLK1) );
	vdp_xnor g5432 (.Z(w5313), .B(1'b0), .A(w5393) );
	vdp_xor g5433 (.Z(w5374), .B(w5382), .A(w5384) );
	vdp_aon22 g5434 (.Z(w6228), .B2(w5391), .B1(M5), .A1(w5398), .A2(w6229) );
	vdp_not g5435 (.nZ(w5400), .A(w5399) );
	vdp_not g5436 (.nZ(w6229), .A(M5) );
	vdp_not g5437 (.nZ(w5329), .A(w5386) );
	vdp_not g5438 (.nZ(w6169), .A(w5389) );
	vdp_not g5439 (.nZ(w5312), .A(w5383) );
	vdp_not g5440 (.nZ(w5319), .A(w5395) );
	vdp_not g5441 (.nZ(w5331), .A(w5386) );
	vdp_comp_we g5442 (.nZ(w5350), .A(w111), .Z(w5332) );
	vdp_comp_we g5443 (.nZ(w5353), .A(w5374), .Z(w5334) );
	vdp_comp_we g5444 (.nZ(w5375), .A(w5386), .Z(w5330) );
	vdp_and g5445 (.Z(w6172), .B(w6217), .A(w5400) );
	vdp_aoi21 g5446 (.Z(w5389), .B(w24), .A1(M5), .A2(w21) );
	vdp_sr_bit g5447 (.Q(w5384), .D(w5444), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_aon22 g5448 (.Z(w5451), .B2(w5446), .B1(w5445), .A1(w5442), .A2(w5392) );
	vdp_aon22 g5449 (.Z(w5450), .B2(w5446), .B1(w5448), .A1(w5447), .A2(w5392) );
	vdp_aon22 g5450 (.Z(w5453), .B2(w5446), .B1(w5447), .A1(w5448), .A2(w5392) );
	vdp_aon22 g5451 (.Z(w5452), .B2(w5446), .B1(w5442), .A1(w5445), .A2(w5392) );
	vdp_not g5452 (.nZ(w5409), .A(w5445) );
	vdp_not g5453 (.nZ(w5410), .A(w5448) );
	vdp_not g5454 (.nZ(w5415), .A(w5447) );
	vdp_not g5455 (.nZ(w5414), .A(w5442) );
	vdp_not g5456 (.nZ(w5345), .A(w5450) );
	vdp_not g5457 (.nZ(w5346), .A(w5451) );
	vdp_not g5458 (.nZ(w5347), .A(w5452) );
	vdp_not g5459 (.nZ(w5348), .A(w5453) );
	vdp_not g5460 (.nZ(w5390), .A(M5) );
	vdp_comp_we g5461 (.nZ(w5446), .A(w5384), .Z(w5392) );
	vdp_not g5462 (.nZ(w5386), .A(w5443) );
	vdp_not g5463 (.nZ(w5441), .A(w5440) );
	vdp_dlatch_inv g5464 (.nQ(w5440), .D(w5439), .nC(nHCLK1), .C(HCLK1) );
	vdp_aon2222 g5465 (.Z(w5344), .B2(w5346), .B1(w5403), .A1(w5402), .A2(w5345), .D2(w5348), .D1(w5420), .C1(w5419), .C2(w5347) );
	vdp_aon2222 g5466 (.Z(w5394), .B2(w5415), .B1(w5407), .A1(w5414), .A2(w5402), .D2(w5409), .D1(w5411), .C1(w5410), .C2(w5454) );
	vdp_aon2222 g5467 (.Z(w5364), .B2(w5346), .B1(w5408), .A1(w5407), .A2(w5345), .D2(w5348), .D1(w5412), .C1(w5455), .C2(w5347) );
	vdp_aon2222 g5468 (.Z(w5355), .B2(w5415), .B1(w5408), .A1(w5414), .A2(w5403), .D2(w5409), .D1(w5422), .C1(w5410), .C2(w5416) );
	vdp_aon2222 g5469 (.Z(w5372), .B2(w5346), .B1(w5416), .A1(w5454), .A2(w5345), .D2(w5348), .D1(w5418), .C1(w5417), .C2(w5347) );
	vdp_aon2222 g5470 (.Z(w5363), .B2(w5415), .B1(w5455), .A1(w5414), .A2(w5419), .D2(w5409), .D1(w5421), .C1(w5410), .C2(w5417) );
	vdp_aon2222 g5471 (.Z(w6196), .B2(w5346), .B1(w5422), .A1(w5411), .A2(w5345), .D2(w5348), .D1(w5423), .C1(w5421), .C2(w5347) );
	vdp_aon2222 g5472 (.Z(w5367), .B2(w5415), .B1(w5412), .A1(w5414), .A2(w5420), .D2(w5409), .D1(w5423), .C1(w5410), .C2(w5418) );
	vdp_aon2222 g5473 (.Z(w5356), .B2(w5346), .B1(w5425), .A1(w5424), .A2(w5345), .D2(w5348), .D1(w5437), .C1(w5426), .C2(w5347) );
	vdp_aon2222 g5474 (.Z(w5371), .B2(w5415), .B1(w5427), .A1(w5414), .A2(w5424), .D2(w5409), .D1(w5428), .C1(w5410), .C2(w5429) );
	vdp_aon2222 g5475 (.Z(w5368), .B2(w5346), .B1(w5431), .A1(w5427), .A2(w5345), .D2(w5348), .D1(w5430), .C1(w5432), .C2(w5347) );
	vdp_aon2222 g5476 (.Z(w5380), .B2(w5415), .B1(w5431), .A1(w5414), .A2(w5425), .D2(w5409), .D1(w5433), .C1(w5410), .C2(w5434) );
	vdp_aon2222 g5477 (.Z(w5379), .B2(w5346), .B1(w5434), .A1(w5429), .A2(w5345), .D2(w5348), .D1(w5435), .C1(w5436), .C2(w5347) );
	vdp_aon2222 g5478 (.Z(w5381), .B2(w5415), .B1(w5432), .A1(w5414), .A2(w5426), .D2(w5409), .D1(w5438), .C1(w5410), .C2(w5436) );
	vdp_aon2222 g5479 (.Z(w5388), .B2(w5346), .B1(w5433), .A1(w5428), .A2(w5345), .D2(w5348), .D1(w5449), .C1(w5438), .C2(w5347) );
	vdp_aon2222 g5480 (.Z(w5387), .B2(w5415), .B1(w5430), .A1(w5414), .A2(w5437), .D2(w5409), .D1(w5449), .C1(w5410), .C2(w5435) );
	vdp_aoi22 g5481 (.Z(w5342), .B2(w5401), .B1(w5344), .A1(w5357), .A2(w5394) );
	vdp_aoi22 g5482 (.Z(w5351), .B2(w5401), .B1(w5356), .A1(w5357), .A2(w5355) );
	vdp_aoi22 g5483 (.Z(w5358), .B2(w5401), .B1(w5364), .A1(w5357), .A2(w5363) );
	vdp_aoi22 g5484 (.Z(w5362), .B2(w5401), .B1(w5368), .A1(w5357), .A2(w5367) );
	vdp_aoi22 g5485 (.Z(w5343), .B2(w5401), .B1(w5372), .A1(w5357), .A2(w5371) );
	vdp_aoi22 g5486 (.Z(w5352), .B2(w5401), .B1(w5379), .A1(w5357), .A2(w5380) );
	vdp_aoi22 g5487 (.Z(w5359), .B2(w5401), .B1(w6196), .A1(w5357), .A2(w5381) );
	vdp_aoi22 g5488 (.Z(w5361), .B2(w5401), .B1(w5388), .A1(w5357), .A2(w5387) );
	vdp_nand g5489 (.Z(w5443), .B(w5441), .A(HCLK2) );
	vdp_nor g5490 (.Z(w5401), .B(w5390), .A(w5300) );
	vdp_nor g5491 (.Z(w5357), .B(M5), .A(w5300) );
	vdp_sr_bit g5492 (.Q(w5445), .D(w5448), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5493 (.Q(w5448), .D(w5447), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5494 (.Q(w5447), .D(w5442), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5495 (.Q(w5442), .D(w5443), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_dlatch_inv g5496 (.nQ(w5294), .D(w5445), .nC(nDCLK1), .C(DCLK1) );
	vdp_comp_str g5497 (.nZ(w5406), .A(w5456), .Z(w5458) );
	vdp_comp_str g5498 (.nZ(w5405), .A(w5456), .Z(w5461) );
	vdp_comp_str g5499 (.nZ(w5413), .A(w5456), .Z(w5462) );
	vdp_comp_str g5500 (.nZ(w5404), .A(w5456), .Z(w5457) );
	vdp_slatch g5501 (.D(w5471), .Q(w5402), .nC(w5404), .C(w5457) );
	vdp_slatch g5502 (.D(w6254), .Q(w5403), .nC(w5413), .C(w5462) );
	vdp_slatch g5503 (.D(w6253), .Q(w5419), .nC(w5405), .C(w5461) );
	vdp_slatch g5504 (.D(w6252), .Q(w5420), .nC(w5406), .C(w5458) );
	vdp_slatch g5505 (.D(w5470), .Q(w5407), .nC(w5404), .C(w5457) );
	vdp_slatch g5506 (.D(w6251), .Q(w5408), .nC(w5413), .C(w5462) );
	vdp_slatch g5507 (.D(w6250), .Q(w5455), .nC(w5405), .C(w5461) );
	vdp_slatch g5508 (.D(w6249), .Q(w5412), .nC(w5406), .C(w5458) );
	vdp_slatch g5509 (.D(w5469), .Q(w5454), .nC(w5404), .C(w5457) );
	vdp_slatch g5510 (.D(w6248), .Q(w5416), .nC(w5413), .C(w5462) );
	vdp_slatch g5511 (.D(w6247), .Q(w5417), .nC(w5405), .C(w5461) );
	vdp_slatch g5512 (.D(w6246), .Q(w5418), .nC(w5406), .C(w5458) );
	vdp_slatch g5513 (.D(w5468), .Q(w5411), .nC(w5404), .C(w5457) );
	vdp_slatch g5514 (.D(w6245), .Q(w5422), .nC(w5413), .C(w5462) );
	vdp_slatch g5515 (.D(w6244), .Q(w5421), .nC(w5405), .C(w5461) );
	vdp_slatch g5516 (.D(w6243), .Q(w5423), .nC(w5406), .C(w5458) );
	vdp_slatch g5517 (.D(w5467), .Q(w5424), .nC(w5404), .C(w5457) );
	vdp_slatch g5518 (.D(w6242), .Q(w5425), .nC(w5413), .C(w5462) );
	vdp_slatch g5519 (.D(w6241), .Q(w5426), .nC(w5405), .C(w5461) );
	vdp_slatch g5520 (.D(w6240), .Q(w5437), .nC(w5406), .C(w5458) );
	vdp_slatch g5521 (.D(w5466), .Q(w5427), .nC(w5404), .C(w5457) );
	vdp_slatch g5522 (.D(w6239), .Q(w5431), .nC(w5413), .C(w5462) );
	vdp_slatch g5523 (.D(w6238), .Q(w5432), .nC(w5405), .C(w5461) );
	vdp_slatch g5524 (.D(w6237), .Q(w5430), .nC(w5406), .C(w5458) );
	vdp_slatch g5525 (.D(w5465), .Q(w5429), .nC(w5404), .C(w5457) );
	vdp_slatch g5526 (.D(w6236), .Q(w5434), .nC(w5413), .C(w5462) );
	vdp_slatch g5527 (.D(w6235), .Q(w5436), .nC(w5405), .C(w5461) );
	vdp_slatch g5528 (.D(w6234), .Q(w5435), .nC(w5406), .C(w5458) );
	vdp_slatch g5529 (.D(w5464), .Q(w5428), .nC(w5404), .C(w5457) );
	vdp_slatch g5530 (.D(w6233), .Q(w5433), .nC(w5413), .C(w5462) );
	vdp_slatch g5531 (.D(w6232), .Q(w5438), .nC(w5405), .C(w5461) );
	vdp_slatch g5532 (.D(w6231), .nC(w5406), .C(w5458), .Q(w5449) );
	vdp_sr_bit g5533 (.Q(w5472), .D(w5473), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g5534 (.Q(w6173), .D(w5472), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g5535 (.Q(w5485), .D(w6173), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_comp_str g5536 (.nZ(w5475), .A(w5486), .Z(w5463) );
	vdp_comp_str g5537 (.nZ(w5478), .A(w5486), .Z(w5460) );
	vdp_comp_str g5538 (.nZ(w5480), .A(w5486), .Z(w5459) );
	vdp_dlatch_inv g5539 (.nQ(w5473), .D(w5481), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g5540 (.Z(w5456), .B(DCLK2), .A(w5485) );
	vdp_and g5541 (.Z(w5486), .B(DCLK2), .A(w5472) );
	vdp_and g5542 (.Z(w5487), .B(DCLK2), .A(w5473) );
	vdp_slatch g5543 (.Q(w6233), .D(w6257), .nC(w5475), .C(w5463) );
	vdp_slatch g5544 (.Q(w6232), .D(w6256), .nC(w5478), .C(w5460) );
	vdp_slatch g5545 (.Q(w6231), .D(w6255), .nC(w5480), .C(w5459) );
	vdp_slatch g5546 (.Q(w6236), .D(w6260), .nC(w5475), .C(w5463) );
	vdp_slatch g5547 (.Q(w6235), .D(w6259), .nC(w5478), .C(w5460) );
	vdp_slatch g5548 (.Q(w6234), .D(w6258), .nC(w5480), .C(w5459) );
	vdp_slatch g5549 (.Q(w6239), .D(w6263), .nC(w5475), .C(w5463) );
	vdp_slatch g5550 (.Q(w6238), .D(w6262), .nC(w5478), .C(w5460) );
	vdp_slatch g5551 (.Q(w6237), .D(w6261), .nC(w5480), .C(w5459) );
	vdp_slatch g5552 (.Q(w6242), .D(w6266), .nC(w5475), .C(w5463) );
	vdp_slatch g5553 (.Q(w6241), .D(w6265), .nC(w5478), .C(w5460) );
	vdp_slatch g5554 (.Q(w6240), .D(w6264), .nC(w5480), .C(w5459) );
	vdp_slatch g5555 (.Q(w6245), .D(w6269), .nC(w5475), .C(w5463) );
	vdp_slatch g5556 (.Q(w6244), .D(w6268), .nC(w5478), .C(w5460) );
	vdp_slatch g5557 (.Q(w6243), .D(w6267), .nC(w5480), .C(w5459) );
	vdp_slatch g5558 (.Q(w6248), .D(w6272), .nC(w5475), .C(w5463) );
	vdp_slatch g5559 (.Q(w6247), .D(w6271), .nC(w5478), .C(w5460) );
	vdp_slatch g5560 (.Q(w6246), .D(w6270), .nC(w5480), .C(w5459) );
	vdp_slatch g5561 (.Q(w6251), .D(w6275), .nC(w5475), .C(w5463) );
	vdp_slatch g5562 (.Q(w6250), .D(w6274), .nC(w5478), .C(w5460) );
	vdp_slatch g5563 (.Q(w6249), .D(w6273), .nC(w5480), .C(w5459) );
	vdp_slatch g5564 (.Q(w6254), .D(w6278), .nC(w5475), .C(w5463) );
	vdp_slatch g5565 (.Q(w6253), .D(w6277), .nC(w5478), .C(w5460) );
	vdp_slatch g5566 (.Q(w6252), .D(w6276), .nC(w5480), .C(w5459) );
	vdp_sr_bit g5567 (.Q(w5484), .D(w5483), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_dlatch_inv g5568 (.nQ(w5483), .D(w5482), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g5569 (.Z(w5494), .B(w5483), .A(DCLK2) );
	vdp_nand g5570 (.Z(w5482), .B(w5391), .A(HCLK1) );
	vdp_nand g5571 (.Z(w5481), .B(w5492), .A(HCLK1) );
	vdp_and g5572 (.Z(w5493), .B(w5484), .A(DCLK2) );
	vdp_comp_str g5573 (.nZ(w5479), .A(w5494), .Z(w5491) );
	vdp_comp_str g5574 (.nZ(w5477), .A(w5493), .Z(w5490) );
	vdp_comp_str g5575 (.nZ(w5476), .A(w5487), .Z(w5489) );
	vdp_comp_str g5576 (.nZ(w5474), .A(w5486), .Z(w5488) );
	vdp_slatch g5577 (.D(S[7]), .Q(w5471), .nC(w5474), .C(w5488) );
	vdp_slatch g5578 (.D(S[7]), .Q(w6278), .nC(w5476), .C(w5489) );
	vdp_slatch g5579 (.D(S[7]), .Q(w6277), .nC(w5477), .C(w5490) );
	vdp_slatch g5580 (.D(S[7]), .Q(w6276), .nC(w5479), .C(w5491) );
	vdp_slatch g5581 (.D(S[5]), .Q(w5470), .nC(w5474), .C(w5488) );
	vdp_slatch g5582 (.D(S[5]), .Q(w6275), .nC(w5476), .C(w5489) );
	vdp_slatch g5583 (.D(S[5]), .Q(w6274), .nC(w5477), .C(w5490) );
	vdp_slatch g5584 (.D(S[5]), .Q(w6273), .nC(w5479), .C(w5491) );
	vdp_slatch g5585 (.D(S[3]), .Q(w5469), .nC(w5474), .C(w5488) );
	vdp_slatch g5586 (.D(S[3]), .Q(w6272), .nC(w5476), .C(w5489) );
	vdp_slatch g5587 (.D(S[3]), .Q(w6271), .nC(w5477), .C(w5490) );
	vdp_slatch g5588 (.D(S[3]), .Q(w6270), .nC(w5479), .C(w5491) );
	vdp_slatch g5589 (.D(S[1]), .Q(w5468), .nC(w5474), .C(w5488) );
	vdp_slatch g5590 (.D(S[1]), .Q(w6269), .nC(w5476), .C(w5489) );
	vdp_slatch g5591 (.D(S[1]), .Q(w6268), .nC(w5477), .C(w5490) );
	vdp_slatch g5592 (.D(S[1]), .Q(w6267), .nC(w5479), .C(w5491) );
	vdp_slatch g5593 (.D(S[6]), .Q(w5467), .nC(w5474), .C(w5488) );
	vdp_slatch g5594 (.D(S[6]), .Q(w6266), .nC(w5476), .C(w5489) );
	vdp_slatch g5595 (.D(S[6]), .Q(w6265), .nC(w5477), .C(w5490) );
	vdp_slatch g5596 (.D(S[6]), .Q(w6264), .nC(w5479), .C(w5491) );
	vdp_slatch g5597 (.D(S[4]), .Q(w5466), .nC(w5474), .C(w5488) );
	vdp_slatch g5598 (.D(S[4]), .Q(w6263), .nC(w5476), .C(w5489) );
	vdp_slatch g5599 (.D(S[4]), .Q(w6262), .nC(w5477), .C(w5490) );
	vdp_slatch g5600 (.D(S[4]), .Q(w6261), .nC(w5479), .C(w5491) );
	vdp_slatch g5601 (.D(S[2]), .Q(w5465), .nC(w5474), .C(w5488) );
	vdp_slatch g5602 (.D(S[2]), .Q(w6260), .nC(w5476), .C(w5489) );
	vdp_slatch g5603 (.D(S[2]), .Q(w6259), .nC(w5477), .C(w5490) );
	vdp_slatch g5604 (.D(S[2]), .Q(w6258), .nC(w5479), .C(w5491) );
	vdp_slatch g5605 (.D(S[0]), .Q(w5464), .nC(w5474), .C(w5488) );
	vdp_slatch g5606 (.D(S[0]), .Q(w6257), .nC(w5476), .C(w5489) );
	vdp_slatch g5607 (.D(S[0]), .Q(w6256), .nC(w5477), .C(w5490) );
	vdp_slatch g5608 (.D(S[0]), .nC(w5479), .C(w5491), .Q(w6255) );
	vdp_aon21_sr g5609 (.Q(w5548), .A1(w5120), .A2(w6439), .B(w6592), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5610 (.Q(w6592), .A1(w5117), .A2(w6439), .B(w6593), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5611 (.Q(w6593), .A1(w5115), .A2(w6439), .B(w6594), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5612 (.Q(w6594), .A1(w5533), .A2(w6439), .B(w6595), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5613 (.Q(w6595), .A1(w5543), .A2(w6439), .B(w6596), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5614 (.Q(w6596), .A1(w5510), .A2(w6439), .B(w6597), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5615 (.Q(w6597), .A1(w5512), .A2(w6439), .B(w6598), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5616 (.Q(w6598), .A1(w5502), .A2(w6439), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5617 (.Q(w6599), .A1(w5507), .A2(w6440), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5618 (.Q(w6600), .A1(w5513), .A2(w6440), .B(w6599), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5619 (.Q(w6601), .A1(w5511), .A2(w6440), .B(w6600), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5620 (.Q(w6602), .A1(w5550), .A2(w6440), .B(w6601), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5621 (.Q(w6603), .A1(w5534), .A2(w6440), .B(w6602), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5622 (.Q(w6604), .A1(w5116), .A2(w6440), .B(w6603), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5623 (.Q(w6605), .A1(w5118), .A2(w6440), .B(w6604), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5624 (.Q(w5553), .A1(w5119), .A2(w6440), .B(w6605), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5625 (.Q(w5558), .A1(w5504), .A2(w6441), .B(w6606), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5626 (.Q(w6606), .A1(w5501), .A2(w6441), .B(w6607), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5627 (.Q(w6607), .A1(w5500), .A2(w6441), .B(w6608), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5628 (.Q(w6608), .A1(w5506), .A2(w6441), .B(w6609), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5629 (.Q(w6609), .A1(w5509), .A2(w6441), .B(w6610), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5630 (.Q(w6610), .A1(w5514), .A2(w6441), .B(w6611), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5631 (.Q(w6611), .A1(w5526), .A2(w6441), .B(w6612), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5632 (.Q(w6612), .A1(w5529), .A2(w6441), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_or4 g5633 (.Z(w5539), .B(w5543), .A(w5191), .C(w5550), .D(w5509) );
	vdp_or4 g5634 (.Z(w5194), .B(w5533), .A(w5189), .C(w5534), .D(w5506) );
	vdp_aon22 g5635 (.Z(w5522), .B2(w4360), .B1(w5527), .A1(w5563), .A2(DB[0]) );
	vdp_aon22 g5636 (.Z(w5521), .B2(w4361), .B1(w5527), .A1(w5563), .A2(DB[1]) );
	vdp_aon22 g5637 (.Z(w5520), .B2(w4369), .B1(w5527), .A1(w5563), .A2(DB[2]) );
	vdp_aon22 g5638 (.Z(w5519), .B2(w4360), .B1(w5527), .A1(w5563), .A2(DB[8]) );
	vdp_aon22 g5639 (.Z(w5518), .B2(w4361), .B1(w5527), .A1(w5563), .A2(DB[9]) );
	vdp_aon22 g5640 (.Z(w5517), .B2(w4369), .B1(w5527), .A1(w5563), .A2(DB[10]) );
	vdp_or4 g5641 (.Z(w5549), .B(w5498), .A(w5499), .C(w5531), .D(w5532) );
	vdp_or4 g5642 (.Z(w5540), .B(w5537), .A(w5538), .C(w5536), .D(w5535) );
	vdp_or4 g5643 (.Z(w5557), .B(w5512), .A(w5183), .C(w5513), .D(w5526) );
	vdp_or4 g5644 (.Z(w5554), .B(w5511), .A(w5514), .C(w5510), .D(w5508) );
	vdp_or4 g5645 (.Z(w5564), .B(w5503), .A(w5505), .C(w5516), .D(w5515) );
	vdp_or4 g5646 (.Z(w5555), .B(w5524), .A(w5525), .C(w5530), .D(w5523) );
	vdp_or4 g5647 (.Z(w5566), .B(w5502), .A(w5184), .C(w5507), .D(w5529) );
	vdp_comp_we g5648 (.nZ(w5527), .A(w111), .Z(w5563) );
	vdp_not g5649 (.nZ(w6439), .A(nSRLOAD) );
	vdp_not g5650 (.nZ(w6440), .A(nSRLOAD) );
	vdp_not g5651 (.nZ(w6441), .A(nSRLOAD) );
	vdp_slatch g5652 (.Q(w5535), .D(w5580), .nC(w5546), .C(w5579) );
	vdp_comp_str g5653 (.nZ(w5546), .A(w5204), .Z(w5579) );
	vdp_slatch g5654 (.Q(w5536), .D(w5582), .nC(w5546), .C(w5579) );
	vdp_slatch g5655 (.Q(w5537), .D(w5583), .nC(w5546), .C(w5579) );
	vdp_slatch g5656 (.Q(w5538), .D(w5584), .nC(w5546), .C(w5579) );
	vdp_slatch g5657 (.Q(w5499), .D(w5585), .nC(w5546), .C(w5579) );
	vdp_slatch g5658 (.Q(w5498), .D(w5587), .nC(w5546), .C(w5579) );
	vdp_slatch g5659 (.Q(w5531), .D(w5588), .nC(w5546), .C(w5579) );
	vdp_slatch g5660 (.Q(w5532), .D(w5589), .nC(w5546), .C(w5579) );
	vdp_slatch g5661 (.Q(w5523), .D(w5598), .nC(w5561), .C(w5597) );
	vdp_comp_str g5662 (.nZ(w5561), .A(w5204), .Z(w5597) );
	vdp_slatch g5663 (.Q(w5530), .D(w5600), .nC(w5561), .C(w5597) );
	vdp_slatch g5664 (.Q(w5524), .D(w5601), .nC(w5561), .C(w5597) );
	vdp_slatch g5665 (.Q(w5525), .D(w5602), .nC(w5561), .C(w5597) );
	vdp_slatch g5666 (.Q(w5505), .D(w5603), .nC(w5561), .C(w5597) );
	vdp_slatch g5667 (.Q(w5503), .D(w5605), .nC(w5561), .C(w5597) );
	vdp_slatch g5668 (.Q(w5516), .D(w5606), .nC(w5561), .C(w5597) );
	vdp_slatch g5669 (.Q(w5515), .D(w5607), .nC(w5561), .C(w5597) );
	vdp_comp_we g5670 (.nZ(w5542), .A(1'b0), .Z(w5192) );
	vdp_aon22 g5671 (.Z(w5609), .B2(w5542), .B1(w5565), .A1(w5564), .A2(w5192) );
	vdp_not g5672 (.nZ(nSRLOAD), .A(w4371) );
	vdp_not g5673 (.nZ(w5565), .A(w5566) );
	vdp_not g5674 (.nZ(w5556), .A(w5557) );
	vdp_not g5675 (.nZ(w5552), .A(w5554) );
	vdp_not g5676 (.nZ(w5541), .A(w5539) );
	vdp_and3 g5677 (.Z(w5569), .B(w5568), .A(w5540), .C(w5539) );
	vdp_aon22 g5678 (.Z(w5577), .B2(w5542), .B1(w5541), .A1(w5540), .A2(w5192) );
	vdp_notif0 g5679 (.A(w5544), .nZ(DB[4]), .nE(w5545) );
	vdp_aon2222 g5680 (.Z(w5544), .B2(w5543), .B1(w5575), .A1(w5576), .A2(w5512), .D2(w5120), .D1(w5573), .C1(w5574), .C2(w5115) );
	vdp_notif0 g5681 (.A(w5547), .nZ(DB[12]), .nE(w5545) );
	vdp_aon2222 g5682 (.Z(w5547), .B2(w5510), .B1(w5575), .A1(w5576), .A2(w5502), .D2(w5117), .D1(w5573), .C1(w5574), .C2(w5533) );
	vdp_notif0 g5683 (.A(w6208), .nZ(DB[13]), .nE(w5545) );
	vdp_aon2222 g5684 (.Z(w6208), .B2(w5511), .B1(w5575), .A1(w5576), .A2(w5507), .D2(w5118), .D1(w5573), .C1(w5574), .C2(w5534) );
	vdp_notif0 g5685 (.A(w5551), .nZ(DB[5]), .nE(w5545) );
	vdp_aon2222 g5686 (.Z(w5551), .B2(w5550), .B1(w5575), .A1(w5576), .A2(w5513), .D2(w5119), .D1(w5573), .C1(w5574), .C2(w5116) );
	vdp_notif0 g5687 (.A(w5560), .nZ(DB[14]), .nE(w5545) );
	vdp_aon2222 g5688 (.Z(w5560), .B2(w5514), .B1(w5575), .A1(w5576), .A2(w5529), .D2(w5501), .D1(w5573), .C1(w5574), .C2(w5506) );
	vdp_notif0 g5689 (.A(w5559), .nZ(DB[6]), .nE(w5545) );
	vdp_aon2222 g5690 (.Z(w5559), .B2(w5509), .B1(w5575), .A1(w5576), .A2(w5526), .D2(w5504), .D1(w5573), .C1(w5574), .C2(w5500) );
	vdp_aon22 g5691 (.Z(w5590), .B2(w5542), .B1(w5552), .A1(w5549), .A2(w5192) );
	vdp_aon22 g5692 (.Z(w5593), .B2(w5542), .B1(w5556), .A1(w5555), .A2(w5192) );
	vdp_and3 g5693 (.Z(w5571), .B(w5592), .A(w5549), .C(w5554) );
	vdp_and3 g5694 (.Z(w5572), .B(w5594), .A(w5555), .C(w5557) );
	vdp_and3 g5695 (.Z(w5570), .B(w5608), .A(w5564), .C(w5566) );
	vdp_not g5696 (.nZ(w5545), .A(w112) );
	vdp_slatch g5697 (.Q(w5603), .D(w5265), .nC(w5637), .C(w5604) );
	vdp_slatch g5698 (.Q(w5605), .D(w5268), .nC(w5637), .C(w5604) );
	vdp_slatch g5699 (.Q(w5606), .D(w5269), .nC(w5637), .C(w5604) );
	vdp_slatch g5700 (.Q(w5607), .D(w5271), .nC(w5637), .C(w5604) );
	vdp_comp_str g5701 (.nZ(w5637), .A(w5638), .Z(w5604) );
	vdp_slatch g5702 (.Q(w5598), .D(w5252), .nC(w5632), .C(w5599) );
	vdp_slatch g5703 (.Q(w5600), .D(w5256), .nC(w5632), .C(w5599) );
	vdp_slatch g5704 (.Q(w5601), .D(w5257), .nC(w5632), .C(w5599) );
	vdp_slatch g5705 (.Q(w5602), .D(w5260), .nC(w5632), .C(w5599) );
	vdp_comp_str g5706 (.nZ(w5632), .A(w5636), .Z(w5599) );
	vdp_slatch g5707 (.Q(w5585), .D(w5265), .nC(w5619), .C(w5586) );
	vdp_slatch g5708 (.Q(w5587), .D(w5268), .nC(w5619), .C(w5586) );
	vdp_slatch g5709 (.Q(w5588), .D(w5269), .nC(w5619), .C(w5586) );
	vdp_slatch g5710 (.Q(w5589), .D(w5271), .nC(w5619), .C(w5586) );
	vdp_comp_str g5711 (.nZ(w5619), .A(w6436), .Z(w5586) );
	vdp_slatch g5712 (.Q(w5580), .D(w5252), .nC(w5618), .C(w5581) );
	vdp_slatch g5713 (.Q(w5582), .D(w5256), .nC(w5618), .C(w5581) );
	vdp_slatch g5714 (.Q(w5583), .D(w5257), .nC(w5618), .C(w5581) );
	vdp_slatch g5715 (.Q(w5584), .D(w5260), .nC(w5618), .C(w5581) );
	vdp_comp_str g5716 (.nZ(w5618), .A(w5616), .Z(w5581) );
	vdp_dlatch_inv g5717 (.nQ(w6207), .D(w5611), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5718 (.Z(w5613), .B(w5243), .A(w6207) );
	vdp_sr_bit g5719 (.Q(COLLISION), .D(w6204), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g5720 (.Q(w5610), .D(w5548), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5721 (.nQ(w5615), .D(w5578), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5722 (.nQ(w6199), .D(w5591), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5723 (.nQ(w6201), .D(w5625), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5724 (.Z(w6200), .B(w6201), .A(w5243) );
	vdp_sr_bit g5725 (.Q(w6210), .D(w5553), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5726 (.nQ(w5595), .D(w6434), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5727 (.Z(w6202), .B(w5595), .A(w5243) );
	vdp_sr_bit g5728 (.Q(w5629), .D(w5558), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5729 (.nQ(w5626), .D(w6206), .nC(nDCLK2), .C(DCLK2) );
	vdp_not g5730 (.nZ(w5642), .A(w5243) );
	vdp_not g5731 (.nZ(w5596), .A(w72) );
	vdp_not g5732 (.nZ(w5630), .A(w71) );
	vdp_dlatch_inv g5733 (.nQ(w5640), .D(w6203), .nC(nDCLK2), .C(DCLK2) );
	vdp_and g5734 (.Z(w5608), .B(w5642), .A(w5244) );
	vdp_aoi21 g5735 (.Z(w6203), .B(w5627), .A1(w5609), .A2(w5608) );
	vdp_and g5736 (.Z(w5495), .B(w5640), .A(DCLK1) );
	vdp_and g5737 (.Z(w5496), .B(w5626), .A(DCLK1) );
	vdp_and g5738 (.Z(w5594), .B(w6202), .A(w5244) );
	vdp_aoi21 g5739 (.Z(w6206), .B(w5627), .A1(w5593), .A2(w5594) );
	vdp_and g5740 (.Z(w5592), .B(w6200), .A(w5244) );
	vdp_aoi21 g5741 (.Z(w5591), .B(w5614), .A1(w5590), .A2(w5592) );
	vdp_and g5742 (.Z(w5568), .B(w5244), .A(w5613) );
	vdp_aoi21 g5743 (.Z(w5578), .B(w5614), .A1(w5577), .A2(w5568) );
	vdp_and g5744 (.Z(w5528), .B(DCLK1), .A(w5615) );
	vdp_and g5745 (.Z(w5497), .B(w6199), .A(DCLK1) );
	vdp_and g5746 (.Z(w5573), .B(w5596), .A(w5630) );
	vdp_and g5747 (.Z(w5575), .B(w72), .A(w5630) );
	vdp_and g5748 (.Z(w5574), .B(w5596), .A(w71) );
	vdp_and g5749 (.Z(w5576), .B(w72), .A(w71) );
	vdp_or8 g5750 (.Z(w6204), .B(w5569), .A(w5238), .C(w5570), .D(w6205), .F(w5572), .E(w5567), .G(w5222), .H(w5571) );
	vdp_sr_bit g5751 (.Q(w5299), .D(w5647), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5752 (.Q(w5612), .D(w5299), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5753 (.Q(w5298), .D(w5624), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5754 (.Q(w5643), .D(w5298), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5755 (.Q(w5316), .D(w6188), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5756 (.Q(w5631), .D(w5316), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_comp_we g5757 (.nZ(w5645), .A(M5), .Z(w5644) );
	vdp_not g5758 (.nZ(w5638), .A(w5639) );
	vdp_or g5759 (.Z(w5321), .B(w5641), .A(w5263) );
	vdp_and3 g5760 (.Z(w5641), .B(w5313), .A(w5319), .C(w5312) );
	vdp_and3 g5761 (.Z(w5634), .B(w5313), .A(w5319), .C(w5324) );
	vdp_and3 g5762 (.Z(w6434), .B(w5317), .A(w5307), .C(w5318) );
	vdp_and3 g5763 (.Z(w5621), .B(w5325), .A(w5319), .C(w5312) );
	vdp_and3 g5764 (.Z(w5623), .B(w5325), .A(w5319), .C(w5324) );
	vdp_aoi21 g5765 (.Z(w5611), .B(w5253), .A1(w5242), .A2(w5323) );
	vdp_aon22 g5766 (.Z(w5647), .B2(w5548), .B1(w5645), .A1(w5644), .A2(w5610) );
	vdp_aon22 g5767 (.Z(w5624), .B2(w5553), .B1(w5645), .A1(w5644), .A2(w6210) );
	vdp_aon22 g5768 (.Z(w6188), .B2(w5558), .B1(w5645), .A1(w5644), .A2(w5629) );
	vdp_bufif0 g5769 (.A(w5643), .Z(COL[2]), .nE(w5646) );
	vdp_oai21 g5770 (.Z(w5622), .B(DCLK2), .A1(w5635), .A2(w5623) );
	vdp_and g5771 (.Z(w5625), .B(w5317), .A(w5307) );
	vdp_or g5772 (.Z(w5635), .B(w5621), .A(w5263) );
	vdp_bufif0 g5773 (.A(w5631), .Z(COL[3]), .nE(w5646) );
	vdp_oai21 g5774 (.Z(w5633), .B(DCLK2), .A1(w5635), .A2(w5634) );
	vdp_oai21 g5775 (.Z(w5639), .B(DCLK2), .A1(w5634), .A2(w5321) );
	vdp_not g5776 (.nZ(w5324), .A(w5312) );
	vdp_not g5777 (.nZ(w5636), .A(w5633) );
	vdp_not g5778 (.nZ(w5322), .A(w71) );
	vdp_not g5779 (.nZ(w5325), .A(w5313) );
	vdp_not g5780 (.nZ(w6436), .A(w5622) );
	vdp_not g5781 (.nZ(w5323), .A(w5318) );
	vdp_not g5782 (.nZ(w5616), .A(w5617) );
	vdp_bufif0 g5783 (.A(w5612), .Z(COL[1]), .nE(w5646) );
	vdp_oai21 g5784 (.Z(w5617), .B(DCLK2), .A1(w5305), .A2(w5623) );
	vdp_not g5785 (.nZ(w5646), .A(SPR_PRIO) );
	vdp_nand3 g5786 (.Z(w5620), .B(w102), .A(w72), .C(w5322) );
	vdp_nand g5787 (.Z(w5614), .B(w5320), .A(w5620) );
	vdp_nand3 g5788 (.Z(w5628), .B(w102), .A(w72), .C(w71) );
	vdp_nand g5789 (.Z(w5627), .B(w5320), .A(w5628) );
	vdp_sr_bit g5790 (.Q(w5670), .D(w5711), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5791 (.Q(w5671), .D(w5709), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5792 (.Q(w5668), .D(w5716), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5793 (.Q(w5669), .D(w5708), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5794 (.Z(w4366), .B2(w5670), .B1(w5705), .A1(w5704), .A2(w70), .C1(w5659), .C2(w5671) );
	vdp_aon222 g5795 (.Z(w4365), .B2(w5668), .B1(w5705), .A1(w5704), .A2(w69), .C1(w5659), .C2(w5669) );
	vdp_sr_bit g5796 (.Q(w5666), .D(w5715), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5797 (.Q(w5667), .D(w5707), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5798 (.Z(w4364), .B2(w5666), .B1(w5705), .A1(w5704), .A2(w68), .C1(w5659), .C2(w5667) );
	vdp_sr_bit g5799 (.Q(w5664), .D(w5714), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5800 (.Q(w5665), .D(w5706), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5801 (.Z(w4363), .B2(w5664), .B1(w5705), .A1(w5704), .A2(w67), .C1(w5659), .C2(w5665) );
	vdp_sr_bit g5802 (.Q(w5660), .D(w5713), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5803 (.Q(w5663), .D(w5717), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5804 (.Z(w4362), .B2(w5660), .B1(w5705), .A1(w5704), .A2(w66), .C1(w5659), .C2(w5663) );
	vdp_sr_bit g5805 (.Q(w5661), .D(w5712), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5806 (.Q(w5662), .D(w5703), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5807 (.Z(w4367), .B2(w5661), .B1(w5705), .A1(w5704), .A2(w65), .C1(w5659), .C2(w5662) );
	vdp_sr_bit g5808 (.Q(w5307), .D(w6413), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_slatch g5809 (.Q(w6413), .D(w5397), .nC(w5695), .C(w5656) );
	vdp_sr_bit g5810 (.Q(w5317), .D(w6411), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_slatch g5811 (.Q(w6411), .D(w5377), .nC(w5695), .C(w5656) );
	vdp_sr_bit g5812 (.Q(w5318), .D(w6412), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_slatch g5813 (.Q(w6412), .D(w5385), .nC(w5695), .C(w5656) );
	vdp_sr_bit g5814 (.Q(w5672), .D(w25), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5815 (.Q(w5655), .D(w5672), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5816 (.Q(w5654), .D(w5700), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5817 (.Q(w5688), .D(w5698), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5818 (.Q(w5687), .D(w5697), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5819 (.Q(w5651), .D(w4371), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5820 (.Q(w5650), .D(w5683), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5821 (.Q(w5678), .D(w6213), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5822 (.Q(w6213), .D(w5719), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_xor g5823 (.Z(w5680), .B(w5678), .A(w5679) );
	vdp_dlatch_inv g5824 (.nQ(w5649), .D(w5683), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5825 (.nQ(w5681), .D(w5680), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5826 (.nQ(w5652), .D(w5653), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5827 (.nQ(w5686), .D(w5685), .nC(nHCLK1), .C(HCLK1) );
	vdp_comp_str g5828 (.nZ(w5695), .A(w5692), .Z(w5656) );
	vdp_oai21 g5829 (.Z(w6212), .B(w5682), .A1(w5719), .A2(w5678) );
	vdp_and g5830 (.Z(w4360), .B(w5676), .A(w5648) );
	vdp_not g5831 (.nZ(w5243), .A(w5681) );
	vdp_not g5832 (.nZ(w5683), .A(w6212) );
	vdp_and g5833 (.Z(w4361), .B(w5675), .A(w5648) );
	vdp_and g5834 (.Z(w4369), .B(w5674), .A(w5648) );
	vdp_or g5835 (.Z(w5684), .B(w5650), .A(w5683) );
	vdp_not g5836 (.nZ(w5702), .A(w111) );
	vdp_not g5837 (.nZ(w4371), .A(w5685) );
	vdp_not g5838 (.nZ(w5718), .A(M5) );
	vdp_not g5839 (.nZ(w5705), .A(w6403) );
	vdp_not g5840 (.nZ(w5657), .A(w5656) );
	vdp_not g5841 (.nZ(w5704), .A(w5702) );
	vdp_not g5842 (.nZ(w5659), .A(w5658) );
	vdp_or4 g5843 (.Z(w4368), .B(w4371), .A(w111), .C(w5651), .D(w5684) );
	vdp_or4 g5844 (.Z(w5685), .B(w5688), .A(w5648), .C(w5654), .D(w5687) );
	vdp_nand g5845 (.Z(w5653), .B(w5686), .A(HCLK2) );
	vdp_nand g5846 (.Z(w5320), .B(w5702), .A(w5652) );
	vdp_nor g5847 (.Z(w5244), .B(w5649), .A(w111) );
	vdp_nand g5848 (.Z(w5658), .B(w5702), .A(w5657) );
	vdp_nand g5849 (.Z(w6403), .B(w5702), .A(w5648) );
	vdp_aoi22 g5850 (.Z(w5648), .B2(w5718), .B1(w25), .A1(M5), .A2(w5655) );
	vdp_cnt_bit_load g5851 (.Q(w5747), .D(w5696), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w35), .CI(w5803), .L(w5694), .nL(w5740) );
	vdp_cnt_bit_load g5852 (.Q(w5693), .D(w5744), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w35), .CI(w5689), .L(w5694), .nL(w5740), .CO(w5803) );
	vdp_sr_bit g5853 (.Q(w5682), .D(w6195), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5854 (.SUM(w5700), .CO(w6391), .CI(1'b1), .A(HPOS[0]), .B(M5) );
	vdp_fa g5855 (.SUM(w5698), .CO(w6392), .CI(w6391), .A(HPOS[1]), .B(1'b0) );
	vdp_fa g5856 (.SUM(w5697), .CO(w6393), .CI(w6392), .A(HPOS[2]), .B(1'b1) );
	vdp_fa g5857 (.SUM(w5703), .CO(w6394), .CI(w6393), .A(HPOS[3]), .B(M5) );
	vdp_fa g5858 (.SUM(w5717), .CO(w6395), .CI(w6394), .A(HPOS[4]), .B(w5755) );
	vdp_fa g5859 (.SUM(w5706), .CO(w6396), .CI(w6395), .A(HPOS[5]), .B(1'b1) );
	vdp_fa g5860 (.SUM(w5707), .CO(w6397), .CI(w6396), .A(HPOS[6]), .B(1'b1) );
	vdp_fa g5861 (.SUM(w5708), .CO(w6398), .CI(w6397), .A(HPOS[7]), .B(1'b1) );
	vdp_fa g5862 (.SUM(w5709), .CI(w6398), .A(HPOS[8]), .B(1'b1) );
	vdp_not g5863 (.nZ(w5755), .A(M5) );
	vdp_aoi33 g5864 (.Z(w6195), .B2(w6410), .B1(w5711), .A1(H40), .A2(w5711), .A3(w5710), .B3(w6410) );
	vdp_not g5865 (.nZ(w6410), .A(H40) );
	vdp_or g5866 (.Z(w5710), .B(w5715), .A(w5716) );
	vdp_and g5867 (.Z(w5691), .B(w5689), .A(w5690) );
	vdp_sr_bit g5868 (.Q(w5689), .D(w6211), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5869 (.Q(w6211), .D(w5439), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5870 (.nQ(w5737), .D(w5294), .nC(nDCLK2), .C(DCLK2) );
	vdp_slatch g5871 (.Q(w5736), .D(w5723), .nC(w5677), .C(w5727) );
	vdp_slatch g5872 (.Q(w5676), .D(w5736), .nC(w5673), .C(w5729) );
	vdp_slatch g5873 (.Q(w5730), .D(w5721), .nC(w5677), .C(w5727) );
	vdp_slatch g5874 (.Q(w5674), .D(w5730), .nC(w5673), .C(w5729) );
	vdp_slatch g5875 (.Q(w5731), .D(w5722), .nC(w5677), .C(w5727) );
	vdp_slatch g5876 (.Q(w5675), .D(w5731), .nC(w5673), .C(w5729) );
	vdp_slatch g5877 (.Q(w6214), .D(w5444), .nC(w5677), .C(w5727) );
	vdp_sr_bit g5878 (.Q(w5679), .D(w6214), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_and g5879 (.Z(w5720), .B(DCLK2), .A(w5294) );
	vdp_comp_str g5880 (.nZ(w5673), .A(w5720), .Z(w5729) );
	vdp_comp_str g5881 (.nZ(w5677), .A(w5692), .Z(w5727) );
	vdp_not g5882 (.nZ(w5719), .A(w5737) );
	vdp_comp_we g5883 (.nZ(w5740), .A(w5691), .Z(w5694) );
	vdp_and3 g5884 (.Z(w5692), .B(HCLK1), .A(w5690), .C(w5689) );
	vdp_nand g5885 (.Z(w5744), .B(w5725), .A(M5) );
	vdp_nand g5886 (.Z(w5696), .B(w5724), .A(M5) );
	vdp_nor g5887 (.Z(w5690), .B(w5747), .A(w5693) );
	vdp_fa g5888 (.SUM(w5711), .CI(w5765), .A(w5764), .B(w5775) );
	vdp_aon22 g5889 (.Z(w5764), .B2(w5767), .B1(w5763), .A1(w5797), .A2(w5733) );
	vdp_sr_bit g5890 (.Q(w5763), .D(w5711), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5891 (.Q(w5797), .D(w5798), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5892 (.SUM(w5798), .CI(w5761), .A(w5762), .B(w5793) );
	vdp_aon22 g5893 (.Z(w5762), .B2(w5772), .B1(w5796), .A1(1'b0), .A2(w5726) );
	vdp_fa g5894 (.SUM(w5716), .CO(w5765), .CI(w5760), .A(w5759), .B(w5775) );
	vdp_aon22 g5895 (.Z(w5759), .B2(w5767), .B1(w5758), .A1(w5794), .A2(w5733) );
	vdp_sr_bit g5896 (.Q(w5758), .D(w5716), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5897 (.Q(w5794), .D(w5800), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5898 (.SUM(w5800), .CO(w5761), .CI(w5757), .A(w5756), .B(w5793) );
	vdp_aon22 g5899 (.Z(w5756), .B2(w5772), .B1(w5791), .A1(w5792), .A2(w5726) );
	vdp_fa g5900 (.SUM(w5715), .CO(w5760), .CI(w5754), .A(w5753), .B(w5775) );
	vdp_aon22 g5901 (.Z(w5753), .B2(w5767), .B1(w5752), .A1(w5790), .A2(w5733) );
	vdp_fa g5902 (.SUM(w5801), .CO(w5757), .CI(w5751), .A(w5750), .B(w5777) );
	vdp_aon22 g5903 (.Z(w5750), .B2(w5772), .B1(w5788), .A1(w5789), .A2(w5726) );
	vdp_sr_bit g5904 (.Q(w5752), .D(w5715), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5905 (.Q(w5790), .D(w5801), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5906 (.SUM(w5714), .CO(w5754), .CI(w5766), .A(w5749), .B(w5775) );
	vdp_aon22 g5907 (.Z(w5749), .B2(w5767), .B1(w5748), .A1(w5787), .A2(w5733) );
	vdp_sr_bit g5908 (.Q(w5748), .D(w5714), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5909 (.Q(w5787), .D(w5786), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5910 (.SUM(w5786), .CO(w5751), .CI(w5745), .A(w5746), .B(w5777) );
	vdp_aon22 g5911 (.Z(w5746), .B2(w5772), .B1(w6407), .A1(w5785), .A2(w5726) );
	vdp_fa g5912 (.SUM(w5713), .CO(w5766), .CI(w5742), .A(w5743), .B(w5775) );
	vdp_aon22 g5913 (.Z(w5743), .B2(w5767), .B1(w5741), .A1(w5784), .A2(w5733) );
	vdp_sr_bit g5914 (.Q(w5741), .D(w5713), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5915 (.Q(w5784), .D(w6399), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5916 (.SUM(w6399), .CO(w5745), .CI(w5739), .A(w5738), .B(w5783) );
	vdp_aon22 g5917 (.Z(w5738), .B2(w5772), .B1(w5802), .A1(w5782), .A2(w5726) );
	vdp_fa g5918 (.SUM(w5712), .CO(w5742), .CI(w5735), .A(w5734), .B(w5775) );
	vdp_aon22 g5919 (.Z(w5734), .B2(w5767), .B1(w5732), .A1(w5781), .A2(w5733) );
	vdp_sr_bit g5920 (.Q(w5732), .D(w5712), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5921 (.Q(w5781), .D(w5780), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5922 (.SUM(w5780), .CO(w5739), .CI(w5444), .A(w5728), .B(w6404) );
	vdp_aon22 g5923 (.Z(w5728), .B2(w5772), .B1(w5778), .A1(w5779), .A2(w5726) );
	vdp_aon22 g5924 (.Z(w5397), .B2(w5772), .B1(w5776), .A1(w5799), .A2(w5726) );
	vdp_aon22 g5925 (.Z(w5377), .B2(w5772), .B1(w5771), .A1(w5774), .A2(w5726) );
	vdp_aon22 g5926 (.Z(w5385), .B2(w5772), .B1(w5770), .A1(w5773), .A2(w5726) );
	vdp_and g5927 (.Z(w5735), .B(w5769), .A(w6406) );
	vdp_comp_we g5928 (.nZ(w5726), .A(M5), .Z(w5772) );
	vdp_comp_we g5929 (.nZ(w5767), .A(w6405), .Z(w5733) );
	vdp_sr_bit g5930 (.Q(w6405), .D(w5692), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5931 (.Q(w5768), .D(w5737), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5932 (.Q(w5813), .D(w5816), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5933 (.Q(w5816), .D(w5817), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5934 (.Q(w5817), .D(w5821), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5935 (.Q(w5821), .D(w5822), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5936 (.Q(w5822), .D(w5823), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5937 (.nQ(w5823), .D(w5826), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5938 (.nZ(w5776), .A(w5813) );
	vdp_sr_bit g5939 (.Q(w5827), .D(w5828), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5940 (.Q(w5828), .D(w5832), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5941 (.Q(w5832), .D(w5833), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5942 (.Q(w5833), .D(w5835), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5943 (.Q(w5835), .D(w5838), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5944 (.nQ(w5838), .D(w5837), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5945 (.nZ(w5778), .A(w5827) );
	vdp_sr_bit g5946 (.Q(w5839), .D(w6215), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5947 (.Q(w6215), .D(w5842), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5948 (.Q(w5842), .D(w5844), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5949 (.Q(w5844), .D(w5845), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5950 (.Q(w5845), .D(w5846), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5951 (.nQ(w5846), .D(w5850), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5952 (.nZ(w5802), .A(w5839) );
	vdp_sr_bit g5953 (.Q(w5851), .D(w5854), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5954 (.Q(w5854), .D(w5858), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5955 (.Q(w5858), .D(w5857), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5956 (.Q(w5857), .D(w5859), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5957 (.Q(w5859), .D(w5862), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5958 (.nQ(w5862), .D(w5863), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5959 (.nZ(w6407), .A(w5851) );
	vdp_sr_bit g5960 (.Q(w5866), .D(w5869), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5961 (.Q(w5869), .D(w5870), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5962 (.Q(w5870), .D(w5871), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5963 (.Q(w5871), .D(w5895), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5964 (.Q(w5895), .D(w5896), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5965 (.nQ(w5896), .D(w5876), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5966 (.nZ(w5788), .A(w5866) );
	vdp_sr_bit g5967 (.Q(w5897), .D(w5891), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5968 (.Q(w5891), .D(w5890), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5969 (.Q(w5890), .D(w5888), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5970 (.Q(w5888), .D(w5887), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5971 (.Q(w5887), .D(w5885), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5972 (.nQ(w5885), .D(w5875), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5973 (.nZ(w5791), .A(w5897) );
	vdp_sr_bit g5974 (.Q(w6408), .D(w5881), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5975 (.Q(w5881), .D(w5882), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5976 (.Q(w5882), .D(w5878), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5977 (.Q(w5878), .D(w5877), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5978 (.Q(w5877), .D(w5873), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5979 (.nQ(w5873), .D(w5874), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5980 (.nZ(w5796), .A(w6408) );
	vdp_and g5981 (.Z(w5775), .B(w5769), .A(w5679) );
	vdp_and g5982 (.Z(w5809), .B(w5444), .A(w5725) );
	vdp_and g5983 (.Z(w5810), .B(w5444), .A(w5724) );
	vdp_or g5984 (.Z(w6404), .B(w5809), .A(w5777) );
	vdp_and g5985 (.B(w5812), .A(M5), .Z(w5444) );
	vdp_or g5986 (.Z(w5783), .B(w5810), .A(w5777) );
	vdp_and g5987 (.Z(w5777), .B(w22), .A(w6417) );
	vdp_or g5988 (.Z(w5793), .B(w5777), .A(M5) );
	vdp_not g5989 (.nZ(w6417), .A(M5) );
	vdp_not g5990 (.nZ(w6406), .A(w5679) );
	vdp_nor g5991 (.Z(w5769), .B(w6405), .A(w5768) );
	vdp_sr_bit g5992 (.Q(w5825), .D(w5829), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5993 (.Q(w5829), .D(w5830), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5994 (.Q(w5830), .D(w5831), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5995 (.Q(w5831), .D(w5834), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5996 (.Q(w5834), .D(w6409), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5997 (.nQ(w6409), .D(w5903), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5998 (.nZ(w5722), .A(w5825) );
	vdp_sr_bit g5999 (.Q(w5814), .D(w5815), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6000 (.Q(w5815), .D(w5818), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6001 (.Q(w5818), .D(w5819), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6002 (.Q(w5819), .D(w5820), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6003 (.Q(w5820), .D(w5824), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6004 (.nQ(w5824), .D(w5902), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6005 (.nZ(w5723), .A(w5814) );
	vdp_sr_bit g6006 (.Q(w5804), .D(w5805), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6007 (.Q(w5805), .D(w5806), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6008 (.Q(w5806), .D(w5808), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6009 (.Q(w5808), .D(w5807), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6010 (.Q(w5807), .D(w5811), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6011 (.nQ(w5811), .D(w5901), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6012 (.nZ(w5812), .A(w5804) );
	vdp_sr_bit g6013 (.Q(w5836), .D(w5840), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6014 (.Q(w5840), .D(w5841), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6015 (.Q(w5841), .D(w5843), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6016 (.Q(w5843), .D(w5847), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6017 (.Q(w5847), .D(w5848), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6018 (.nQ(w5848), .D(w5908), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6019 (.nZ(w5721), .A(w5836) );
	vdp_sr_bit g6020 (.Q(w5849), .D(w5852), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6021 (.Q(w5852), .D(w5853), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6022 (.Q(w5853), .D(w5855), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6023 (.Q(w5855), .D(w5856), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6024 (.Q(w5856), .D(w5860), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6025 (.nQ(w5860), .D(w5904), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6026 (.nZ(w5725), .A(w5849) );
	vdp_sr_bit g6027 (.Q(w5861), .D(w5864), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6028 (.Q(w5864), .D(w5865), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6029 (.Q(w5865), .D(w5867), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6030 (.Q(w5867), .D(w5868), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6031 (.Q(w5868), .D(w5872), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6032 (.nQ(w5872), .D(w5905), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6033 (.nZ(w5724), .A(w5861) );
	vdp_sr_bit g6034 (.Q(w5893), .D(w5894), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6035 (.Q(w5894), .D(w5898), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6036 (.Q(w5898), .D(w5899), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6037 (.Q(w5899), .D(w5892), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6038 (.Q(w5892), .D(w5889), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6039 (.nQ(w5889), .D(w5906), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6040 (.nZ(w5770), .A(w5893) );
	vdp_sr_bit g6041 (.Q(w5884), .D(w5886), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6042 (.Q(w5886), .D(w5883), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6043 (.Q(w5883), .D(w5880), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6044 (.Q(w5880), .D(w5879), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6045 (.Q(w5879), .D(w5900), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6046 (.nQ(w5900), .D(w5907), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6047 (.nZ(w5771), .A(w5884) );
	vdp_slatch g6048 (.D(w5933), .nC(w5970), .C(w5911), .nQ(w5773) );
	vdp_slatch g6049 (.D(S[1]), .nC(w5971), .C(w5915), .Q(w5932) );
	vdp_slatch g6050 (.D(S[1]), .nC(w5972), .C(w5914), .Q(w5931) );
	vdp_aoi22 g6051 (.Z(w5930), .B2(w5976), .B1(w5932), .A1(w5931), .A2(w5912) );
	vdp_slatch g6052 (.D(S[0]), .nC(w5971), .C(w5915), .Q(w5935) );
	vdp_slatch g6053 (.D(S[0]), .nC(w5972), .C(w5914), .Q(w5934) );
	vdp_aoi22 g6054 (.Z(w5933), .B2(w5976), .B1(w5935), .A1(w5934), .A2(w5912) );
	vdp_slatch g6055 (.D(w5930), .nC(w5970), .C(w5911), .nQ(w5774) );
	vdp_slatch g6056 (.D(S[2]), .nC(w5971), .C(w5915), .Q(w5929) );
	vdp_slatch g6057 (.D(S[2]), .nC(w5972), .C(w5914), .Q(w5928) );
	vdp_aoi22 g6058 (.Z(w6012), .B2(w5976), .B1(w5929), .A1(w5928), .A2(w5912) );
	vdp_slatch g6059 (.D(w6012), .nC(w5970), .C(w5911), .nQ(w5799) );
	vdp_slatch g6060 (.D(S[3]), .nC(w5971), .C(w5915), .Q(w5927) );
	vdp_slatch g6061 (.D(S[3]), .nC(w5972), .C(w5914), .Q(w5926) );
	vdp_aoi22 g6062 (.Z(w5925), .B2(w5976), .B1(w5927), .A1(w5926), .A2(w5912) );
	vdp_slatch g6063 (.D(w5925), .nC(w5970), .C(w5911), .nQ(w5779) );
	vdp_slatch g6064 (.D(S[4]), .nC(w5971), .C(w5915), .Q(w5924) );
	vdp_slatch g6065 (.D(S[4]), .nC(w5972), .C(w5914), .Q(w5923) );
	vdp_aoi22 g6066 (.Z(w5922), .B2(w5976), .B1(w5924), .A1(w5923), .A2(w5912) );
	vdp_slatch g6067 (.D(w5922), .nC(w5970), .C(w5911), .nQ(w5782) );
	vdp_slatch g6068 (.D(S[5]), .nC(w5971), .C(w5915), .Q(w5921) );
	vdp_slatch g6069 (.D(S[5]), .nC(w5972), .C(w5914), .Q(w5920) );
	vdp_aoi22 g6070 (.Z(w5919), .B2(w5976), .B1(w5921), .A1(w5920), .A2(w5912) );
	vdp_slatch g6071 (.D(w5919), .nC(w5970), .C(w5911), .nQ(w5785) );
	vdp_slatch g6072 (.D(S[6]), .nC(w5971), .C(w5915), .Q(w5918) );
	vdp_slatch g6073 (.D(S[6]), .nC(w5972), .C(w5914), .Q(w5916) );
	vdp_aoi22 g6074 (.Z(w5917), .B2(w5976), .B1(w5918), .A1(w5916), .A2(w5912) );
	vdp_slatch g6075 (.D(w5917), .nC(w5970), .C(w5911), .nQ(w5789) );
	vdp_slatch g6076 (.D(S[7]), .nC(w5971), .C(w5915), .Q(w5913) );
	vdp_slatch g6077 (.D(S[7]), .nC(w5972), .C(w5914), .Q(w5909) );
	vdp_aoi22 g6078 (.Z(w5910), .B2(w5976), .B1(w5913), .A1(w5909), .A2(w5912) );
	vdp_slatch g6079 (.D(w5910), .nC(w5970), .C(w5911), .nQ(w5792) );
	vdp_comp_str g6080 (.nZ(w5970), .A(w5439), .Z(w5911) );
	vdp_comp_str g6081 (.nZ(w5971), .A(w4802), .Z(w5915) );
	vdp_comp_str g6082 (.nZ(w5972), .A(w4806), .Z(w5914) );
	vdp_comp_we g6083 (.nZ(w5976), .A(w5969), .Z(w5912) );
	vdp_sr_bit g6084 (.Q(w5967), .D(w5963), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6085 (.Z(w5963), .B(w5968), .A(w5936) );
	vdp_fa g6086 (.SUM(w5968), .CI(w5938), .A(w5967), .B(1'b0) );
	vdp_sr_bit g6087 (.Q(w6002), .D(w5958), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6088 (.Z(w5958), .B(w5964), .A(w5936) );
	vdp_fa g6089 (.SUM(w5964), .CO(w5938), .CI(w5939), .A(w6002), .B(1'b0) );
	vdp_sr_bit g6090 (.Q(w5959), .D(w5982), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6091 (.Z(w5982), .B(w5960), .A(w5936) );
	vdp_fa g6092 (.SUM(w5960), .CO(w5939), .CI(w5941), .A(w5959), .B(w5940) );
	vdp_sr_bit g6093 (.Q(w5955), .D(w5954), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6094 (.Z(w5954), .B(w5956), .A(w5936) );
	vdp_fa g6095 (.SUM(w5956), .CO(w5941), .CI(w5943), .A(w5955), .B(w5942) );
	vdp_sr_bit g6096 (.Q(w5946), .D(w6414), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6097 (.Q(w6414), .D(w21), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6098 (.nQ(w5944), .D(w5946), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g6099 (.nQ(w5936), .D(w5945), .nC(nHCLK1), .C(HCLK1) );
	vdp_and g6100 (.Z(w5940), .B(w5943), .A(w5951) );
	vdp_and g6101 (.Z(w5942), .B(w5943), .A(w5950) );
	vdp_and g6102 (.Z(w4446), .B(w6414), .A(w6026) );
	vdp_or g6103 (.Z(w5945), .B(w5948), .A(w6013) );
	vdp_not g6104 (.nZ(w5947), .A(M5) );
	vdp_not g6105 (.nZ(w5943), .A(w5944) );
	vdp_fa g6106 (.SUM(w5987), .CO(w5990), .CI(w5988), .A(w6040), .B(w5961) );
	vdp_aoi22 g6107 (.Z(w6051), .B2(w5973), .B1(w5989), .A1(w5987), .A2(w6036) );
	vdp_notif0 g6108 (.A(w6051), .nZ(VRAMA[9]), .nE(w6029) );
	vdp_fa g6109 (.SUM(w5978), .CO(w5988), .CI(w5984), .A(w6039), .B(w5965) );
	vdp_aoi22 g6110 (.Z(w5986), .B2(w5973), .B1(w5987), .A1(w5978), .A2(w6036) );
	vdp_notif0 g6111 (.A(w5986), .nZ(VRAMA[8]), .nE(w6029) );
	vdp_fa g6112 (.SUM(w5974), .CO(w5984), .CI(w5977), .A(w6038), .B(w5957) );
	vdp_aoi22 g6113 (.Z(w5985), .B2(w5973), .B1(w5978), .A1(w5974), .A2(w6036) );
	vdp_notif0 g6114 (.A(w5985), .nZ(VRAMA[7]), .nE(w6029) );
	vdp_fa g6115 (.SUM(w5980), .CO(w5977), .CI(1'b0), .A(w6037), .B(w5953) );
	vdp_aoi22 g6116 (.Z(w5975), .B2(w5973), .B1(w5974), .A1(w5980), .A2(w6036) );
	vdp_notif0 g6117 (.A(w5975), .nZ(VRAMA[6]), .nE(w6029) );
	vdp_not g6118 (.nZ(w6029), .A(w6043) );
	vdp_ha g6119 (.SUM(w5989), .B(w6041), .A(w5990), .CO(w5991) );
	vdp_aoi22 g6120 (.Z(w5993), .B2(w5973), .B1(w5992), .A1(w5989), .A2(w6036) );
	vdp_notif0 g6121 (.A(w5993), .nZ(VRAMA[10]), .nE(w6046) );
	vdp_ha g6122 (.SUM(w5992), .B(w6042), .A(w5991), .CO(w5994) );
	vdp_aoi22 g6123 (.Z(w5995), .B2(w5973), .B1(w6003), .A1(w5992), .A2(w6036) );
	vdp_notif0 g6124 (.A(w5995), .nZ(VRAMA[11]), .nE(w6046) );
	vdp_ha g6125 (.SUM(w6003), .B(w6045), .A(w5994), .CO(w5996) );
	vdp_aoi22 g6126 (.Z(w5998), .B2(w5973), .B1(w5997), .A1(w6003), .A2(w6036) );
	vdp_notif0 g6127 (.A(w5998), .nZ(VRAMA[12]), .nE(w6046) );
	vdp_ha g6128 (.SUM(w5997), .B(w6044), .A(w5996), .CO(w6000) );
	vdp_aoi22 g6129 (.Z(w6001), .B2(w5973), .B1(w5999), .A1(w5997), .A2(w6036) );
	vdp_notif0 g6130 (.A(w6001), .nZ(VRAMA[13]), .nE(w6046) );
	vdp_ha g6131 (.SUM(w5999), .B(w6048), .A(w6000), .CO(w6006) );
	vdp_aoi22 g6132 (.Z(w6004), .B2(w5973), .B1(w6005), .A1(w5999), .A2(w6036) );
	vdp_notif0 g6133 (.A(w6004), .nZ(VRAMA[14]), .nE(w6046) );
	vdp_ha g6134 (.SUM(w6005), .B(w6047), .A(w6006), .CO(w6007) );
	vdp_aoi22 g6135 (.Z(w6010), .B2(w5973), .B1(w6011), .A1(w6005), .A2(w6036) );
	vdp_notif0 g6136 (.A(w6010), .nZ(VRAMA[15]), .nE(w6046) );
	vdp_ha g6137 (.SUM(w6011), .B(w6050), .A(w6007) );
	vdp_aoi22 g6138 (.Z(w6009), .B2(w5973), .B1(w5068), .A1(w6011), .A2(w6036) );
	vdp_notif0 g6139 (.A(w6009), .nZ(VRAMA[16]), .nE(w6046) );
	vdp_not g6140 (.nZ(w6046), .A(w6043) );
	vdp_sr_bit g6141 (.Q(w6043), .D(w6194), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6142 (.nQ(w4370), .D(w6008), .nC(nHCLK2), .C(HCLK2) );
	vdp_and g6143 (.Z(w6194), .B(M5), .A(w21) );
	vdp_or9 g6144 (.Z(w6008), .B(w5907), .A(w5906), .C(w5826), .D(w5837), .F(w5863), .E(w5850), .G(w5876), .H(w5875), .I(w5874) );
	vdp_sr_bit g6145 (.Q(w4440), .D(w6294), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_sr_bit g6146 (.D(w6415), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_fa g6147 (.SUM(w5953), .CO(w6400), .CI(1'b0), .A(w6024), .B(w5954) );
	vdp_fa g6148 (.SUM(w5957), .CO(w6401), .CI(w6400), .A(w6025), .B(w5982) );
	vdp_fa g6149 (.SUM(w5965), .CO(w6402), .CI(w6401), .A(1'b0), .B(w5958) );
	vdp_fa g6150 (.SUM(w5961), .CI(w6402), .A(1'b0), .B(w5963) );
	vdp_notif0 g6151 (.A(1'b1), .nZ(VRAMA[0]), .nE(w6029) );
	vdp_notif0 g6152 (.A(1'b1), .nZ(VRAMA[1]), .nE(w6029) );
	vdp_not g6153 (.nZ(w5962), .A(w6030) );
	vdp_notif0 g6154 (.A(w5962), .nZ(VRAMA[2]), .nE(w6029) );
	vdp_not g6155 (.nZ(w5966), .A(w6032) );
	vdp_notif0 g6156 (.A(w5966), .nZ(VRAMA[3]), .nE(w6029) );
	vdp_not g6157 (.nZ(w5979), .A(w6031) );
	vdp_notif0 g6158 (.A(w5979), .nZ(VRAMA[4]), .nE(w6029) );
	vdp_notif0 g6159 (.A(w5981), .nZ(VRAMA[5]), .nE(w6029) );
	vdp_aoi22 g6160 (.Z(w5981), .B2(w5973), .B1(w5980), .A1(w6022), .A2(w6036) );
	vdp_comp_we g6161 (.nZ(w5973), .A(w1), .Z(w6036) );
	vdp_aon22 g6162 (.Z(w6024), .B2(w5949), .B1(w6022), .A1(w6020), .A2(w6023) );
	vdp_aon22 g6163 (.Z(w6025), .B2(w5949), .B1(w6020), .A1(w6019), .A2(w6023) );
	vdp_comp_we g6164 (.nZ(w5949), .A(w1), .Z(w6023) );
	vdp_or g6165 (.Z(w6415), .B(w6013), .A(w4446) );
	vdp_nor g6166 (.Z(w6294), .B(w5948), .A(w5947) );
	vdp_comp_str g6167 (.nZ(w6076), .A(w6033), .Z(w6049) );
	vdp_slatch g6168 (.D(w6079), .nC(w6076), .C(w6049), .Q(w5906) );
	vdp_aon22 g6169 (.Z(w6080), .B2(w6052), .B1(w5934), .A1(DB[0]), .A2(w6034) );
	vdp_slatch g6170 (.D(w6081), .nC(w6076), .C(w6049), .Q(w5907) );
	vdp_aon22 g6171 (.Z(w6082), .B2(w6052), .B1(w5931), .A1(DB[1]), .A2(w6034) );
	vdp_slatch g6172 (.D(w6083), .nC(w6076), .C(w6049), .Q(w5826) );
	vdp_aon22 g6173 (.Z(w6084), .B2(w6052), .B1(w5928), .A1(DB[2]), .A2(w6034) );
	vdp_slatch g6174 (.D(w6085), .nC(w6076), .C(w6049), .Q(w5837) );
	vdp_aon22 g6175 (.Z(w6086), .B2(w6052), .B1(w5926), .A1(DB[3]), .A2(w6034) );
	vdp_slatch g6176 (.D(w6087), .nC(w6076), .C(w6049), .Q(w5850) );
	vdp_aon22 g6177 (.Z(w6088), .B2(w6052), .B1(w5923), .A1(DB[4]), .A2(w6034) );
	vdp_slatch g6178 (.D(w6089), .nC(w6076), .C(w6049), .Q(w5863) );
	vdp_aon22 g6179 (.Z(w6090), .B2(w6052), .B1(w5920), .A1(DB[5]), .A2(w6034) );
	vdp_slatch g6180 (.D(w6091), .nC(w6076), .C(w6049), .Q(w5876) );
	vdp_aon22 g6181 (.Z(w6092), .B2(w6052), .B1(w5916), .A1(DB[6]), .A2(w6034) );
	vdp_slatch g6182 (.D(w6094), .nC(w6076), .C(w6049), .Q(w5875) );
	vdp_aon22 g6183 (.Z(w6137), .B2(w6052), .B1(w5909), .A1(DB[7]), .A2(w6034) );
	vdp_slatch g6184 (.D(w6093), .nC(w6076), .C(w6049), .Q(w5874) );
	vdp_aon22 g6185 (.Z(w6095), .B2(w6052), .B1(w4915), .A1(DB[8]), .A2(w6034) );
	vdp_slatch g6186 (.D(w6067), .nC(w6063), .C(w6035), .Q(w6039) );
	vdp_aon22 g6187 (.Z(w6102), .B2(w6052), .B1(w5929), .A1(DB[2]), .A2(w6034) );
	vdp_slatch g6188 (.D(w6066), .nC(w6063), .C(w6035), .Q(w6040) );
	vdp_aon22 g6189 (.Z(w6097), .B2(w6052), .B1(w5927), .A1(DB[3]), .A2(w6034) );
	vdp_slatch g6190 (.D(w6073), .nC(w6063), .C(w6035), .Q(w6041) );
	vdp_aon22 g6191 (.Z(w6098), .B2(w6052), .B1(w5924), .A1(DB[4]), .A2(w6034) );
	vdp_slatch g6192 (.D(w6072), .nC(w6063), .C(w6035), .Q(w6042) );
	vdp_aon22 g6193 (.Z(w6101), .B2(w6052), .B1(w5921), .A1(DB[5]), .A2(w6034) );
	vdp_slatch g6194 (.D(w6070), .nC(w6063), .C(w6035), .Q(w6045) );
	vdp_aon22 g6195 (.Z(w6103), .B2(w6052), .B1(w5918), .A1(DB[6]), .A2(w6034) );
	vdp_slatch g6196 (.D(w6071), .nC(w6063), .C(w6035), .Q(w6044) );
	vdp_aon22 g6197 (.Z(w6104), .B2(w6052), .B1(w5913), .A1(DB[7]), .A2(w6034) );
	vdp_slatch g6198 (.D(w6069), .nC(w6063), .C(w6035), .Q(w6048) );
	vdp_aon22 g6199 (.Z(w6105), .B2(w6052), .B1(w4856), .A1(DB[8]), .A2(w6034) );
	vdp_slatch g6200 (.D(w6061), .nC(w6063), .C(w6035), .Q(w6047) );
	vdp_aon22 g6201 (.Z(w6060), .B2(w6052), .B1(w4916), .A1(DB[9]), .A2(w6034) );
	vdp_slatch g6202 (.D(w6077), .nC(w6063), .C(w6035), .Q(w6050) );
	vdp_aon22 g6203 (.Z(w6078), .B2(w6052), .B1(w4923), .A1(DB[10]), .A2(w6034) );
	vdp_slatch g6204 (.D(w6064), .nC(w6063), .C(w6035), .Q(w6037) );
	vdp_aon22 g6205 (.Z(w6099), .B2(w6052), .B1(w5935), .A1(w6065), .A2(w6034) );
	vdp_slatch g6206 (.D(w6106), .nC(w6063), .C(w6035), .Q(w6038) );
	vdp_aon22 g6207 (.Z(w6100), .B2(w6052), .B1(w5932), .A1(DB[1]), .A2(w6034) );
	vdp_comp_str g6208 (.nZ(w6063), .A(w6033), .Z(w6035) );
	vdp_not g6209 (.nZ(w6033), .A(w6189) );
	vdp_oai21 g6210 (.Z(w6189), .B(HCLK1), .A1(w5948), .A2(w109) );
	vdp_sr_bit g6211 (.Q(w6190), .D(w6192), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6212 (.Q(w5439), .D(w6191), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6213 (.Q(w5969), .D(w6193), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6214 (.Q(w6096), .D(w5492), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g6215 (.Q(w6016), .D(w6021), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w6013), .CI(w21), .L(w6018), .nL(w6055), .CO(w6056) );
	vdp_cnt_bit_load g6216 (.Q(w6054), .D(w6017), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w6013), .CI(w6056), .L(w6018), .nL(w6055) );
	vdp_comp_we g6217 (.nZ(w6055), .A(w5948), .Z(w6018) );
	vdp_not g6218 (.nZ(w6021), .A(w6057) );
	vdp_not g6219 (.nZ(w6017), .A(w6053) );
	vdp_not g6220 (.nZ(w6014), .A(w108) );
	vdp_nand g6221 (.Z(w6107), .B(w108), .A(w4440) );
	vdp_nand g6222 (.Z(w6015), .B(w6014), .A(w4440) );
	vdp_not g6223 (.nZ(w6052), .A(w6015) );
	vdp_nor g6224 (.Z(w6026), .B(w6054), .A(w6016) );
	vdp_and g6225 (.Z(w5948), .B(w6026), .A(w21) );
	vdp_rs_ff g6226 (.Q(w6192), .R(w6027), .S(w6013) );
	vdp_and3 g6227 (.Z(w6191), .B(w5492), .A(w4447), .C(w6190) );
	vdp_cnt_bit g6228 (.Q(w6193), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w35), .CI(w6096) );
	vdp_not g6229 (.nZ(w6034), .A(w6107) );
	vdp_not g6230 (.nZ(w6059), .A(w4405) );
	vdp_not g6231 (.nZ(w6062), .A(w4406) );
	vdp_comp_str g6232 (.nZ(w6058), .A(w6033), .Z(w6109) );
	vdp_not g6233 (.nZ(w6117), .A(w109) );
	vdp_aon22 g6234 (.Z(w6119), .B2(w6052), .B1(w4974), .A1(DB[0]), .A2(w6034) );
	vdp_slatch g6235 (.D(w6108), .nC(w6058), .C(w6109), .Q(w5901) );
	vdp_bufif0 g6236 (.A(w6116), .Z(DB[0]), .nE(w6117) );
	vdp_aon222 g6237 (.Z(w6116), .B2(w4407), .B1(w5906), .A1(w5901), .A2(w6059), .C1(w6037), .C2(w6062) );
	vdp_aon22 g6238 (.Z(w6122), .B2(w6052), .B1(w5050), .A1(DB[1]), .A2(w6034) );
	vdp_slatch g6239 (.D(w6118), .nC(w6058), .C(w6109), .Q(w5902) );
	vdp_bufif0 g6240 (.A(w6120), .Z(DB[1]), .nE(w6117) );
	vdp_aon222 g6241 (.Z(w6120), .B2(w4407), .B1(w5907), .A1(w5902), .A2(w6059), .C1(w6038), .C2(w6062) );
	vdp_aon22 g6242 (.Z(w6124), .B2(w6052), .B1(w5069), .A1(DB[2]), .A2(w6034) );
	vdp_slatch g6243 (.D(w6121), .nC(w6058), .C(w6109), .Q(w5903) );
	vdp_bufif0 g6244 (.A(w6123), .Z(DB[2]), .nE(w6117) );
	vdp_aon222 g6245 (.Z(w6123), .B2(w4407), .B1(w5826), .A1(w5903), .A2(w6059), .C1(w6039), .C2(w6062) );
	vdp_aon22 g6246 (.Z(w6133), .B2(w6052), .B1(w5036), .A1(DB[3]), .A2(w6034) );
	vdp_slatch g6247 (.D(w6125), .nC(w6058), .C(w6109), .Q(w5908) );
	vdp_bufif0 g6248 (.A(w6132), .Z(DB[3]), .nE(w6117) );
	vdp_aon222 g6249 (.Z(w6132), .B2(w4407), .B1(w5837), .A1(w5908), .A2(w6059), .C1(w6040), .C2(w6062) );
	vdp_aon22 g6250 (.Z(w6130), .B2(w6052), .B1(w4386), .A1(DB[4]), .A2(w6034) );
	vdp_slatch g6251 (.D(w6057), .nC(w6058), .C(w6109), .Q(w5904) );
	vdp_bufif0 g6252 (.A(w6131), .Z(DB[4]), .nE(w6117) );
	vdp_aon222 g6253 (.Z(w6131), .B2(w4407), .B1(w5850), .A1(w5904), .A2(w6059), .C1(w6041), .C2(w6062) );
	vdp_aon22 g6254 (.Z(w6128), .B2(w6052), .B1(w4430), .A1(DB[5]), .A2(w6034) );
	vdp_slatch g6255 (.D(w6053), .nC(w6058), .C(w6109), .Q(w5905) );
	vdp_bufif0 g6256 (.A(w6129), .Z(DB[5]), .nE(w6117) );
	vdp_aon222 g6257 (.Z(w6129), .B2(w4407), .B1(w5863), .A1(w5905), .A2(w6059), .C1(w6042), .C2(w6062) );
	vdp_aon22 g6258 (.Z(w6126), .B2(w6052), .B1(w4387), .A1(DB[6]), .A2(w6034) );
	vdp_slatch g6259 (.D(w6127), .nC(w6058), .C(w6109), .Q(w5950) );
	vdp_bufif0 g6260 (.A(w6150), .Z(DB[6]), .nE(w6117) );
	vdp_aon222 g6261 (.Z(w6150), .B2(w4407), .B1(w5876), .A1(w5950), .A2(w6059), .C1(w6045), .C2(w6062) );
	vdp_aon22 g6262 (.Z(w6146), .B2(w6052), .B1(w4383), .A1(DB[7]), .A2(w6034) );
	vdp_slatch g6263 (.D(w6147), .nC(w6068), .C(w6148), .Q(w5951) );
	vdp_bufif0 g6264 (.A(w6149), .Z(DB[7]), .nE(w6117) );
	vdp_aon222 g6265 (.Z(w6149), .B2(w4407), .B1(w5875), .A1(w5951), .A2(w6059), .C1(w6044), .C2(w6062) );
	vdp_aon22 g6266 (.Z(w6144), .B2(w6052), .B1(w6110), .A1(DB[8]), .A2(w6034) );
	vdp_slatch g6267 (.D(w6145), .nC(w6068), .C(w6148), .Q(w6030) );
	vdp_bufif0 g6268 (.A(w6416), .Z(DB[8]), .nE(w6117) );
	vdp_aon222 g6269 (.Z(w6416), .B2(w4407), .B1(w5874), .A1(w6030), .A2(w6059), .C1(w6048), .C2(w6062) );
	vdp_aon22 g6270 (.Z(w6142), .B2(w6052), .B1(w6115), .A1(DB[9]), .A2(w6034) );
	vdp_slatch g6271 (.D(w6143), .nC(w6068), .C(w6148), .Q(w6032) );
	vdp_bufif0 g6272 (.A(w6151), .Z(DB[9]), .nE(w6117) );
	vdp_aon222 g6273 (.Z(w6151), .B2(w4407), .B1(1'b0), .A1(w6032), .A2(w6059), .C1(w6047), .C2(w6062) );
	vdp_aon22 g6274 (.Z(w6140), .B2(w6052), .B1(w6114), .A1(DB[10]), .A2(w6034) );
	vdp_slatch g6275 (.D(w6141), .nC(w6068), .C(w6148), .Q(w6031) );
	vdp_bufif0 g6276 (.A(w6152), .Z(DB[10]), .nE(w6117) );
	vdp_aon222 g6277 (.Z(w6152), .B2(w4407), .B1(1'b0), .A1(w6031), .A2(w6059), .C1(w6050), .C2(w6062) );
	vdp_aon22 g6278 (.Z(w6138), .B2(w6052), .B1(w6113), .A1(DB[11]), .A2(w6034) );
	vdp_slatch g6279 (.D(w6139), .nC(w6068), .C(w6148), .Q(w6022) );
	vdp_bufif0 g6280 (.A(w6022), .Z(DB[11]), .nE(w6117) );
	vdp_aon22 g6281 (.Z(w6136), .B2(w6052), .B1(w6112), .A1(DB[12]), .A2(w6034) );
	vdp_slatch g6282 (.D(w6153), .nC(w6068), .C(w6148), .Q(w6020) );
	vdp_bufif0 g6283 (.A(w6020), .Z(DB[12]), .nE(w6117) );
	vdp_aon22 g6284 (.Z(w6134), .B2(w6052), .B1(w6111), .A1(DB[13]), .A2(w6034) );
	vdp_slatch g6285 (.D(w6135), .nC(w6068), .C(w6148), .Q(w6019) );
	vdp_bufif0 g6286 (.A(w6019), .Z(DB[13]), .nE(w6117) );
	vdp_comp_str g6287 (.nZ(w6068), .A(w6033), .Z(w6148) );
	vdp_sr_bit g6288 (.Q(w4542), .D(w116), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6289 (.Q(w4546), .D(VRAMA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6290 (.Q(w6161), .D(w6154), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6291 (.Q(w4535), .D(VRAMA[3]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6292 (.Q(w4537), .D(VRAMA[4]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6293 (.Q(w4538), .D(VRAMA[5]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6294 (.Q(w4539), .D(VRAMA[6]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6295 (.Q(w4540), .D(VRAMA[7]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6296 (.Q(w4541), .D(VRAMA[8]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6297 (.Q(w4482), .D(w6158), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6298 (.Q(w4481), .D(w6159), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_and g6299 (.Z(w6158), .B(w119), .A(w6160) );
	vdp_and g6300 (.Z(w6159), .B(w118), .A(w6160) );
	vdp_sr_bit g6301 (.Q(w6174), .D(RD_DATA[0]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6302 (.Q(w6175), .D(RD_DATA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6303 (.Q(w6177), .D(w300), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6304 (.Q(w6176), .D(RD_DATA[2]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_V_PLA g6305 (.o0(w1807), .o1(w1808), .o2(w1809), .o3(w1810), .o4(w1811), .o5(w1812), .o6(w1813), .o7(w1814), .o8(w1815), .o9(w1816), .o10(w1817), .o11(w6614), .o12(w6615), .o13(w6613), .o14(w1818), .o15(w6534), .o16(w6535), .o17(w6536), .o18(w1819), .o19(w1820), .o20(w1821), .o21(w1822), .o22(w6537), .o23(w1823), .o24(w1902), .o25(w1824), .o26(w1825), .o27(w1903), .o28(w1918), .o29(w1917), .o30(w1938), .o31(w1841), .o32(w1806), .o33(w1805), .o34(w1842), .o35(w1826), .o36(w1843), .o37(w1844), .o38(w1804), .o39(w1803), .o40(w1847), .o41(w1845), .o42(w1846), .o43(w1802), .o44(w1801), .o45(w1800), .o46(w1799), .o47(w6423), .Vcnt0(w1637), .Vcnt1(w1775), .Vcnt2(w1857), .Vcnt3(w1760), .Vcnt4(w1856), .Vcnt5(w1855), .Vcnt6(w1680), .Vcnt7(w1854), .Vcnt8(w1777), .ODD_EVEN(ODD_EVEN), .LS0(w1016), .PAL(PAL), .nPAL(w1768), .i2(w1767), .i3(w1756), .M5(M5) );
	vdp_not g6306 (.A(w757), .nZ(w6421) );
	vdp_not g6307 (.A(w924), .nZ(w6422) );
	vdp_not g6308 (.nZ(w2367), .A(w6421) );
	vdp_not g6309 (.nZ(w2368), .A(w6422) );
	vdp_cram g6310 (.q8(w2654), .D8(w2659), .q7(w2756), .D7(w2655), .q6(w2653), .D6(w2656), .q5(w2658), .D5(w2657), .q4(w2652), .D4(w2660), .q3(w2661), .D3(w2878), .q2(w2651), .D2(w2662), .q1(w2650), .D1(w2663), .q0(w2648), .D0(w2664), .A0(w2683), .A1(w2687), .CLK(HCLK1), .A2(w2693), .A3(w2703), .A4(w2724), .A5(w2723), .WE(w2730), .RD(w2729) );
	vdp_linebuf_ram g6311 (.q0(w5172), .D0(w5522), .q1(w5152), .D1(w5521), .q2(w5114), .D2(w5520), .q3(w5191), .D3(w5535), .q4(w5543), .D4(w5536), .q5(w5550), .D5(w5537), .q6(w5509), .D6(w5538), .q7(w5171), .D7(w5519), .q8(w5155), .D8(w5518), .q9(w5135), .D9(w5517), .q10(w5508), .D10(w5499), .q11(w5510), .D11(w5498), .q12(w5511), .D12(w5531), .q13(w5514), .D13(w5532), .q14(w5170), .D14(w5522), .q15(w5153), .D15(w5521), .q16(w5137), .D16(w5520), .q17(w5183), .D17(w5523), .q18(w5512), .D18(w5530), .q19(w5513), .D19(w5524), .q20(w5526), .D20(w5525), .q21(w5169), .D21(w5519), .q22(w5159), .D22(w5518), .q23(w5132), .D23(w5517), .q24(w5184), .D24(w5505), .q25(w5502), .D25(w5503), .q26(w5507), .D26(w5516), .q27(w5529), .D27(w5515), .CLK(w4368), .A5(w4362), .A4(w4363), .A3(w4364), .A2(w4365), .A1(w4366), .A0(w4367), .Ai(w5528), .Bi(w5497), .Ci(w5496), .Di(w5495) );
	vdp_linebuf_ram g6312 (.q0(w5178), .D0(w5522), .q1(w5149), .D1(w5521), .q2(w5140), .D2(w5520), .q3(w5121), .D3(w5167), .q4(w5120), .D4(w5165), .q5(w5119), .D5(w5166), .q6(w5504), .D6(w6156), .q7(w5173), .D7(w5519), .q8(w5151), .D8(w5518), .q9(w5138), .D9(w5517), .q10(w5188), .D10(w5161), .q11(w5117), .D11(w5162), .q12(w5118), .D12(w5163), .q13(w5501), .D13(w5156), .q14(w5174), .D14(w5522), .q15(w5150), .D15(w5521), .q16(w5141), .D16(w5520), .q17(w5195), .D17(w5130), .q18(w5115), .D18(w5113), .q19(w5116), .D19(w5128), .q20(w5500), .D20(w5129), .q21(w5123), .D21(w5519), .q22(w5122), .D22(w5518), .q23(w5136), .D23(w5517), .q24(w5189), .D24(w6157), .q25(w5533), .D25(w5124), .q26(w5534), .D26(w5125), .q27(w5506), .D27(w5126), .A0(w4367), .CLK(w4368), .A5(w4362), .A3(w4364), .A4(w4363), .A2(w4365), .A1(w4366), .Ai(w5237), .Bi(w5221), .Ci(w5233), .Di(w5223) );
	vdp_att_cashe_ram2 g6313 (.q0(w4559), .D0(FIFOo[0]), .q1(w4558), .D1(FIFOo[1]), .q2(w4557), .D2(FIFOo[2]), .q3(w4556), .D3(FIFOo[3]), .q4(w4532), .D4(FIFOo[4]), .q5(w4531), .D5(FIFOo[5]), .q6(w4526), .D6(FIFOo[6]), .q7(w4702), .D7(w6174), .q8(w4741), .D8(w6175), .q9(w4725), .D9(w6176), .q10(w4722), .D10(w6177), .CLK(HCLK1), .A6(w6181), .A5(w6182), .A1(w6187), .A0(w6186), .A4(w6183), .A3(w6184), .A2(w6185), .Ai(w6178), .Bi(w4544) );
	vdp_att_cashe_ram1 g6314 (.q0(w4591), .D0(FIFOo[0]), .q1(w4594), .D1(FIFOo[1]), .q2(w4587), .D2(FIFOo[2]), .q3(w4588), .D3(FIFOo[3]), .q4(w4570), .D4(FIFOo[4]), .q5(w4562), .D5(FIFOo[5]), .q6(w4563), .D6(FIFOo[6]), .q7(w4561), .D7(FIFOo[7]), .q8(w4560), .D8(w6174), .q9(w4555), .D9(w6175), .CLK(HCLK1), .A0(w6186), .A1(w6187), .A2(w6185), .A3(w6184), .A4(w6183), .A5(w6182), .A6(w6181), .Ai(w6180), .Bi(w6179) );
	vdp_att_temp_ram g6315 (.A4(w4464), .A0(w4468), .A1(w4467), .A2(w4466), .A3(w4465), .q0(w6064), .D0(w6099), .q1(w6106), .D1(w6100), .q2(w6067), .D2(w6102), .q3(w6066), .D3(w6097), .q4(w6073), .D4(w6098), .q5(w6072), .D5(w6101), .q6(w6070), .D6(w6103), .q7(w6071), .D7(w6104), .q8(w6069), .D8(w6105), .q9(w6061), .D9(w6060), .q10(w6077), .D10(w6078), .q11(w6079), .D11(w6080), .q12(w6081), .D12(w6082), .q13(w6083), .D13(w6084), .q14(w6085), .D14(w6086), .q15(w6087), .D15(w6088), .q16(w6089), .D16(w6090), .q17(w6091), .D17(w6092), .q18(w6094), .D18(w6137), .q19(w6093), .D19(w6095), .q20(w6108), .D20(w6119), .q21(w6118), .D21(w6122), .q22(w6121), .D22(w6124), .q23(w6125), .D23(w6133), .q24(w6057), .D24(w6130), .q25(w6053), .D25(w6128), .q26(w6127), .D26(w6126), .q26(w6147), .D26(w6146), .q27(w6145), .D27(w6144), .q28(w6143), .D28(w6142), .q29(w6141), .D29(w6140), .q30(w6139), .D30(w6138), .q31(w6153), .D[31](w6136), .q32(w6135), .D32(w6134), .CLK(HCLK1), .Ai(w4439), .Bi(w4431), .Ci(w4435) );
	vdp_vsram g6316 (.CLK(HCLK1), .D10(w3864), .q10(w3827), .D9(w3868), .q9(w3820), .D8(w3866), .q8(w3842), .D7(w3865), .q7(w3812), .D6(w3854), .q6(w3808), .D5(w3852), .q5(w3800), .D4(w3859), .q4(w3796), .D3(w3861), .q3(w3793), .D2(w3863), .q2(w3847), .D1(w3826), .q1(w3788), .D0(w3840), .q0(w3783), .A1(w3607), .A2(w3579), .A3(w3578), .A4(w3577), .A5(w3576), .A0(w3608), .Ai(w3575), .Bi(w3574) );
	vdp_not g6317 (.nZ(w1750), .A(w6423) );
	vdp_not g6318 (.nZ(PAL), .A(w6424) );
	vdp_H_PLA g6319 (.HPLA0(HPLA0), .HPLA1(HPLA1), .HPLA2(HPLA2), .HPLA3(HPLA3), .HPLA4(HPLA4), .HPLA5(HPLA5), .HPLA7(HPLA7), .HPLA8(HPLA8), .HPLA9(HPLA9), .HPLA6(HPLA6), .HPLA10(HPLA10), .HPLA11(HPLA11), .HPLA16(HPLA16), .HPLA15(HPLA15), .HPLA14(HPLA14), .HPLA13(HPLA13), .HPLA12(HPLA12), .i0(w56), .HPLA17(HPLA17), .HPLA18(HPLA18), .HPLA19(HPLA19), .HPLA20(HPLA20), .HPLA21(HPLA21), .HPLA22(HPLA22), .Hcnt0(w1860), .Hcnt1(w1625), .Hcnt2(w1626), .Hcnt3(w1624), .Hcnt4(w1668), .Hcnt5(w1700), .Hcnt6(w1833), .Hcnt7(w1677), .Hcnt8(w1873), .H40(H40), .M5(M5), .B(w1862), .C(w1776), .A(w1673), .HPLA23(HPLA23), .HPLA24(HPLA24), .HPLA25(HPLA25), .HPLA26(HPLA26), .HPLA27(HPLA27), .HPLA28(HPLA28), .HPLA29(HPLA29), .HPLA30(HPLA30), .HPLA31(HPLA31), .HPLA32(HPLA32), .HPLA33(HPLA33), .i3(w1837), .HPLA35(HPLA35), .HPLA36(HPLA36), .HPLA34(HPLA34) );
	vdp_slatch g5073 (.D(S[4]), .nC(w4861), .C(w4862), .Q(w5049) );
endmodule // VDP

// Module Definitions [It is possible to wrap here on your primitives]

module vdp_slatch (  nQ, D, C, nC);

	output wire nQ;
	input wire D;
	input wire C;
	input wire nC;

endmodule // vdp_slatch

module vdp_sr_bit (  D, C2, C1, Q, nC2, nC1);

	input wire D;
	input wire C2;
	input wire C1;
	output wire Q;
	input wire nC2;
	input wire nC1;

endmodule // vdp_sr_bit

module vdp_notif0 (  A, nZ, nE);

	input wire A;
	output wire nZ;
	input wire nE;

endmodule // vdp_notif0

module vdp_aon22 (  Z, A1, A2, B1, B2);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire B1;
	input wire B2;

endmodule // vdp_aon22

module vdp_not (  A, nZ);

	input wire A;
	output wire nZ;

endmodule // vdp_not

module vdp_comp_str (  A, Z, nZ);

	input wire A;
	output wire Z;
	output wire nZ;

endmodule // vdp_comp_str

module vdp_comp_we (  A, Z, nZ);

	input wire A;
	output wire Z;
	output wire nZ;

endmodule // vdp_comp_we

module vdp_and (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_and

module vdp_nand (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_nand

module vdp_and3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_and3

module vdp_fa (  SUM, A, B, CO, CI);

	output wire SUM;
	input wire A;
	input wire B;
	output wire CO;
	input wire CI;

endmodule // vdp_fa

module vdp_comp_dff (  D, C2, C1, Q, nC2, nC1);

	input wire D;
	input wire C2;
	input wire C1;
	output wire Q;
	input wire nC2;
	input wire nC1;

endmodule // vdp_comp_dff

module vdp_or (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_or

module vdp_xor (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_xor

module vdp_aoi21 (  Z, B, A1, A2);

	output wire Z;
	input wire B;
	input wire A1;
	input wire A2;

endmodule // vdp_aoi21

module vdp_nor (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_nor

module vdp_and5 (  Z, A, B, C, D, E);

	output wire Z;
	input wire A;
	input wire B;
	input wire C;
	input wire D;
	input wire E;

endmodule // vdp_and5

module vdp_aon2222 (  C2, B2, A2, C1, B1, A1, Z, D2, D1);

	input wire C2;
	input wire B2;
	input wire A2;
	input wire C1;
	input wire B1;
	input wire A1;
	output wire Z;
	input wire D2;
	input wire D1;

endmodule // vdp_aon2222

module vdp_cnt_bit (  R, Q, C1, C2, nC1, nC2, CI);

	input wire R;
	output wire Q;
	input wire C1;
	input wire C2;
	input wire nC1;
	input wire nC2;
	input wire CI;

endmodule // vdp_cnt_bit

module vdp_oai21 (  A1, Z, A2, B);

	input wire A1;
	output wire Z;
	input wire A2;
	input wire B;

endmodule // vdp_oai21

module vdp_comb1 (  Z, C1, B, C2, A);

	output wire Z;
	input wire C1;
	input wire B;
	input wire C2;
	input wire A;

endmodule // vdp_comb1

module vdp_rs_ff (  Q, R, S);

	output wire Q;
	input wire R;
	input wire S;

endmodule // vdp_rs_ff

module vdp_and4 (  A, Z, B, C, D);

	input wire A;
	output wire Z;
	input wire B;
	input wire C;
	input wire D;

endmodule // vdp_and4

module vdp_or3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_or3

module vdp_bufif0 (  A, Z, nE);

	input wire A;
	output wire Z;
	input wire nE;

endmodule // vdp_bufif0

module vdp_aoi221 (  Z, A2, B1, B2, A1, C);

	output wire Z;
	input wire A2;
	input wire B1;
	input wire B2;
	input wire A1;
	input wire C;

endmodule // vdp_aoi221

module vdp_aon33 (  Z, A2, B1, B2, A1, A3, B3);

	output wire Z;
	input wire A2;
	input wire B1;
	input wire B2;
	input wire A1;
	input wire A3;
	input wire B3;

endmodule // vdp_aon33

module vdp_dlatch_inv (  D, C, Q, nC);

	input wire D;
	input wire C;
	output wire Q;
	input wire nC;

endmodule // vdp_dlatch_inv

module vdp_cnt_bit_load (  D, nL, L, R, Q, C1, C2, nC1, nC2, CI, CO);

	input wire D;
	input wire nL;
	input wire L;
	input wire R;
	output wire Q;
	input wire C1;
	input wire C2;
	input wire nC1;
	input wire nC2;
	input wire CI;
	output wire CO;

endmodule // vdp_cnt_bit_load

module vdp_nand3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_nand3

module vdp_nor3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_nor3

module vdp_dff (  Q, R, C, D);

	output wire Q;
	input wire R;
	input wire C;
	input wire D;

endmodule // vdp_dff

module vdp_ha (  SUM, A, B, CO);

	output wire SUM;
	input wire A;
	input wire B;
	output wire CO;

endmodule // vdp_ha

module vdp_slatch_r (  Q, D, R, C, nC);

	output wire Q;
	input wire D;
	input wire R;
	input wire C;
	input wire nC;

endmodule // vdp_slatch_r

module vdp_or5 (  C, A, B, Z, D, E);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;
	input wire E;

endmodule // vdp_or5

module vdp_2a3oi (  A1, B, Z, A2, C);

	input wire A1;
	input wire B;
	output wire Z;
	input wire A2;
	input wire C;

endmodule // vdp_2a3oi

module vdp_nor5 (  C, A, B, Z, D, E);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;
	input wire E;

endmodule // vdp_nor5

module vdp_or4 (  C, A, B, Z, D);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;

endmodule // vdp_or4

module vdp_aoi22 (  Z, A1, A2, B1, B2);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire B1;
	input wire B2;

endmodule // vdp_aoi22

module vdp_aon222 (  C2, B2, A2, C1, B1, A1, Z);

	input wire C2;
	input wire B2;
	input wire A2;
	input wire C1;
	input wire B1;
	input wire A1;
	output wire Z;

endmodule // vdp_aon222

module vdp_dlatch (  D, C, Q, nC);

	input wire D;
	input wire C;
	output wire Q;
	input wire nC;

endmodule // vdp_dlatch

module vdp_nor4 (  C, A, B, Z, D);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;

endmodule // vdp_nor4

module vdp_and6 (  C, A, B, Z, D, E, F);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;
	input wire E;
	input wire F;

endmodule // vdp_and6

module vdp_n_fet (  Z, A);

	output wire Z;
	input wire A;

endmodule // vdp_n_fet

module vdp_tff (  C2, C1, nC2, nC1, CI, R, A, Q);

	input wire C2;
	input wire C1;
	input wire nC2;
	input wire nC1;
	input wire CI;
	input wire R;
	input wire A;
	output wire Q;

endmodule // vdp_tff

module vdp_sdelay8 (  Q, D, nC1, C1, nC2, C2, nC3, C3, nC4, C4, nC5, C5, nC6, C6, nC7, C7, nC8, C8, nC9, C9, nC10, C10, nC11, C11, nC12, C12, nC13, C13, nC14, C14, nC15, C15, nC16, C16);

	output wire Q;
	input wire D;
	input wire nC1;
	input wire C1;
	input wire nC2;
	input wire C2;
	input wire nC3;
	input wire C3;
	input wire nC4;
	input wire C4;
	input wire nC5;
	input wire C5;
	input wire nC6;
	input wire C6;
	input wire nC7;
	input wire C7;
	input wire nC8;
	input wire C8;
	input wire nC9;
	input wire C9;
	input wire nC10;
	input wire C10;
	input wire nC11;
	input wire C11;
	input wire nC12;
	input wire C12;
	input wire nC13;
	input wire C13;
	input wire nC14;
	input wire C14;
	input wire nC15;
	input wire C15;
	input wire nC16;
	input wire C16;

endmodule // vdp_sdelay8

module vdp_sdelay7 (  Q, D, C1, nC1, C2, nC2, nC3, C4, nC4, C5, nC5, C6, nC6, C7, nC7, C8, nC8, C9, nC9, C10, nC10, C11, nC11, C12, nC12, C13, nC13, C14, nC14, C3);

	output wire Q;
	input wire D;
	input wire C1;
	input wire nC1;
	input wire C2;
	input wire nC2;
	input wire nC3;
	input wire C4;
	input wire nC4;
	input wire C5;
	input wire nC5;
	input wire C6;
	input wire nC6;
	input wire C7;
	input wire nC7;
	input wire C8;
	input wire nC8;
	input wire C9;
	input wire nC9;
	input wire C10;
	input wire nC10;
	input wire C11;
	input wire nC11;
	input wire C12;
	input wire nC12;
	input wire C13;
	input wire nC13;
	input wire C14;
	input wire nC14;
	input wire C3;

endmodule // vdp_sdelay7

module vdp_or8 (  Z, A, B, C, D, E, F, G, H);

	output wire Z;
	input wire A;
	input wire B;
	input wire C;
	input wire D;
	input wire E;
	input wire F;
	input wire G;
	input wire H;

endmodule // vdp_or8

module vdp_or7 (  Z, A, B, C, D, E, F, G);

	output wire Z;
	input wire A;
	input wire B;
	input wire C;
	input wire D;
	input wire E;
	input wire F;
	input wire G;

endmodule // vdp_or7

module vdp_clkgen (  PH, CLK1, nCLK1, CLK2, nCLK2);

	input wire PH;
	output wire CLK1;
	output wire nCLK1;
	output wire CLK2;
	output wire nCLK2;

endmodule // vdp_clkgen

module vdp_cgi2a (  Z, A, C, B);

	output wire Z;
	input wire A;
	input wire C;
	input wire B;

endmodule // vdp_cgi2a

module vdp_nand4 (  Z, A, B, D, C);

	output wire Z;
	input wire A;
	input wire B;
	input wire D;
	input wire C;

endmodule // vdp_nand4

module vdp_lfsr_bit (  Q, A, C2, C1, nC2, nC1, C, B);

	output wire Q;
	input wire A;
	input wire C2;
	input wire C1;
	input wire nC2;
	input wire nC1;
	input wire C;
	input wire B;

endmodule // vdp_lfsr_bit

module vdp_aoi222 (  Z, A1, B1, B2, A2, C1, C2);

	output wire Z;
	input wire A1;
	input wire B1;
	input wire B2;
	input wire A2;
	input wire C1;
	input wire C2;

endmodule // vdp_aoi222

module vdp_aon333 (  Z, A1, A2, A3, B1, B2, B3, C1, C2, C3);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire A3;
	input wire B1;
	input wire B2;
	input wire B3;
	input wire C1;
	input wire C2;
	input wire C3;

endmodule // vdp_aon333

module vdp_aoi33 (  Z, A1, A2, A3, B1, B2, B3);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire A3;
	input wire B1;
	input wire B2;
	input wire B3;

endmodule // vdp_aoi33

module vdp_comp_strong (  nZ, Z, A);

	output wire nZ;
	output wire Z;
	input wire A;

endmodule // vdp_comp_strong

module vdp_neg_dff (  Q, C, D, R);

	output wire Q;
	input wire C;
	input wire D;
	input wire R;

endmodule // vdp_neg_dff

module vdp_aon2x8 (  Z, A1, B1, C1, D2, A2, B2, C2, D1, E2, F1, E1, F2, G1, H2, G2, H1);

	output wire Z;
	input wire A1;
	input wire B1;
	input wire C1;
	input wire D2;
	input wire A2;
	input wire B2;
	input wire C2;
	input wire D1;
	input wire E2;
	input wire F1;
	input wire E1;
	input wire F2;
	input wire G1;
	input wire H2;
	input wire G2;
	input wire H1;

endmodule // vdp_aon2x8

module vdp_xnor (  Z, A, B);

	output wire Z;
	input wire A;
	input wire B;

endmodule // vdp_xnor

module vdp_oai211 (  Z, A1, A2, B, C);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire B;
	input wire C;

endmodule // vdp_oai211

module vdp_aoi31 (  Z, B3, B2, B1, A);

	output wire Z;
	input wire B3;
	input wire B2;
	input wire B1;
	input wire A;

endmodule // vdp_aoi31

module vdp_cnt_bit_rev (  nC2, nC1, C2, C1, Q, CI, B, A);

	input wire nC2;
	input wire nC1;
	input wire C2;
	input wire C1;
	output wire Q;
	input wire CI;
	input wire B;
	input wire A;

endmodule // vdp_cnt_bit_rev

module vdp_2x_sr_bit (  Q, D, nC2, nC1, C2, C1, nC4, nC3, C4, C3);

	output wire Q;
	input wire D;
	input wire nC2;
	input wire nC1;
	input wire C2;
	input wire C1;
	input wire nC4;
	input wire nC3;
	input wire C4;
	input wire C3;

endmodule // vdp_2x_sr_bit

module vdp_and9 (  Z, B, A, C, D, F, E, G, H, I);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;
	input wire I;

endmodule // vdp_and9

module vdp_nor12 (  Z, B, A, C, D, F, E, G, H, J, I, K, L);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;
	input wire J;
	input wire I;
	input wire K;
	input wire L;

endmodule // vdp_nor12

module vdp_nor8 (  Z, B, A, C, D, F, E, G, H);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;

endmodule // vdp_nor8

module vdp_aon21_sr (  Q, A1, A2, B, nC2, nC1, C2, C1);

	output wire Q;
	input wire A1;
	input wire A2;
	input wire B;
	input wire nC2;
	input wire nC1;
	input wire C2;
	input wire C1;

endmodule // vdp_aon21_sr

module vdp_or9 (  Z, B, A, C, D, F, E, G, H, I);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;
	input wire I;

endmodule // vdp_or9

module vdp_V_PLA (  o0, o1, o2, o3, o4, o5, o6, o7, o8, o9, o10, o11, o12, o13, o14, o15, o16, o17, o18, o19, o20, o21, o22, o23, o24, o25, o26, o27, o28, o29, o30, o31, o32, o33, o34, o35, o36, o37, o38, o39, o40, o41, o42, o43, o44, o45, o46, o47, Vcnt0, Vcnt1, Vcnt2, Vcnt3, Vcnt4, Vcnt5, Vcnt6, Vcnt7, Vcnt8, ODD_EVEN, LS0, PAL, nPAL, i2, i3, M5);

	output wire o0;
	output wire o1;
	output wire o2;
	output wire o3;
	output wire o4;
	output wire o5;
	output wire o6;
	output wire o7;
	output wire o8;
	output wire o9;
	output wire o10;
	output wire o11;
	output wire o12;
	output wire o13;
	output wire o14;
	output wire o15;
	output wire o16;
	output wire o17;
	output wire o18;
	output wire o19;
	output wire o20;
	output wire o21;
	output wire o22;
	output wire o23;
	output wire o24;
	output wire o25;
	output wire o26;
	output wire o27;
	output wire o28;
	output wire o29;
	output wire o30;
	output wire o31;
	output wire o32;
	output wire o33;
	output wire o34;
	output wire o35;
	output wire o36;
	output wire o37;
	output wire o38;
	output wire o39;
	output wire o40;
	output wire o41;
	output wire o42;
	output wire o43;
	output wire o44;
	output wire o45;
	output wire o46;
	output wire o47;
	input wire Vcnt0;
	input wire Vcnt1;
	input wire Vcnt2;
	input wire Vcnt3;
	input wire Vcnt4;
	input wire Vcnt5;
	input wire Vcnt6;
	input wire Vcnt7;
	input wire Vcnt8;
	input wire ODD_EVEN;
	input wire LS0;
	input wire PAL;
	input wire nPAL;
	input wire i2;
	input wire i3;
	input wire M5;

endmodule // vdp_V_PLA

module vdp_cram (  q8, D8, q7, D7, q6, D6, q5, D5, q4, D4, q3, D3, q2, D2, q1, D1, q0, D0, A0, A1, CLK, A2, A3, A4, A5, WE, RD);

	output wire q8;
	input wire D8;
	output wire q7;
	input wire D7;
	output wire q6;
	input wire D6;
	output wire q5;
	input wire D5;
	output wire q4;
	input wire D4;
	output wire q3;
	input wire D3;
	output wire q2;
	input wire D2;
	output wire q1;
	input wire D1;
	output wire q0;
	input wire D0;
	input wire A0;
	input wire A1;
	input wire CLK;
	input wire A2;
	input wire A3;
	input wire A4;
	input wire A5;
	input wire WE;
	input wire RD;

endmodule // vdp_cram

module vdp_linebuf_ram (  q0, D0, q1, D1, q2, D2, q3, D3, q4, D4, q5, D5, q6, D6, q7, D7, q8, D8, q9, D9, q10, D10, q11, D11, q12, D12, q13, D13, q14, D14, q15, D15, q16, D16, q17, D17, q18, D18, q19, D19, q20, D20, q21, D21, q22, D22, q23, D23, q24, D24, q25, D25, q26, D26, q27, D27, CLK, A5, A4, A3, A2, A1, A0, Ai, Bi, Ci, Di);

	output wire q0;
	input wire D0;
	output wire q1;
	input wire D1;
	output wire q2;
	input wire D2;
	output wire q3;
	input wire D3;
	output wire q4;
	input wire D4;
	output wire q5;
	input wire D5;
	output wire q6;
	input wire D6;
	output wire q7;
	input wire D7;
	output wire q8;
	input wire D8;
	output wire q9;
	input wire D9;
	output wire q10;
	input wire D10;
	output wire q11;
	input wire D11;
	output wire q12;
	input wire D12;
	output wire q13;
	input wire D13;
	output wire q14;
	input wire D14;
	output wire q15;
	input wire D15;
	output wire q16;
	input wire D16;
	output wire q17;
	input wire D17;
	output wire q18;
	input wire D18;
	output wire q19;
	input wire D19;
	output wire q20;
	input wire D20;
	output wire q21;
	input wire D21;
	output wire q22;
	input wire D22;
	output wire q23;
	input wire D23;
	output wire q24;
	input wire D24;
	output wire q25;
	input wire D25;
	output wire q26;
	input wire D26;
	output wire q27;
	input wire D27;
	input wire CLK;
	input wire A5;
	input wire A4;
	input wire A3;
	input wire A2;
	input wire A1;
	input wire A0;
	input wire Ai;
	input wire Bi;
	input wire Ci;
	input wire Di;

endmodule // vdp_linebuf_ram

module vdp_att_cashe_ram2 (  q0, D0, q1, D1, q2, D2, q3, D3, q4, D4, q5, D5, q6, D6, q7, D7, q8, D8, q9, D9, q10, D10, CLK, A6, A5, A1, A0, A4, A3, A2, Ai, Bi);

	output wire q0;
	input wire D0;
	output wire q1;
	input wire D1;
	output wire q2;
	input wire D2;
	output wire q3;
	input wire D3;
	output wire q4;
	input wire D4;
	output wire q5;
	input wire D5;
	output wire q6;
	input wire D6;
	output wire q7;
	input wire D7;
	output wire q8;
	input wire D8;
	output wire q9;
	input wire D9;
	output wire q10;
	input wire D10;
	input wire CLK;
	input wire A6;
	input wire A5;
	input wire A1;
	input wire A0;
	input wire A4;
	input wire A3;
	input wire A2;
	input wire Ai;
	input wire Bi;

endmodule // vdp_att_cashe_ram2

module vdp_att_cashe_ram1 (  q0, D0, q1, D1, q2, D2, q3, D3, q4, D4, q5, D5, q6, D6, q7, D7, q8, D8, q9, D9, CLK, A0, A1, A2, A3, A4, A5, A6, Ai, Bi);

	output wire q0;
	input wire D0;
	output wire q1;
	input wire D1;
	output wire q2;
	input wire D2;
	output wire q3;
	input wire D3;
	output wire q4;
	input wire D4;
	output wire q5;
	input wire D5;
	output wire q6;
	input wire D6;
	output wire q7;
	input wire D7;
	output wire q8;
	input wire D8;
	output wire q9;
	input wire D9;
	input wire CLK;
	input wire A0;
	input wire A1;
	input wire A2;
	input wire A3;
	input wire A4;
	input wire A5;
	input wire A6;
	input wire Ai;
	input wire Bi;

endmodule // vdp_att_cashe_ram1

module vdp_att_temp_ram (  A4, A0, A1, A2, A3, q0, D0, q1, D1, q2, D2, q3, D3, q4, D4, q5, D5, q6, D6, q7, D7, q8, D8, q9, D9, q10, D10, q11, D11, q12, D12, q13, D13, q14, D14, q15, D15, q16, D16, q17, D17, q18, D18, q19, D19, q20, D20, q21, D21, q22, D22, q23, D23, q24, D24, q25, D25, q26, D26, q26, D26, q27, D27, q28, D28, q29, D29, q30, D30, q31, D[31], q32, D32, CLK, Ai, Bi, Ci);

	input wire A4;
	input wire A0;
	input wire A1;
	input wire A2;
	input wire A3;
	output wire q0;
	input wire D0;
	output wire q1;
	input wire D1;
	output wire q2;
	input wire D2;
	output wire q3;
	input wire D3;
	output wire q4;
	input wire D4;
	output wire q5;
	input wire D5;
	output wire q6;
	input wire D6;
	output wire q7;
	input wire D7;
	output wire q8;
	input wire D8;
	output wire q9;
	input wire D9;
	output wire q10;
	input wire D10;
	output wire q11;
	input wire D11;
	output wire q12;
	input wire D12;
	output wire q13;
	input wire D13;
	output wire q14;
	input wire D14;
	output wire q15;
	input wire D15;
	output wire q16;
	input wire D16;
	output wire q17;
	input wire D17;
	output wire q18;
	input wire D18;
	output wire q19;
	input wire D19;
	output wire q20;
	input wire D20;
	output wire q21;
	input wire D21;
	output wire q22;
	input wire D22;
	output wire q23;
	input wire D23;
	output wire q24;
	input wire D24;
	output wire q25;
	input wire D25;
	output wire q26;
	input wire D26;
	output wire q26;
	input wire D26;
	output wire q27;
	input wire D27;
	output wire q28;
	input wire D28;
	output wire q29;
	input wire D29;
	output wire q30;
	input wire D30;
	output wire q31;
	input wire D[31];
	output wire q32;
	input wire D32;
	input wire CLK;
	input wire Ai;
	input wire Bi;
	input wire Ci;

endmodule // vdp_att_temp_ram

module vdp_vsram (  CLK, D10, q10, D9, q9, D8, q8, D7, q7, D6, q6, D5, q5, D4, q4, D3, q3, D2, q2, D1, q1, D0, q0, A1, A2, A3, A4, A5, A0, Ai, Bi);

	input wire CLK;
	input wire D10;
	output wire q10;
	input wire D9;
	output wire q9;
	input wire D8;
	output wire q8;
	input wire D7;
	output wire q7;
	input wire D6;
	output wire q6;
	input wire D5;
	output wire q5;
	input wire D4;
	output wire q4;
	input wire D3;
	output wire q3;
	input wire D2;
	output wire q2;
	input wire D1;
	output wire q1;
	input wire D0;
	output wire q0;
	input wire A1;
	input wire A2;
	input wire A3;
	input wire A4;
	input wire A5;
	input wire A0;
	input wire Ai;
	input wire Bi;

endmodule // vdp_vsram

module vdp_H_PLA (  HPLA0, HPLA1, HPLA2, HPLA3, HPLA4, HPLA5, HPLA7, HPLA8, HPLA9, HPLA6, HPLA10, HPLA11, HPLA16, HPLA15, HPLA14, HPLA13, HPLA12, i0, HPLA17, HPLA18, HPLA19, HPLA20, HPLA21, HPLA22, Hcnt0, Hcnt1, Hcnt2, Hcnt3, Hcnt4, Hcnt5, Hcnt6, Hcnt7, Hcnt8, H40, M5, B, C, A, HPLA23, HPLA24, HPLA25, HPLA26, HPLA27, HPLA28, HPLA29, HPLA30, HPLA31, HPLA32, HPLA33, i3, HPLA35, HPLA36, HPLA34);

	output wire HPLA0;
	output wire HPLA1;
	output wire HPLA2;
	output wire HPLA3;
	output wire HPLA4;
	output wire HPLA5;
	output wire HPLA7;
	output wire HPLA8;
	output wire HPLA9;
	output wire HPLA6;
	output wire HPLA10;
	output wire HPLA11;
	output wire HPLA16;
	output wire HPLA15;
	output wire HPLA14;
	output wire HPLA13;
	output wire HPLA12;
	input wire i0;
	output wire HPLA17;
	output wire HPLA18;
	output wire HPLA19;
	output wire HPLA20;
	output wire HPLA21;
	output wire HPLA22;
	input wire Hcnt0;
	input wire Hcnt1;
	input wire Hcnt2;
	input wire Hcnt3;
	input wire Hcnt4;
	input wire Hcnt5;
	input wire Hcnt6;
	input wire Hcnt7;
	input wire Hcnt8;
	input wire H40;
	input wire M5;
	input wire B;
	input wire C;
	input wire A;
	output wire HPLA23;
	output wire HPLA24;
	output wire HPLA25;
	output wire HPLA26;
	output wire HPLA27;
	output wire HPLA28;
	output wire HPLA29;
	output wire HPLA30;
	output wire HPLA31;
	output wire HPLA32;
	output wire HPLA33;
	input wire i3;
	output wire HPLA35;
	output wire HPLA36;
	output wire HPLA34;

endmodule // vdp_H_PLA



// ERROR: conflicting wire AD_DATA[7]
// ERROR: conflicting wire AD_DATA[6]
// ERROR: conflicting wire AD_DATA[4]
// ERROR: conflicting wire RD_DATA[2]
// ERROR: conflicting wire RD_DATA[1]
// ERROR: conflicting wire RD_DATA[0]
// ERROR: conflicting wire AD_DATA[5]
// ERROR: conflicting wire DB[0]
// ERROR: conflicting wire DB[1]
// ERROR: conflicting wire DB[2]
// ERROR: conflicting wire DB[3]
// ERROR: conflicting wire DB[4]
// ERROR: conflicting wire DB[5]
// ERROR: conflicting wire DB[6]
// ERROR: conflicting wire DB[7]
// ERROR: conflicting wire DB[8]
// ERROR: conflicting wire DB[9]
// ERROR: conflicting wire AD_DATA[3]
// ERROR: conflicting wire AD_DATA[2]
// ERROR: conflicting wire AD_DATA[1]
// ERROR: conflicting wire AD_DATA[0]
// ERROR: conflicting wire DB[14]
// ERROR: conflicting wire DB[13]
// ERROR: conflicting wire DB[12]
// ERROR: conflicting wire DB[11]
// ERROR: conflicting wire DB[10]
// ERROR: floating wire w172
// ERROR: conflicting wire RD_DATA[4]
// ERROR: floating wire w203
// ERROR: conflicting wire RD_DATA[6]
// ERROR: floating wire w219
// ERROR: conflicting wire w235
// ERROR: conflicting wire w242
// ERROR: conflicting wire w276
// ERROR: conflicting wire w284
// ERROR: conflicting wire w300
// ERROR: floating wire w313
// ERROR: conflicting wire RD_DATA[5]
// ERROR: floating wire w329
// ERROR: conflicting wire DB[15]
// ERROR: conflicting wire w334
// ERROR: floating wire w427
// ERROR: conflicting wire VRAMA[0]
// ERROR: floating wire w540
// ERROR: conflicting wire VRAMA[8]
// ERROR: conflicting wire VRAMA[7]
// ERROR: conflicting wire VRAMA[9]
// ERROR: conflicting wire VRAMA[10]
// ERROR: conflicting wire VRAMA[6]
// ERROR: conflicting wire VRAMA[5]
// ERROR: conflicting wire VRAMA[11]
// ERROR: conflicting wire VRAMA[12]
// ERROR: conflicting wire VRAMA[4]
// ERROR: conflicting wire VRAMA[13]
// ERROR: conflicting wire VRAMA[3]
// ERROR: conflicting wire VRAMA[14]
// ERROR: conflicting wire VRAMA[2]
// ERROR: conflicting wire VRAMA[15]
// ERROR: conflicting wire VRAMA[1]
// ERROR: conflicting wire VRAMA[16]
// ERROR: floating wire w752
// ERROR: floating wire w754
// ERROR: floating wire w772
// ERROR: floating wire w773
// ERROR: floating wire w1032
// ERROR: conflicting wire COL[1]
// ERROR: conflicting wire COL[0]
// ERROR: conflicting wire COL[2]
// ERROR: conflicting wire COL[3]
// ERROR: conflicting wire COL[4]
// ERROR: conflicting wire COL[6]
// ERROR: conflicting wire COL[5]
// ERROR: floating wire w1051
// ERROR: floating wire w1052
// ERROR: floating wire w1173
// ERROR: floating wire w1243
// ERROR: floating wire w1250
// ERROR: floating wire w1258
// ERROR: floating wire w1302
// ERROR: floating wire w1324
// ERROR: conflicting wire w1396
// ERROR: conflicting wire w1465
// ERROR: conflicting wire w1466
// ERROR: floating wire w1516
// ERROR: conflicting wire w1549
// ERROR: floating wire w1553
// ERROR: floating wire w1619
// ERROR: floating wire w1716
// ERROR: floating wire w1747
// ERROR: floating wire w1759
// ERROR: floating wire w1769
// ERROR: floating wire w1906
// ERROR: floating wire w1998
// ERROR: floating wire w2184
// ERROR: floating wire w2219
// ERROR: floating wire w2396
// ERROR: floating wire w2540
// ERROR: floating wire w2546
// ERROR: floating wire w2700
// ERROR: floating wire w3003
// ERROR: floating wire w3013
// ERROR: floating wire w3345
// ERROR: floating wire w3404
// ERROR: floating wire w3484
// ERROR: floating wire w3540
// ERROR: floating wire w3581
// ERROR: floating wire w3621
// ERROR: floating wire w3626
// ERROR: floating wire w3680
// ERROR: floating wire w3682
// ERROR: floating wire w3755
// ERROR: floating wire w3781
// ERROR: floating wire w3832
// ERROR: floating wire w3948
// ERROR: floating wire w4280
// ERROR: floating wire w4290
// ERROR: floating wire w4441
// ERROR: floating wire w4503
// ERROR: floating wire w4508
// ERROR: floating wire w4545
// ERROR: floating wire w4604
// ERROR: floating wire w4609
// ERROR: floating wire w4638
// ERROR: floating wire w4683
// ERROR: floating wire w4742
// ERROR: floating wire w4748
// ERROR: floating wire w4793
// ERROR: floating wire w4978
// ERROR: floating wire w5033
// ERROR: floating wire w5160
// ERROR: floating wire w5168
// ERROR: floating wire w5182
// ERROR: floating wire w5328
// ERROR: floating wire w5376
// ERROR: floating wire w5562
// ERROR: floating wire w5699
// ERROR: floating wire w5701
// ERROR: floating wire w5795
// ERROR: floating wire w5937
// ERROR: floating wire w5952
// ERROR: floating wire w5983
// ERROR: floating wire w6028
// ERROR: floating wire w6065
// ERROR: floating wire w6074
// ERROR: floating wire w6075
// ERROR: floating wire w6319
// ERROR: floating wire w6435
// ERROR: floating wire w6437
// ERROR: floating wire w6438
// ERROR: floating wire w6584
// WARNING: Cell vdp_fa:g385 port CO not connected.
// WARNING: Cell vdp_and:g527 port Z not connected.
// WARNING: Cell vdp_cnt_bit_load:g871 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g873 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g1405 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g1406 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1407 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1408 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1409 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1410 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1411 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1412 port Q not connected.
// WARNING: Cell vdp_or:g1576 port Z not connected.
// WARNING: Cell vdp_cnt_bit_load:g1959 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g1960 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2145 port CO not connected.
// WARNING: Cell vdp_ha:g2278 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2280 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2282 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2284 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2286 port CO not connected.
// WARNING: Cell vdp_rs_ff:g2380 port nQ not connected.
// WARNING: Cell vdp_rs_ff:g2381 port nQ not connected.
// WARNING: Cell vdp_comp_we:g2612 port nZ not connected.
// WARNING: Cell vdp_comp_we:g2701 port nZ not connected.
// WARNING: Cell vdp_fa:g3842 port CO not connected.
// WARNING: Cell vdp_fa:g4058 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g4437 port CO not connected.
// WARNING: Cell vdp_fa:g4453 port CO not connected.
// WARNING: Cell vdp_fa:g4463 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g5851 port CO not connected.
// WARNING: Cell vdp_fa:g5862 port CO not connected.
// WARNING: Cell vdp_fa:g5888 port CO not connected.
// WARNING: Cell vdp_fa:g5892 port CO not connected.
// WARNING: Cell vdp_fa:g6086 port CO not connected.
// WARNING: Cell vdp_ha:g6137 port CO not connected.
// WARNING: Cell vdp_sr_bit:g6146 port Q not connected.
// WARNING: Cell vdp_fa:g6150 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g6216 port CO not connected.
