module IO (  VD15_i, VD15_d, VD15_o, VA1_i, VA1_d, VA1_o, VA2_i, VA2_d, VA2_o, VA3_i, VA3_d, VA3_o, VA4_i, VA4_d, VA4_o, VA5_i, VA5_d, VA5_o, VA6_i, VA6_d, VA6_o, VA7_i, VA7_d, VA7_o, n_FRES, n_DISK, PC0_i, PC0_d, PC0_o, PC1_i, PC1_d, PC1_o, PC2_i, PC2_d, PC2_o, PC3_i, PC3_d, PC3_o, PC4_i, PC4_d, PC4_o, PC5_i, PC5_d, PC5_o, PC6_i, PC6_d, PC6_o, TEST, n_HL, n_LWR, n_CAS0, VCLK, n_JAP, NTSC, n_M3, n_IO, n_SRES, n_ZTOV, n_VTOZ, ZD7_i, ZD7_d, ZD7_o, ZD6_i, ZD6_d, ZD6_o, ZD5_i, ZD5_d, ZD5_o, ZD4_i, ZD4_d, ZD4_o, ZD3_i, ZD3_d, ZD3_o, ZD2_i, ZD2_d, ZD2_o, ZD1_i, ZD1_d, ZD1_o, ZD0_i, ZD0_d, ZD0_o, ZA0, ZA1_i, ZA1_d, ZA1_o, ZA2_i, ZA2_d, ZA2_o, ZA3_i, ZA3_d, ZA3_o, ZA4_i, ZA4_d, ZA4_o, ZA5_i, ZA5_d, ZA5_o, ZA6_i, ZA6_d, ZA6_o, ZA7_i, ZA7_d, ZA7_o, PA0_i, PA0_d, PA0_o, PA1_i, PA1_d, PA1_o, PA2_i, PA2_d, PA2_o, PA3_i, PA3_d, PA3_o, PA4_i, PA4_d, PA4_o, PA5_i, PA5_d, PA5_o, PA6_i, PA6_d, PA6_o, PB0_i, PB0_d, PB0_o, PB1_i, PB1_d, PB1_o, PB2_i, PB2_d, PB2_o, PB3_i, PB3_d, PB3_o, PB4_i, PB4_d, PB4_o, PB5_i, PB5_d, PB5_o, PB6_i, PB6_d, PB6_o, VD0_i, VD0_d, VD0_o, VD1_i, VD1_d, VD1_o, VD2_i, VD2_d, VD2_o, VD3_i, VD3_d, VD3_o, VD4_i, VD4_d, VD4_o, VD5_i, VD5_d, VD5_o, VD6_i, VD6_d, VD6_o, VD7_i, VD7_d, VD7_o, VD8_i, VD8_d, VD8_o, VD9_i, VD9_d, VD9_o, VD10_i, VD10_d, VD10_o, VD11_i, VD11_d, VD11_o, VD12_i, VD12_d, VD12_o, VD13_i, VD13_d, VD13_o, VD14_i, VD14_d, VD14_o);

	input wire VD15_i;
	output wire VD15_d;
	output wire VD15_o;
	input wire VA1_i;
	output wire VA1_d;
	output wire VA1_o;
	input wire VA2_i;
	output wire VA2_d;
	output wire VA2_o;
	input wire VA3_i;
	output wire VA3_d;
	output wire VA3_o;
	input wire VA4_i;
	output wire VA4_d;
	output wire VA4_o;
	input wire VA5_i;
	output wire VA5_d;
	output wire VA5_o;
	input wire VA6_i;
	output wire VA6_d;
	output wire VA6_o;
	input wire VA7_i;
	output wire VA7_d;
	output wire VA7_o;
	output wire n_FRES;
	input wire n_DISK;
	input wire PC0_i;
	output wire PC0_d;
	output wire PC0_o;
	input wire PC1_i;
	output wire PC1_d;
	output wire PC1_o;
	input wire PC2_i;
	output wire PC2_d;
	output wire PC2_o;
	input wire PC3_i;
	output wire PC3_d;
	output wire PC3_o;
	input wire PC4_i;
	output wire PC4_d;
	output wire PC4_o;
	input wire PC5_i;
	output wire PC5_d;
	output wire PC5_o;
	input wire PC6_i;
	output wire PC6_d;
	output wire PC6_o;
	input wire TEST;
	output wire n_HL;
	input wire n_LWR;
	input wire n_CAS0;
	input wire VCLK;
	input wire n_JAP;
	input wire NTSC;
	input wire n_M3;
	input wire n_IO;
	input wire n_SRES;
	input wire n_ZTOV;
	input wire n_VTOZ;
	input wire ZD7_i;
	output wire ZD7_d;
	output wire ZD7_o;
	input wire ZD6_i;
	output wire ZD6_d;
	output wire ZD6_o;
	input wire ZD5_i;
	output wire ZD5_d;
	output wire ZD5_o;
	input wire ZD4_i;
	output wire ZD4_d;
	output wire ZD4_o;
	input wire ZD3_i;
	output wire ZD3_d;
	output wire ZD3_o;
	input wire ZD2_i;
	output wire ZD2_d;
	output wire ZD2_o;
	input wire ZD1_i;
	output wire ZD1_d;
	output wire ZD1_o;
	input wire ZD0_i;
	output wire ZD0_d;
	output wire ZD0_o;
	input wire ZA0;
	input wire ZA1_i;
	output wire ZA1_d;
	output wire ZA1_o;
	input wire ZA2_i;
	output wire ZA2_d;
	output wire ZA2_o;
	input wire ZA3_i;
	output wire ZA3_d;
	output wire ZA3_o;
	input wire ZA4_i;
	output wire ZA4_d;
	output wire ZA4_o;
	input wire ZA5_i;
	output wire ZA5_d;
	output wire ZA5_o;
	input wire ZA6_i;
	output wire ZA6_d;
	output wire ZA6_o;
	input wire ZA7_i;
	output wire ZA7_d;
	output wire ZA7_o;
	input wire PA0_i;
	output wire PA0_d;
	output wire PA0_o;
	input wire PA1_i;
	output wire PA1_d;
	output wire PA1_o;
	input wire PA2_i;
	output wire PA2_d;
	output wire PA2_o;
	input wire PA3_i;
	output wire PA3_d;
	output wire PA3_o;
	input wire PA4_i;
	output wire PA4_d;
	output wire PA4_o;
	input wire PA5_i;
	output wire PA5_d;
	output wire PA5_o;
	input wire PA6_i;
	output wire PA6_d;
	output wire PA6_o;
	input wire PB0_i;
	output wire PB0_d;
	output wire PB0_o;
	input wire PB1_i;
	output wire PB1_d;
	output wire PB1_o;
	input wire PB2_i;
	output wire PB2_d;
	output wire PB2_o;
	input wire PB3_i;
	output wire PB3_d;
	output wire PB3_o;
	input wire PB4_i;
	output wire PB4_d;
	output wire PB4_o;
	input wire PB5_i;
	output wire PB5_d;
	output wire PB5_o;
	input wire PB6_i;
	output wire PB6_d;
	output wire PB6_o;
	input wire VD0_i;
	output wire VD0_d;
	output wire VD0_o;
	input wire VD1_i;
	output wire VD1_d;
	output wire VD1_o;
	input wire VD2_i;
	output wire VD2_d;
	output wire VD2_o;
	input wire VD3_i;
	output wire VD3_d;
	output wire VD3_o;
	input wire VD4_i;
	output wire VD4_d;
	output wire VD4_o;
	input wire VD5_i;
	output wire VD5_d;
	output wire VD5_o;
	input wire VD6_i;
	output wire VD6_d;
	output wire VD6_o;
	input wire VD7_i;
	output wire VD7_d;
	output wire VD7_o;
	input wire VD8_i;
	output wire VD8_d;
	output wire VD8_o;
	input wire VD9_i;
	output wire VD9_d;
	output wire VD9_o;
	input wire VD10_i;
	output wire VD10_d;
	output wire VD10_o;
	input wire VD11_i;
	output wire VD11_d;
	output wire VD11_o;
	input wire VD12_i;
	output wire VD12_d;
	output wire VD12_o;
	input wire VD13_i;
	output wire VD13_d;
	output wire VD13_o;
	input wire VD14_i;
	output wire VD14_d;
	output wire VD14_o;

	// Wires

	wire w1;
	wire w2;
	wire w3;
	wire w4;
	wire w5;
	wire w6;
	wire w7;
	wire w8;
	wire w9;
	wire w10;
	wire w11;
	wire w12;
	wire w13;
	wire w14;
	wire w15;
	wire w16;
	wire w17;
	wire w18;
	wire w19;
	wire w20;
	wire w21;
	wire w22;
	wire w23;
	wire w24;
	wire w25;
	wire w26;
	wire w27;
	wire w28;
	wire w29;
	wire w30;
	wire w31;
	wire w32;
	wire w33;
	wire w34;
	wire w35;
	wire w36;
	wire w37;
	wire w38;
	wire w39;
	wire w40;
	wire w41;
	wire w42;
	wire w43;
	wire w44;
	wire w45;
	wire w46;
	wire w47;
	wire w48;
	wire w49;
	wire w50;
	wire w51;
	wire w52;
	wire w53;
	wire w54;
	wire w55;
	wire w56;
	wire w57;
	wire w58;
	wire w59;
	wire w60;
	wire w61;
	wire w62;
	wire w63;
	wire w64;
	wire w65;
	wire w66;
	wire w67;
	wire w68;
	wire w69;
	wire w70;
	wire w71;
	wire w72;
	wire w73;
	wire w74;
	wire w75;
	wire w76;
	wire w77;
	wire w78;
	wire w79;
	wire w80;
	wire w81;
	wire w82;
	wire w83;
	wire w84;
	wire w85;
	wire w86;
	wire w87;
	wire w88;
	wire w89;
	wire w90;
	wire w91;
	wire w92;
	wire w93;
	wire w94;
	wire w95;
	wire w96;
	wire w97;
	wire w98;
	wire w99;
	wire w100;
	wire w101;
	wire w102;
	wire w103;
	wire w104;
	wire w105;
	wire w106;
	wire w107;
	wire w108;
	wire w109;
	wire w110;
	wire w111;
	wire w112;
	wire w113;
	wire w114;
	wire w115;
	wire w116;
	wire w117;
	wire w118;
	wire w119;
	wire w120;
	wire w121;
	wire w122;
	wire w123;
	wire w124;
	wire w125;
	wire w126;
	wire w127;
	wire w128;
	wire w129;
	wire w130;
	wire w131;
	wire w132;
	wire w133;
	wire w134;
	wire w135;
	wire w136;
	wire w137;
	wire w138;
	wire w139;
	wire w140;
	wire w141;
	wire w142;
	wire w143;
	wire w144;
	wire w145;
	wire w146;
	wire w147;
	wire w148;
	wire w149;
	wire w150;
	wire w151;
	wire w152;
	wire w153;
	wire w154;
	wire w155;
	wire w156;
	wire w157;
	wire w158;
	wire w159;
	wire w160;
	wire w161;
	wire w162;
	wire w163;
	wire w164;
	wire w165;
	wire w166;
	wire w167;
	wire w168;
	wire w169;
	wire w170;
	wire w171;
	wire w172;
	wire w173;
	wire w174;
	wire w175;
	wire w176;
	wire w177;
	wire w178;
	wire w179;
	wire w180;
	wire w181;
	wire w182;
	wire w183;
	wire w184;
	wire w185;
	wire w186;
	wire w187;
	wire w188;
	wire w189;
	wire w190;
	wire w191;
	wire w192;
	wire w193;
	wire w194;
	wire w195;
	wire w196;
	wire w197;
	wire w198;
	wire w199;
	wire w200;
	wire w201;
	wire w202;
	wire w203;
	wire w204;
	wire w205;
	wire w206;
	wire w207;
	wire w208;
	wire w209;
	wire w210;
	wire w211;
	wire w212;
	wire w213;
	wire w214;
	wire w215;
	wire w216;
	wire w217;
	wire w218;
	wire w219;
	wire w220;
	wire w221;
	wire w222;
	wire w223;
	wire w224;
	wire w225;
	wire w226;
	wire w227;
	wire w228;
	wire w229;
	wire w230;
	wire w231;
	wire w232;
	wire w233;
	wire w234;
	wire w235;
	wire w236;
	wire w237;
	wire w238;
	wire w239;
	wire w240;
	wire w241;
	wire w242;
	wire w243;
	wire w244;
	wire w245;
	wire w246;
	wire w247;
	wire w248;
	wire w249;
	wire w250;
	wire w251;
	wire w252;
	wire w253;
	wire w254;
	wire w255;
	wire w256;
	wire w257;
	wire w258;
	wire w259;
	wire w260;
	wire w261;
	wire w262;
	wire w263;
	wire w264;
	wire w265;
	wire w266;
	wire w267;
	wire w268;
	wire w269;
	wire w270;
	wire w271;
	wire w272;
	wire w273;
	wire w274;
	wire w275;
	wire w276;
	wire w277;
	wire w278;
	wire w279;
	wire w280;
	wire w281;
	wire w282;
	wire w283;
	wire w284;
	wire w285;
	wire w286;
	wire w287;
	wire w288;
	wire w289;
	wire w290;
	wire w291;
	wire w292;
	wire w293;
	wire w294;
	wire w295;
	wire w296;
	wire w297;
	wire w298;
	wire w299;
	wire w300;
	wire w301;
	wire w302;
	wire w303;
	wire w304;
	wire w305;
	wire w306;
	wire w307;
	wire w308;
	wire w309;
	wire w310;
	wire w311;
	wire w312;
	wire w313;
	wire w314;
	wire w315;
	wire w316;
	wire w317;
	wire w318;
	wire w319;
	wire w320;
	wire w321;
	wire w322;
	wire w323;
	wire w324;
	wire w325;
	wire w326;
	wire w327;
	wire w328;
	wire w329;
	wire w330;
	wire w331;
	wire w332;
	wire w333;
	wire w334;
	wire w335;
	wire w336;
	wire w337;
	wire w338;
	wire w339;
	wire w340;
	wire w341;
	wire w342;
	wire w343;
	wire w344;
	wire w345;
	wire w346;
	wire w347;
	wire w348;
	wire w349;
	wire w350;
	wire w351;
	wire w352;
	wire w353;
	wire w354;
	wire w355;
	wire w356;
	wire w357;
	wire w358;
	wire w359;
	wire w360;
	wire w361;
	wire w362;
	wire w363;
	wire w364;
	wire w365;
	wire w366;
	wire w367;
	wire w368;
	wire w369;
	wire w370;
	wire w371;
	wire w372;
	wire w373;
	wire w374;
	wire w375;
	wire w376;
	wire w377;
	wire w378;
	wire w379;
	wire w380;
	wire w381;
	wire w382;
	wire w383;
	wire w384;
	wire w385;
	wire w386;
	wire w387;
	wire w388;
	wire w389;
	wire w390;
	wire w391;
	wire w392;
	wire w393;
	wire w394;
	wire w395;
	wire w396;
	wire w397;
	wire w398;
	wire w399;
	wire w400;
	wire w401;
	wire w402;
	wire w403;
	wire w404;
	wire w405;
	wire w406;
	wire w407;
	wire w408;
	wire w409;
	wire w410;
	wire w411;
	wire w412;
	wire w413;
	wire w414;
	wire w415;
	wire w416;
	wire w417;
	wire w418;
	wire w419;
	wire w420;
	wire w421;
	wire w422;
	wire w423;
	wire w424;
	wire w425;
	wire w426;
	wire w427;
	wire w428;
	wire w429;
	wire w430;
	wire w431;
	wire w432;
	wire w433;
	wire w434;
	wire w435;
	wire w436;
	wire w437;
	wire w438;
	wire w439;
	wire w440;
	wire w441;
	wire w442;
	wire w443;
	wire w444;
	wire w445;
	wire w446;
	wire w447;
	wire w448;
	wire w449;
	wire w450;
	wire w451;
	wire w452;
	wire w453;
	wire w454;
	wire w455;
	wire w456;
	wire w457;
	wire w458;
	wire w459;
	wire w460;
	wire w461;
	wire w462;
	wire w463;
	wire w464;
	wire w465;
	wire w466;
	wire w467;
	wire w468;
	wire w469;
	wire w470;
	wire w471;
	wire w472;
	wire w473;
	wire w474;
	wire w475;
	wire w476;
	wire w477;
	wire w478;
	wire w479;
	wire w480;
	wire w481;
	wire w482;
	wire w483;
	wire w484;
	wire w485;
	wire w486;
	wire w487;
	wire w488;
	wire w489;
	wire w490;
	wire w491;
	wire w492;
	wire w493;
	wire w494;
	wire w495;
	wire w496;
	wire w497;
	wire w498;
	wire w499;
	wire w500;
	wire w501;
	wire w502;
	wire w503;
	wire w504;
	wire w505;
	wire w506;
	wire w507;
	wire w508;
	wire w509;
	wire w510;
	wire w511;
	wire w512;
	wire w513;
	wire w514;
	wire w515;
	wire w516;
	wire w517;
	wire w518;
	wire w519;
	wire w520;
	wire w521;
	wire w522;
	wire w523;
	wire w524;
	wire w525;
	wire w526;
	wire w527;
	wire w528;
	wire w529;
	wire w530;
	wire w531;
	wire w532;
	wire w533;
	wire w534;
	wire w535;
	wire w536;
	wire w537;
	wire w538;
	wire w539;
	wire w540;
	wire w541;
	wire w542;
	wire w543;
	wire w544;
	wire w545;
	wire w546;
	wire w547;
	wire w548;
	wire w549;
	wire w550;
	wire w551;
	wire w552;
	wire w553;
	wire w554;
	wire w555;
	wire w556;
	wire w557;
	wire w558;
	wire w559;
	wire w560;
	wire w561;
	wire w562;
	wire w563;
	wire w564;
	wire w565;
	wire w566;
	wire w567;
	wire w568;
	wire w569;
	wire w570;
	wire w571;
	wire w572;
	wire w573;
	wire w574;
	wire w575;
	wire w576;
	wire w577;
	wire w578;
	wire w579;
	wire w580;
	wire w581;
	wire w582;
	wire w583;
	wire w584;
	wire w585;
	wire w586;
	wire w587;
	wire w588;
	wire w589;
	wire w590;
	wire w591;
	wire w592;
	wire w593;
	wire w594;
	wire w595;
	wire w596;
	wire w597;
	wire w598;
	wire w599;
	wire w600;
	wire w601;
	wire w602;
	wire w603;
	wire w604;
	wire w605;
	wire w606;
	wire w607;
	wire w608;
	wire w609;
	wire w610;
	wire w611;
	wire w612;
	wire w613;
	wire w614;
	wire w615;
	wire w616;
	wire w617;
	wire w618;
	wire w619;
	wire w620;
	wire w621;
	wire w622;
	wire w623;
	wire w624;
	wire w625;
	wire w626;
	wire w627;
	wire w628;
	wire w629;
	wire w630;
	wire w631;
	wire w632;
	wire w633;
	wire w634;
	wire w635;
	wire w636;
	wire w637;
	wire w638;
	wire w639;
	wire w640;
	wire w641;
	wire w642;
	wire w643;
	wire w644;
	wire w645;
	wire w646;
	wire w647;
	wire w648;
	wire w649;
	wire w650;
	wire w651;
	wire w652;
	wire w653;
	wire w654;
	wire w655;
	wire w656;
	wire w657;
	wire w658;
	wire w659;
	wire w660;
	wire w661;
	wire w662;
	wire w663;
	wire w664;
	wire w665;
	wire w666;
	wire w667;
	wire w668;
	wire w669;
	wire w670;
	wire w671;
	wire w672;
	wire w673;
	wire w674;
	wire w675;
	wire w676;
	wire w677;
	wire w678;
	wire w679;
	wire w680;
	wire w681;
	wire w682;
	wire w683;
	wire w684;
	wire w685;
	wire w686;
	wire w687;
	wire w688;
	wire w689;
	wire w690;
	wire w691;
	wire w692;
	wire w693;
	wire w694;
	wire w695;
	wire w696;
	wire w697;
	wire w698;
	wire w699;
	wire w700;
	wire w701;
	wire w702;
	wire w703;
	wire w704;
	wire w705;
	wire w706;
	wire w707;
	wire w708;
	wire w709;
	wire w710;
	wire w711;
	wire w712;
	wire w713;
	wire w714;
	wire w715;
	wire w716;
	wire w717;
	wire w718;
	wire w719;
	wire w720;
	wire w721;
	wire w722;
	wire w723;
	wire w724;
	wire w725;
	wire w726;
	wire w727;
	wire w728;
	wire w729;
	wire w730;
	wire w731;
	wire w732;
	wire w733;
	wire w734;
	wire w735;
	wire w736;
	wire w737;
	wire w738;
	wire w739;
	wire w740;
	wire w741;
	wire w742;
	wire w743;
	wire w744;
	wire w745;
	wire w746;
	wire w747;
	wire w748;
	wire w749;
	wire w750;
	wire w751;
	wire w752;
	wire w753;
	wire w754;
	wire w755;
	wire w756;
	wire w757;
	wire w758;
	wire w759;
	wire w760;
	wire w761;
	wire w762;
	wire w763;
	wire w764;
	wire w765;
	wire w766;
	wire w767;
	wire w768;
	wire w769;
	wire w770;
	wire w771;
	wire w772;
	wire w773;
	wire w774;
	wire w775;
	wire w776;
	wire w777;
	wire w778;
	wire w779;
	wire w780;
	wire w781;
	wire w782;
	wire w783;
	wire w784;
	wire w785;
	wire w786;
	wire w787;
	wire w788;
	wire w789;
	wire w790;
	wire w791;
	wire w792;
	wire w793;
	wire w794;
	wire w795;
	wire w796;
	wire w797;
	wire w798;
	wire w799;
	wire w800;
	wire w801;
	wire w802;
	wire w803;
	wire w804;
	wire w805;
	wire w806;
	wire w807;
	wire w808;
	wire w809;
	wire w810;
	wire w811;
	wire w812;
	wire w813;
	wire w814;
	wire w815;
	wire w816;
	wire w817;
	wire w818;
	wire w819;
	wire w820;
	wire w821;
	wire w822;
	wire w823;
	wire w824;
	wire w825;
	wire w826;
	wire w827;
	wire w828;
	wire w829;
	wire w830;
	wire w831;
	wire w832;
	wire w833;
	wire w834;
	wire w835;
	wire w836;
	wire w837;
	wire w838;
	wire w839;
	wire w840;
	wire w841;
	wire w842;
	wire w843;
	wire w844;
	wire w845;
	wire w846;
	wire w847;
	wire w848;
	wire w849;
	wire w850;
	wire w851;
	wire w852;
	wire w853;
	wire w854;
	wire w855;
	wire w856;
	wire w857;
	wire w858;
	wire w859;
	wire w860;
	wire w861;
	wire w862;
	wire w863;
	wire w864;
	wire w865;
	wire w866;
	wire w867;
	wire w868;
	wire w869;
	wire w870;
	wire w871;
	wire w872;
	wire w873;
	wire w874;
	wire w875;
	wire w876;
	wire w877;
	wire w878;
	wire w879;
	wire w880;
	wire w881;
	wire w882;
	wire w883;
	wire w884;
	wire w885;
	wire w886;
	wire w887;
	wire w888;
	wire w889;
	wire w890;
	wire w891;
	wire w892;
	wire w893;
	wire w894;
	wire w895;
	wire w896;
	wire w897;
	wire w898;
	wire w899;
	wire w900;
	wire w901;
	wire w902;
	wire w903;
	wire w904;
	wire w905;
	wire w906;
	wire w907;
	wire w908;
	wire w909;
	wire w910;
	wire w911;
	wire w912;
	wire w913;
	wire w914;
	wire w915;
	wire w916;
	wire w917;
	wire w918;
	wire w919;
	wire w920;
	wire w921;
	wire w922;
	wire w923;
	wire w924;
	wire w925;
	wire w926;
	wire w927;
	wire w928;
	wire w929;
	wire w930;
	wire w931;
	wire w932;
	wire w933;
	wire w934;
	wire w935;
	wire w936;

	assign w217 = VD15_i;
	assign VD15_d = w208;
	assign VD15_o = w205;
	assign w57 = VA1_i;
	assign VA1_d = w291;
	assign VA1_o = w224;
	assign w54 = VA2_i;
	assign VA2_d = w291;
	assign VA2_o = w223;
	assign w66 = VA3_i;
	assign VA3_d = w291;
	assign VA3_o = w55;
	assign w102 = VA4_i;
	assign VA4_d = w291;
	assign VA4_o = w222;
	assign w103 = VA5_i;
	assign VA5_d = w291;
	assign VA5_o = w88;
	assign w104 = VA6_i;
	assign VA6_d = w291;
	assign VA6_o = w246;
	assign w106 = VA7_i;
	assign VA7_d = w291;
	assign VA7_o = w259;
	assign n_FRES = w300;
	assign w306 = n_DISK;
	assign w307 = PC0_i;
	assign PC0_d = w308;
	assign PC0_o = w330;
	assign w157 = PC1_i;
	assign PC1_d = w310;
	assign PC1_o = w309;
	assign w257 = PC2_i;
	assign PC2_d = w331;
	assign PC2_o = w311;
	assign w314 = PC3_i;
	assign PC3_d = w313;
	assign PC3_o = w312;
	assign w317 = PC4_i;
	assign PC4_d = w316;
	assign PC4_o = w315;
	assign w318 = PC5_i;
	assign PC5_d = w319;
	assign PC5_o = w320;
	assign w321 = PC6_i;
	assign PC6_d = w322;
	assign PC6_o = w323;
	assign w324 = TEST;
	assign n_HL = w245;
	assign w325 = n_LWR;
	assign w268 = n_CAS0;
	assign w115 = VCLK;
	assign w153 = n_JAP;
	assign w293 = NTSC;
	assign w8 = n_M3;
	assign w266 = n_IO;
	assign w292 = n_SRES;
	assign w291 = n_ZTOV;
	assign w98 = n_VTOZ;
	assign w289 = ZD7_i;
	assign ZD7_d = w232;
	assign ZD7_o = w290;
	assign w288 = ZD6_i;
	assign ZD6_d = w232;
	assign ZD6_o = w287;
	assign w286 = ZD5_i;
	assign ZD5_d = w232;
	assign ZD5_o = w285;
	assign w283 = ZD4_i;
	assign ZD4_d = w232;
	assign ZD4_o = w284;
	assign w229 = ZD3_i;
	assign ZD3_d = w232;
	assign ZD3_o = w278;
	assign w280 = ZD2_i;
	assign ZD2_d = w232;
	assign ZD2_o = w279;
	assign w228 = ZD1_i;
	assign ZD1_d = w232;
	assign ZD1_o = w281;
	assign w226 = ZD0_i;
	assign ZD0_d = w232;
	assign ZD0_o = w282;
	assign w188 = ZA0;
	assign w35 = ZA1_i;
	assign ZA1_d = w98;
	assign ZA1_o = w57;
	assign w99 = ZA2_i;
	assign ZA2_d = w98;
	assign ZA2_o = w54;
	assign w100 = ZA3_i;
	assign ZA3_d = w98;
	assign ZA3_o = w66;
	assign w101 = ZA4_i;
	assign ZA4_d = w98;
	assign ZA4_o = w102;
	assign w90 = ZA5_i;
	assign ZA5_d = w98;
	assign ZA5_o = w103;
	assign w91 = ZA6_i;
	assign ZA6_d = w98;
	assign ZA6_o = w104;
	assign w105 = ZA7_i;
	assign ZA7_d = w98;
	assign ZA7_o = w106;
	assign w107 = PA0_i;
	assign PA0_d = w84;
	assign PA0_o = w85;
	assign w160 = PA1_i;
	assign PA1_d = w79;
	assign PA1_o = w934;
	assign w258 = PA2_i;
	assign PA2_d = w80;
	assign PA2_o = w81;
	assign w76 = PA3_i;
	assign PA3_d = w83;
	assign PA3_o = w82;
	assign w73 = PA4_i;
	assign PA4_d = w155;
	assign PA4_o = w74;
	assign w71 = PA5_i;
	assign PA5_d = w72;
	assign PA5_o = w75;
	assign w70 = PA6_i;
	assign PA6_d = w69;
	assign PA6_o = w68;
	assign w65 = PB0_i;
	assign PB0_d = w64;
	assign PB0_o = w67;
	assign w63 = PB1_i;
	assign PB1_d = w62;
	assign PB1_o = w58;
	assign w61 = PB2_i;
	assign PB2_d = w60;
	assign PB2_o = w59;
	assign w28 = PB3_i;
	assign PB3_d = w26;
	assign PB3_o = w27;
	assign w242 = PB4_i;
	assign PB4_d = w13;
	assign PB4_o = w15;
	assign w23 = PB5_i;
	assign PB5_d = w25;
	assign PB5_o = w24;
	assign w189 = PB6_i;
	assign PB6_d = w96;
	assign PB6_o = w190;
	assign w191 = VD0_i;
	assign VD0_d = w192;
	assign VD0_o = w193;
	assign w195 = VD1_i;
	assign VD1_d = w192;
	assign VD1_o = w194;
	assign w197 = VD2_i;
	assign VD2_d = w192;
	assign VD2_o = w196;
	assign w198 = VD3_i;
	assign VD3_d = w192;
	assign VD3_o = w213;
	assign w199 = VD4_i;
	assign VD4_d = w192;
	assign VD4_o = w200;
	assign w202 = VD5_i;
	assign VD5_d = w192;
	assign VD5_o = w201;
	assign w204 = VD6_i;
	assign VD6_d = w192;
	assign VD6_o = w203;
	assign w206 = VD7_i;
	assign VD7_d = w192;
	assign VD7_o = w205;
	assign w209 = VD8_i;
	assign VD8_d = w208;
	assign VD8_o = w207;
	assign w210 = VD9_i;
	assign VD9_d = w208;
	assign VD9_o = w194;
	assign w211 = VD10_i;
	assign VD10_d = w208;
	assign VD10_o = w196;
	assign w212 = VD11_i;
	assign VD11_d = w208;
	assign VD11_o = w213;
	assign w214 = VD12_i;
	assign VD12_d = w208;
	assign VD12_o = w200;
	assign w215 = VD13_i;
	assign VD13_d = w208;
	assign VD13_o = w201;
	assign w216 = VD14_i;
	assign VD14_d = w208;
	assign VD14_o = w203;

	// Instances

	io_AND g_1 (.Z(w1), .B(w2), .A(w8) );
	io_OR g_2 (.A(w1), .Z(w129), .B(w10) );
	io_NOR g_3 (.Z(w10), .B(w8), .A(w5) );
	io_NOT g_4 (.A(w9), .nZ(w5) );
	io_OR g_5 (.B(w5), .Z(w12), .A(w6) );
	io_AND g_6 (.Z(w173), .B(w6), .A(w11) );
	io_OR4 g_7 (.Z(w11), .D(w8), .C(w4), .B(w3), .A(w7) );
	io_OR g_8 (.B(w2), .Z(w4), .A(w20) );
	io_OR3 g_9 (.Z(w6), .C(w8), .B(w14), .A(w16) );
	io_NAND g_10 (.A(w161), .B(w932), .Z(w3) );
	io_NOT g_11 (.A(w161), .nZ(w22) );
	io_NOT g_12 (.A(w932), .nZ(w21) );
	io_NAND8 g_13 (.Z(w14), .D(w22), .C(w21), .B(w20), .A(1'b1), .E(w2), .F(w18), .G(w17), .H(w32) );
	io_AND3 g_14 (.Z(w31), .C(w32), .B(w17), .A(w18) );
	io_NOR g_15 (.Z(w7), .B(w31), .A(w30) );
	io_NOR3 g_16 (.Z(w30), .C(w17), .B(w32), .A(w18) );
	io_DFFRPOS g_17 (.Q(w29), .nRES(1'b1), .D(w186), .C(w33) );
	io_DFFRPOS g_18 (.Q(w27), .nRES(1'b1), .D(w156), .C(w33) );
	io_NOT g_19 (.A(w221), .nZ(w26) );
	io_DFFRPOS g_20 (.Q(w59), .nRES(1'b1), .D(w108), .C(w33) );
	io_DFFRPOS g_21 (.Q(w58), .nRES(1'b1), .D(w337), .C(w33) );
	io_NOT g_22 (.A(w120), .nZ(w62) );
	io_MUX4BIT g_23 (.C(w8), .Z0(w32), .B0(w100), .A0(w102), .B1(w99), .A1(w66), .Z1(w17), .Z2(w2), .A2(w54), .B2(w35), .B3(w188), .A3(w57), .Z3(w9) );
	io_NOT g_24 (.A(w166), .nZ(w60) );
	io_NOT g_25 (.A(w134), .nZ(w64) );
	io_DFFRPOS g_26 (.Q(w67), .nRES(1'b1), .D(w143), .C(w33) );
	io_DFFSPOS g_27 (.C(w12), .D(w130), .nSET(w122), .Q(w131) );
	io_MUX4BIT g_28 (.C(w8), .Z0(w190), .B0(w163), .A0(w133), .B1(w131), .A1(w124), .Z1(w24), .Z2(w68), .A2(w126), .B2(w162), .B3(w132), .A3(w123), .Z3(w75) );
	io_DFFSPOS g_29 (.C(w12), .D(w138), .nSET(w122), .Q(w163) );
	io_DFFSPOS g_30 (.C(w12), .D(w165), .nSET(w122), .Q(w162) );
	io_OR g_31 (.B(w153), .Z(w145), .A(w72) );
	io_AND g_32 (.Z(w147), .B(w145), .A(w71) );
	io_OR g_33 (.B(w153), .Z(w931), .A(w25) );
	io_MUX4BIT g_34 (.C(w8), .Z0(w154), .B0(w151), .A0(w28), .B1(w242), .A1(w61), .Z1(w150), .Z2(w149), .A2(w63), .B2(w28), .B3(w61), .A3(w65), .Z3(w152) );
	io_AND g_35 (.Z(w151), .A(w23), .B(w931) );
	io_DFFRPOS g_36 (.Q(w82), .nRES(1'b1), .D(w156), .C(w142) );
	io_NOT g_37 (.A(w77), .nZ(w83) );
	io_DFFRPOS g_38 (.Q(w81), .nRES(1'b1), .D(w108), .C(w142) );
	io_DFFRPOS g_39 (.Q(w85), .nRES(1'b1), .D(w143), .C(w142) );
	io_DFFRPOS g_40 (.Q(w934), .nRES(1'b1), .D(w337), .C(w142) );
	io_NOT g_41 (.A(w249), .nZ(w84) );
	io_DFFRPOS g_42 (.nRES(w112), .D(1'b0), .C(w86) );
	io_MUX4BIT g_43 (.C(w8), .B0(1'b0), .A0(1'b0), .B1(w91), .A1(w105), .Z1(w259), .Z2(w246), .A2(w91), .B2(w90), .B3(w101), .A3(w90), .Z3(w88) );
	io_DFFRPOS g_44 (.nRES(w112), .D(1'b0), .C(w86) );
	io_MUX4BIT g_45 (.C(w8), .Z0(w161), .B0(w105), .A0(1'b0), .B1(w91), .A1(w106), .Z1(w932), .Z2(w20), .A2(w104), .B2(w90), .B3(w101), .A3(w103), .Z3(w18) );
	io_NOR4 g_46 (.Z(w174), .D(w161), .C(w932), .B(w20), .A(w18) );
	io_DFFRPOS g_47 (.Q(w50), .nRES(w112), .D(w186), .C(w176) );
	io_DFFRPOS g_48 (.Q(w184), .nRES(w112), .D(w186), .C(w86) );
	io_DFFRPOS g_49 (.nRES(w112), .D(1'b0), .C(w176) );
	io_DFFRPOS g_50 (.nRES(w112), .D(1'b0), .C(w176) );
	io_DFFRPOS g_51 (.nRES(w112), .D(1'b0), .C(w137) );
	io_DFFRPOS g_52 (.nRES(w112), .D(1'b0), .C(w137) );
	io_DFFRPOS g_53 (.nRES(w112), .D(1'b0), .C(w137) );
	io_NAND4 g_54 (.B(w92), .C(w175), .A(w93), .D(w170) );
	io_NAND4 g_55 (.B(w94), .C(w93), .A(w92), .D(w170), .Z(w862) );
	io_NOT g_56 (.A(w2), .nZ(w168) );
	io_NAND4 g_57 (.B(w94), .C(w170), .A(w93), .D(w168) );
	io_NOT g_58 (.A(w170), .nZ(w95) );
	io_NAND4 g_59 (.B(w95), .C(w168), .A(w94), .D(w93) );
	io_NOT g_60 (.A(w175), .nZ(w94) );
	io_NAND4 g_61 (.B(w92), .C(w93), .A(w95), .D(w94) );
	io_NAND4 g_62 (.B(w95), .C(w175), .A(w92), .D(w93), .Z(w167) );
	io_NAND4 g_63 (.B(w95), .C(w175), .A(w93), .D(w168) );
	io_NOT g_64 (.A(w168), .nZ(w92) );
	io_NOT g_65 (.A(w96), .nZ(w46) );
	io_NOT g_66 (.A(w69), .nZ(w97) );
	io_AND3 g_67 (.Z(w192), .C(w237), .B(w236), .A(w881) );
	io_OR g_68 (.B(w291), .Z(w881), .A(w235) );
	io_NOT g_69 (.A(w268), .nZ(w235) );
	io_OR g_70 (.B(w268), .Z(w236), .A(w98) );
	io_OR g_71 (.B(w235), .Z(w234), .A(w98) );
	io_AND g_72 (.Z(w232), .B(w233), .A(w234) );
	io_OR g_73 (.B(w291), .Z(w233), .A(w268) );
	io_MUX4BIT g_74 (.C(w227), .Z0(w895), .B0(w198), .A0(w212), .B1(w197), .A1(w211), .Z1(w231), .Z2(w238), .A2(w210), .B2(w195), .B3(w191), .A3(w209), .Z3(w888) );
	io_NOT g_75 (.A(w816), .nZ(w933) );
	io_MUX4BIT g_76 (.C(w754), .Z0(w156), .B0(w198), .A0(w229), .B1(w197), .A1(w280), .Z1(w108), .Z2(w337), .A2(w228), .B2(w195), .B3(w191), .A3(w226), .Z3(w143) );
	io_MUX4BIT g_77 (.C(w53), .Z0(w213), .B0(w229), .A0(w904), .B1(w280), .A1(w903), .Z1(w196), .Z2(w194), .A2(w930), .B2(w228), .B3(w226), .A3(w225), .Z3(w193) );
	io_CNT_BIT g_78 (.nQ(w889), .C(w115), .RES(1'b1), .D(1'b1), .nLD(w119), .CI(w218) );
	io_NOR4 g_79 (.Z(w395), .D(w889), .C(w912), .B(w890), .A(w891) );
	io_CNT_BIT g_80 (.nQ(w890), .C(w115), .RES(1'b1), .D(1'b0), .nLD(w119), .CO(w892), .CI(w219) );
	io_CNT_BIT g_81 (.Q(w878), .nQ(w912), .C(w115), .RES(1'b1), .D(1'b0), .nLD(w119), .CO(w218), .CI(w892) );
	io_DFFRPOS g_82 (.Q(w134), .nRES(w112), .D(w143), .C(w855) );
	io_DFFRPOS g_83 (.Q(w126), .nRES(1'b1), .D(w130), .C(w142) );
	io_DFFRPOS g_84 (.Q(w123), .nRES(1'b1), .D(w165), .C(w142) );
	io_DFFRPOS g_85 (.Q(w124), .nRES(1'b1), .D(w165), .C(w33) );
	io_NOT g_86 (.A(w241), .nZ(w146) );
	io_DFFRPOS g_87 (.Q(w254), .nRES(1'b1), .D(w138), .C(w142) );
	io_MUX4BIT g_88 (.C(w8), .Z0(w798), .B0(w63), .A0(w254), .B1(w65), .A1(w70), .Z1(w762), .Z2(w243), .A2(w71), .B2(w147), .B3(w73), .A3(w73), .Z3(w244) );
	io_MUX8TO1 g_89 (.S0(w250), .S2(w247), .S1(w251), .G(w252), .H(w253), .F(w134), .E(w249), .Z(w894), .C(w152), .D(w307), .B(w107), .A(w893) );
	io_MUX8TO1 g_90 (.S0(w250), .S2(w247), .S1(w251), .G(w255), .H(w248), .F(w221), .E(w77), .Z(w896), .C(w154), .D(w314), .B(w76), .A(w897) );
	io_MUX8TO1 g_91 (.S0(w250), .S2(w247), .S1(w251), .G(w478), .H(w651), .F(w166), .E(w139), .Z(w905), .C(w150), .D(w257), .B(w258), .A(w790) );
	io_DFFSPOS g_92 (.C(w367), .D(w71), .nSET(w276), .nQ(w260), .Q(w557) );
	io_DFFRPOS g_93 (.Q(w906), .nRES(w907), .D(w260), .C(w437) );
	io_MUX8TO1 g_94 (.S0(w250), .S2(w247), .S1(w251), .G(w927), .H(w265), .F(w677), .E(w270), .Z(w901), .C(w880), .D(w262), .B(w269), .A(w264) );
	io_DFFRPOS g_95 (.Q(w265), .nRES(w112), .D(w156), .C(w86) );
	io_NOR3 g_96 (.Z(w53), .C(w268), .B(w266), .A(w267) );
	io_AND g_97 (.Z(w272), .B(1'b1), .A(w557) );
	io_DFFRPOS g_98 (.Q(w841), .nRES(w907), .D(1'b1), .C(w437) );
	io_DFFRPOS g_99 (.Q(w264), .nRES(1'b1), .D(w922), .C(w437) );
	io_DFFRPOS g_100 (.Q(w825), .nRES(1'b1), .D(w910), .C(w437) );
	io_NOT g_101 (.A(w275), .nZ(w182) );
	io_SIPO_4BIT g_102 (.i1(w356), .D(w272), .i9(w276), .o12(w923), .o13(w274), .o26(w852), .Q3(w911) );
	io_SIPO_4BIT g_103 (.i1(w356), .i2(w911), .i9(w276), .o12(w916), .o13(w918), .o26(w854), .o27(w750) );
	io_AND g_104 (.Z(w907), .B(w861), .A(w171) );
	io_DFFRPOS g_105 (.Q(w921), .nRES(1'b1), .D(w917), .C(w437) );
	io_DFFRPOS g_106 (.Q(w840), .nRES(1'b1), .D(w919), .C(w437) );
	io_NOT g_107 (.A(w32), .nZ(w857) );
	io_OR g_108 (.B(w268), .Z(w277), .A(w266) );
	io_NOR g_109 (.Z(w47), .B(w46), .A(w189) );
	io_NOR g_110 (.Z(w48), .B(w49), .A(w47) );
	io_NAND g_111 (.B(w240), .A(w53), .Z(w237) );
	io_NOR g_112 (.Z(w40), .B(w8), .A(w48) );
	io_DFFSPOS g_113 (.C(w230), .D(w52), .nSET(w50), .Q(w45) );
	io_AND g_114 (.Z(w43), .B(w50), .A(w45) );
	io_NOT g_115 (.A(w51), .nZ(w44) );
	io_NOR g_116 (.Z(w239), .B(w189), .A(w44) );
	io_NOT g_117 (.A(w50), .nZ(w42) );
	io_AND g_118 (.Z(w13), .B(w42), .A(w933) );
	io_OR g_119 (.B(w41), .Z(w15), .A(w43) );
	io_OR g_120 (.B(w42), .Z(w41), .A(w29) );
	io_NOT g_121 (.A(w8), .nZ(w38) );
	io_NOR g_122 (.Z(w39), .B(w56), .A(w38) );
	io_NOR g_123 (.Z(w245), .B(w40), .A(w39) );
	io_BUF g_124 (.Z(w240), .A(w8) );
	io_AND g_125 (.Z(w227), .B(w36), .A(w240) );
	io_NOT g_126 (.A(w188), .nZ(w36) );
	io_MUX4BIT g_127 (.C(w8), .Z0(w222), .B0(w100), .A0(w101), .B1(w99), .A1(w100), .Z1(w55), .Z2(w223), .A2(w99), .B2(w35), .B3(w188), .A3(w35), .Z3(w224) );
	io_AND3 g_128 (.Z(w37), .C(1'b1), .B(w119), .A(1'b1) );
	io_CNT_BIT g_129 (.nQ(w109), .C(w115), .RES(1'b1), .D(w121), .nLD(w119), .CO(w110), .CI(w37) );
	io_CNT_BIT g_130 (.nQ(w113), .C(w115), .RES(1'b1), .D(1'b0), .nLD(w119), .CO(w111), .CI(w110) );
	io_AND g_131 (.Z(w112), .B(w8), .A(w127) );
	io_NOR4 g_132 (.Z(w524), .D(w113), .C(w109), .B(w117), .A(w116) );
	io_CNT_BIT g_133 (.nQ(w116), .C(w115), .RES(1'b1), .D(1'b1), .nLD(w119), .CO(w118), .CI(w111) );
	io_CNT_BIT g_134 (.nQ(w117), .C(w115), .RES(1'b1), .D(1'b1), .nLD(w119), .CI(w118) );
	io_BUF g_135 (.Z(w128), .A(w129) );
	io_BUF g_136 (.Z(w122), .A(w127) );
	io_NOR g_137 (.Z(w49), .B(w70), .A(w97) );
	io_NOT g_138 (.A(w819), .nZ(w164) );
	io_DFFSPOS g_139 (.C(w12), .D(w337), .nSET(w122), .Q(w125) );
	io_DFFSPOS g_140 (.C(w12), .D(w108), .nSET(w122), .Q(w136) );
	io_MUX4BIT g_141 (.C(w8), .Z0(w96), .B0(w135), .A0(w146), .B1(w136), .A1(w180), .Z1(w25), .Z2(w69), .A2(w164), .B2(w125), .B3(w144), .A3(w148), .Z3(w72) );
	io_DFFSPOS g_142 (.C(w12), .D(w143), .nSET(w122), .Q(w144) );
	io_DFFSPOS g_143 (.C(w12), .D(w156), .nSET(w122), .Q(w135) );
	io_BUF g_144 (.Z(w251), .A(w129) );
	io_DFFRPOS g_145 (.Q(w249), .nRES(w112), .D(w143), .C(w140) );
	io_DFFRPOS g_146 (.Q(w77), .nRES(w112), .D(w156), .C(w140) );
	io_MUX8TO1 g_147 (.SO(w250), .S1(w251), .S2(w247), .G(w352), .H(w159), .F(w120), .E(w141), .Z(w158), .C(w149), .D(w157), .B(w160), .A(w256) );
	io_NOT g_148 (.A(w139), .nZ(w80) );
	io_NOT g_149 (.A(w141), .nZ(w79) );
	io_DFFRPOS g_150 (.Q(w139), .nRES(w112), .D(w108), .C(w140) );
	io_DFFRPOS g_151 (.Q(w789), .nRES(w112), .D(w138), .C(w137) );
	io_DFFRPOS g_152 (.Q(w261), .nRES(w112), .D(w186), .C(w137) );
	io_DFFRPOS g_153 (.Q(w141), .nRES(w112), .D(w337), .C(w140) );
	io_DFFRPOS g_154 (.nRES(w112), .D(1'b0), .C(w86) );
	io_DFFRPOS g_155 (.Q(w269), .nRES(w112), .D(w156), .C(w137) );
	io_DFFRPOS g_156 (.Q(w270), .nRES(w112), .D(w156), .C(w176) );
	io_OR g_157 (.A(w178), .Z(w180), .B(w179) );
	io_NOT g_158 (.A(w263), .nZ(w179) );
	io_DFFRPOS g_159 (.Q(w271), .nRES(w112), .D(w165), .C(w86) );
	io_DFFRPOS g_160 (.Q(w275), .nRES(w112), .D(w165), .C(w140) );
	io_OR g_161 (.B(w276), .Z(w148), .A(w182) );
	io_BUF g_162 (.Z(w247), .A(w181) );
	io_BUF g_163 (.Z(w183), .A(w181) );
	io_DFFRPOS g_164 (.nRES(w112), .D(1'b0), .C(w176) );
	io_DFFRPOS g_165 (.Q(w178), .nRES(w112), .D(w165), .C(w176) );
	io_DFFRPOS g_166 (.Q(w276), .nRES(w112), .D(w165), .C(w137) );
	io_AND g_167 (.Z(w181), .B(w17), .A(w8) );
	io_NOT g_168 (.A(w17), .nZ(w170) );
	io_NAND g_169 (.A(w8), .B(w174), .Z(w172) );
	io_AND g_170 (.Z(w267), .B(w173), .A(w172) );
	io_NOT g_171 (.A(w9), .nZ(w175) );
	io_NAND4 g_172 (.B(w175), .C(w170), .A(w168), .D(w93), .Z(w171) );
	io_NOR3 g_173 (.Z(w93), .C(w172), .B(w277), .A(w169) );
	io_NOT g_174 (.A(w32), .nZ(w169) );
	io_AND g_175 (.Z(w52), .B(w590), .A(w882) );
	io_NOT g_176 (.A(w883), .nZ(w882) );
	io_DFFRPOS g_177 (.Q(w883), .nRES(w50), .D(w884), .C(w729) );
	io_AON22 g_178 (.Z(w884), .B2(w733), .A2(w730), .B1(w885), .A1(w876) );
	io_DFFRPOS g_179 (.Q(w885), .nRES(w50), .D(w886), .C(w729) );
	io_NOT g_180 (.A(w730), .Z(w733) );
	io_AON22 g_181 (.Z(w886), .B2(w733), .A2(w730), .B1(w887), .A1(w767) );
	io_DFFRPOS g_182 (.Q(w887), .nRES(w50), .D(w877), .C(w729) );
	io_DFFRPOS g_183 (.Q(w221), .nRES(w112), .D(w156), .C(w855) );
	io_DFFRPOS g_184 (.Q(w166), .nRES(w112), .D(w108), .C(w855) );
	io_DFFRPOS g_185 (.Q(w120), .nRES(w112), .D(w337), .C(w855) );
	io_DFFRPOS g_186 (.Q(w51), .nRES(w112), .D(w138), .C(w855) );
	io_AND g_187 (.Z(w897), .B(w230), .A(w324) );
	io_CNT_BIT g_188 (.nQ(w891), .C(w115), .RES(1'b1), .D(1'b1), .nLD(w119), .CO(w219), .CI(w879) );
	io_DFFRPOS g_189 (.Q(w816), .nRES(w112), .D(w186), .C(w855) );
	io_DFFRPOS g_190 (.Q(w241), .nRES(w112), .D(w130), .C(w855) );
	io_DFFRPOS g_191 (.Q(w133), .nRES(1'b1), .D(w130), .C(w33) );
	io_DFFRPOS g_192 (.Q(w824), .nRES(1'b1), .D(w138), .C(w33) );
	io_DFFRPOS g_193 (.Q(w819), .nRES(w112), .D(w130), .C(w140) );
	io_DFFRPOS g_194 (.Q(w815), .nRES(w112), .D(w186), .C(w140) );
	io_DFFRPOS g_195 (.Q(w805), .nRES(w112), .D(w138), .C(w140) );
	io_AND g_196 (.Z(w893), .B(w367), .A(w324) );
	io_DFFRPOS g_197 (.Q(w869), .nRES(1'b1), .D(w186), .C(w142) );
	io_AND g_198 (.Z(w873), .B(w32), .A(w8) );
	io_MUX4BIT g_199 (.C(w53), .Z0(w278), .B0(w895), .A0(w904), .B1(w231), .A1(w903), .Z1(w279), .Z2(w281), .A2(w930), .B2(w238), .B3(w888), .A3(w225), .Z3(w282) );
	io_DFFRPOS g_200 (.Q(w263), .nRES(w112), .D(w165), .C(w855) );
	io_MUX4BIT g_201 (.C(w873), .Z0(w904), .B0(w896), .A0(w901), .B1(w905), .A1(w899), .Z1(w903), .Z2(w930), .A2(w829), .B2(w158), .B3(w894), .A3(w671), .Z3(w225) );
	io_DFFRPOS g_202 (.Q(w898), .nRES(1'b1), .D(w902), .C(w714) );
	io_NOR6 g_203 (.Z(w56), .F(w796), .E(w239), .D(w870), .C(w909), .B(w908), .A(w872) );
	io_MUX8TO1 g_204 (.S0(w250), .S2(w247), .S1(w251), .G(w860), .H(w868), .F(w749), .E(w900), .Z(w899), .C(w871), .D(w898), .B(w906), .A(w921) );
	io_AND g_205 (.Z(w909), .B(w831), .A(w265) );
	io_AND g_206 (.Z(w872), .B(w841), .A(w269) );
	io_AND g_207 (.Z(w908), .B(w830), .A(w270) );
	io_DFFRPOS g_208 (.Q(w672), .nSET(1'b1), .D(w929), .C(w714) );
	io_SIPO_4BIT g_209 (.i1(w363), .i2(w753), .i9(w178), .o12(w924), .o13(w926), .o26(w844), .o27(w867) );
	io_DFFRPOS g_210 (.Q(w927), .nRES(1'b1), .D(w866), .C(w638) );
	io_DFFRPOS g_211 (.Q(w900), .nRES(w920), .D(w928), .C(w714) );
	io_DFFSPOS g_212 (.C(w624), .D(w23), .nSET(w178), .nQ(w928), .Q(w846) );
	io_DFFRPOS g_213 (.Q(w847), .nRES(1'b1), .D(w273), .C(w437) );
	io_DFFRPOS g_214 (.Q(w865), .nRES(1'b1), .D(w864), .C(w437) );
	io_DFFRPOS g_215 (.Q(w830), .nRES(w920), .D(1'b1), .C(w714) );
	io_DFFRPOS g_216 (.Q(w262), .nRES(1'b1), .D(w863), .C(w714) );
	io_AND g_217 (.Z(w920), .B(w861), .A(w862) );
	io_NAND4 g_218 (.A(w858), .D(w739), .B(w915), .C(w447), .Z(w365) );
	io_AND g_219 (.Z(w859), .B(w739), .A(w447) );
	io_DFFRPOS g_220 (.nQ(w915), .nRES(w462), .D(w856), .C(w624) );
	io_NAND g_221 (.A(w874), .B(w914), .Z(w856) );
	io_OR g_222 (.A(w915), .Z(w914), .B(w702) );
	io_OR g_223 (.A(w701), .Z(w874), .B(w702) );
	io_NOR3 g_224 (.Z(w702), .C(w915), .B(w846), .A(w913) );
	io_NOT g_225 (.A(w859), .nZ(w913) );
	io_NOT g_226 (.A(w846), .nZ(w858) );
	io_NOT g_227 (.A(w857), .nZ(w851) );
	io_NOT g_228 (.A(w590), .nZ(w730) );
	io_DFFRPOS g_229 (.Q(w779), .nRES(w50), .D(w780), .C(w729) );
	io_AON22 g_230 (.Z(w780), .B2(w733), .A2(w730), .B1(w781), .A1(w770) );
	io_DFFRPOS g_231 (.Q(w781), .nRES(w50), .D(w778), .C(w729) );
	io_AON22 g_232 (.Z(w877), .B2(w733), .A2(w772), .B1(w779), .A1(w730) );
	io_AON22 g_233 (.Z(w778), .B2(w733), .A2(w730), .B1(w777), .A1(w774) );
	io_DFFRPOS g_234 (.Q(w777), .nRES(w50), .D(w776), .C(w729) );
	io_AON22 g_235 (.Z(w776), .B2(w775), .A2(w730), .B1(w733), .A1(w759) );
	io_DFFRPOS g_236 (.Q(w775), .nRES(w50), .D(w757), .C(w729) );
	io_BUF g_237 (.Z(w610), .A(w127) );
	io_TFF g_238 (.Q(w616), .T(w610), .C(w771) );
	io_TFF g_239 (.Q(w761), .T(w610), .C(w760) );
	io_TFF g_240 (.Q(w724), .T(w610), .C(w761) );
	io_DFFSPOS g_241 (.C(w413), .D(w615), .nSET(w261), .Q(w763) );
	io_AND3 g_242 (.Z(w879), .C(1'b1), .B(w119), .A(w391) );
	io_TFF g_243 (.Q(w771), .T(w610), .C(w764) );
	io_TFF g_244 (.Q(w764), .T(w610), .C(w724) );
	io_MUX g_245 (.C(w324), .Z(w769), .A(w121), .B(w878) );
	io_SLATCH g_246 (.nQ(w770), .C(w674), .Q(w880), .D(w156) );
	io_AND g_247 (.Z(w765), .B(w261), .A(w763) );
	io_MUX g_248 (.C(w324), .Z(w760), .A(w878), .B(w115) );
	io_SLATCH g_249 (.nQ(w876), .C(w674), .Q(w673), .D(w143) );
	io_SLATCH g_250 (.nQ(w772), .C(w674), .Q(w871), .D(w108) );
	io_SLATCH g_251 (.nQ(w773), .C(w674), .Q(w766), .D(w130) );
	io_SLATCH g_252 (.nQ(w774), .C(w674), .Q(w823), .D(w186) );
	io_MUX4BIT g_253 (.C(w873), .Z0(w755), .BO(w809), .A0(w811), .B1(w768), .A1(w820), .Z1(w758), .Z2(w821), .A2(w822), .B2(w808), .B3(w814), .A3(w807), .Z3(w727) );
	io_OR g_254 (.A(w96), .Z(w806), .B(w153) );
	io_AND g_255 (.Z(w804), .B(w189), .A(w806) );
	io_MUX4BIT g_256 (.C(w8), .Z0(w936), .B0(w804), .A0(w824), .B1(w803), .A1(w189), .Z1(w802), .Z2(w797), .A2(w23), .B2(1'b0), .B3(1'b1), .A3(w242), .Z3(w795) );
	io_MUX8TO1 g_257 (.S0(w799), .S2(w183), .S1(w128), .G(w679), .H(w736), .F(w263), .E(w275), .Z(w808), .C(w797), .D(w318), .B(w243), .A(w347) );
	io_OR g_258 (.B(w69), .Z(w787), .A(w153) );
	io_AND g_259 (.Z(w803), .B(w70), .A(w787) );
	io_NOT g_260 (.A(w815), .nZ(w785) );
	io_DFFRPOS g_261 (.Q(w792), .nRES(w112), .D(w186), .C(w431) );
	io_BUF g_262 (.Z(w861), .A(w127) );
	io_NOT g_263 (.A(w805), .nZ(w788) );
	io_NOR g_264 (.Z(w870), .B(w788), .A(w70) );
	io_AND g_265 (.Z(w155), .B(w785), .A(w786) );
	io_AND g_266 (.Z(w790), .B(w324), .A(w624) );
	io_NOT g_267 (.A(w261), .nZ(w786) );
	io_AND g_268 (.Z(w784), .B(w869), .A(w786) );
	io_AND g_269 (.Z(w256), .B(w324), .A(w413) );
	io_OR g_270 (.B(w784), .Z(w74), .A(w765) );
	io_MUX8TO1 g_271 (.S0(w799), .S2(w183), .S1(w128), .G(w654), .H(w818), .F(w748), .E(w723), .Z(w820), .C(w766), .D(w837), .B(w817), .A(w840) );
	io_DFFRPOS g_272 (.Q(w868), .nRES(w838), .D(w678), .C(w638) );
	io_DFFRPOS g_273 (.Q(w817), .nRES(w112), .D(w130), .C(w137) );
	io_DFFRPOS g_274 (.Q(w837), .nRES(1'b1), .D(w839), .C(w714) );
	io_SIPO_4BIT g_275 (.i1(w380), .i2(w656), .i9(w271), .o12(w875), .o13(w836), .o26(w842), .o27(w668) );
	io_MUX8TO1 g_276 (.S0(w799), .S2(w183), .S1(w128), .G(w704), .H(w271), .F(w558), .E(w178), .Z(w822), .C(w835), .D(w718), .B(w276), .A(w865) );
	io_DFFRPOS g_277 (.Q(w723), .nRES(w112), .D(w130), .C(w176) );
	io_DFFRPOS g_278 (.Q(w860), .nRES(1'b1), .D(w849), .C(w638) );
	io_AND g_279 (.Z(w838), .B(w167), .A(w861) );
	io_DFFRPOS g_280 (.Q(w831), .nRES(w838), .D(1'b1), .C(w638) );
	io_DFFRPOS g_281 (.Q(w827), .nRES(1'b1), .D(w853), .C(w437) );
	io_NOR3 g_282 (.Z(w741), .C(w851), .B(w172), .A(w16) );
	io_NAND4 g_283 (.A(w741), .D(w740), .B(w743), .C(w742), .Z(w333) );
	io_NAND4 g_284 (.A(w742), .D(w744), .B(w741), .C(w745), .Z(w855) );
	io_NAND4 g_285 (.A(w741), .D(w746), .B(w743), .C(w740), .Z(w33) );
	io_NAND4 g_286 (.B(w743), .C(w742), .A(w741), .D(w745), .Z(w142) );
	io_NAND4 g_287 (.B(w744), .C(w746), .A(w741), .D(w745), .Z(w140) );
	io_NOT g_288 (.A(w240), .nZ(w754) );
	io_MUX4BIT g_289 (.C(w53), .Z0(w205), .B0(w289), .A0(w755), .B1(w288), .A1(w758), .Z1(w203), .Z2(w201), .A2(w821), .B2(w286), .B3(w283), .A3(w727), .Z3(w200) );
	io_MUX4BIT g_290 (.C(w227), .Z0(w728), .B0(w206), .A0(w217), .B1(w204), .A1(w216), .Z1(w756), .Z2(w725), .A2(w215), .B2(w202), .B3(w199), .A3(w214), .Z3(w726) );
	io_AON22 g_291 (.Z(w757), .B2(w733), .A2(w730), .B1(w732), .A1(w773) );
	io_MUX4BIT g_292 (.C(w754), .Z0(w138), .B0(w206), .A0(w289), .B1(w204), .A1(w288), .Z1(w130), .Z2(w165), .A2(w286), .B2(w202), .B3(w199), .A3(w283), .Z3(w186) );
	io_MUX4BIT g_293 (.C(w53), .Z0(w290), .B0(w728), .A0(w755), .B1(w756), .A1(w758), .Z1(w287), .Z2(w285), .A2(w821), .B2(w725), .B3(w726), .A3(w727), .Z3(w284) );
	io_MUX2BIT4TO1 g_294 (.i2(w771), .i3(w612), .o5(w413), .i8(w722), .i9(w616), .i12(w760), .i13(w724), .o15(w367), .i18(w771), .i19(w761), .i21(w817), .i23(w789) );
	io_MUX2BIT4TO1 g_295 (.i2(w771), .i3(w612), .o5(w230), .i8(w722), .i9(w616), .i12(w760), .i13(w724), .o15(w624), .i18(w771), .i19(w761), .i21(w723), .i23(w810) );
	io_MUX2BIT4TO1 g_296 (.i2(w771), .i3(w612), .o5(w346), .i8(w722), .i9(w616), .i12(w760), .i13(w724), .o15(w427), .i18(w771), .i19(w761), .i21(w818), .i23(w793) );
	io_SLATCH g_297 (.nQ(w721), .C(w674), .Q(w791), .D(w138) );
	io_MUX8TO1 g_298 (.S0(w799), .S2(w183), .S1(w128), .G(w353), .H(w731), .F(w241), .E(w819), .Z(w768), .C(w802), .D(w321), .B(w762), .A(w769) );
	io_MUX8TO1 g_299 (.S0(w799), .S2(w183), .S1(w128), .G(w792), .H(w720), .F(w816), .E(w815), .Z(w814), .C(w795), .D(w317), .B(w244), .A(w605) );
	io_NOT g_300 (.A(w735), .nZ(w794) );
	io_NOR g_301 (.Z(w796), .B(w321), .A(w794) );
	io_DFFRPOS g_302 (.Q(w735), .nRES(w112), .D(w138), .C(w431) );
	io_MUX8TO1 g_303 (.S0(w799), .S2(w183), .S1(w128), .G(w735), .H(w734), .F(w51), .E(w805), .Z(w809), .C(w936), .D(w369), .B(w798), .A(w153) );
	io_SLATCH g_304 (.nQ(w767), .C(w674), .Q(w813), .D(w337) );
	io_NOT g_305 (.A(w792), .nZ(w812) );
	io_AND g_306 (.Z(w316), .B(w783), .A(w812) );
	io_NOT g_307 (.A(w184), .nZ(w783) );
	io_AND g_308 (.Z(w782), .B(w783), .A(w351) );
	io_MUX8TO1 g_309 (.S0(w799), .S2(w183), .S1(w128), .G(w463), .H(w793), .F(w565), .E(w810), .Z(w811), .C(w791), .D(w715), .B(w789), .A(w825) );
	io_AND g_310 (.Z(w826), .B(w184), .A(w737) );
	io_OR g_311 (.B(w782), .Z(w315), .A(w826) );
	io_DFFRPOS g_312 (.Q(w793), .nRES(w112), .D(w138), .C(w86) );
	io_MUX8TO1 g_313 (.S0(w250), .S2(w247), .S1(w251), .G(w832), .H(w831), .F(w719), .E(w830), .Z(w829), .C(w813), .D(w828), .B(w841), .A(w827) );
	io_DFFRPOS g_314 (.Q(w818), .nRES(w112), .D(w130), .C(w86) );
	io_DFFRPOS g_315 (.Q(w828), .nRES(1'b1), .D(w843), .C(w714) );
	io_DFFRPOS g_316 (.Q(w832), .nRES(1'b1), .D(w848), .C(w638) );
	io_MUX8TO1 g_317 (.S0(w799), .S2(w183), .S1(w128), .G(w834), .H(w184), .F(w682), .E(w50), .Z(w807), .C(w823), .D(w833), .B(w261), .A(w847) );
	io_DFFRPOS g_318 (.Q(w833), .nRES(1'b1), .D(w752), .C(w714) );
	io_SLATCH g_319 (.nQ(w759), .C(w674), .Q(w835), .D(w165) );
	io_DFFRPOS g_320 (.Q(w834), .nRES(1'b1), .D(w845), .C(w638) );
	io_DFFRPOS g_321 (.Q(w810), .nRES(w112), .D(w138), .C(w176) );
	io_BUF g_322 (.Z(w250), .A(w850) );
	io_BUF g_323 (.Z(w799), .A(w850) );
	io_XNOR g_324 (.A(w9), .B(w8), .Z(w850) );
	io_NOT g_325 (.A(w2), .nZ(w713) );
	io_NOT g_326 (.A(w17), .nZ(w712) );
	io_NOT g_327 (.A(w17), .nZ(w743) );
	io_NOT g_328 (.A(w9), .nZ(w746) );
	io_NAND4 g_329 (.B(w746), .C(w740), .A(w744), .D(w741), .Z(w431) );
	io_NOT g_330 (.A(w2), .nZ(w745) );
	io_NAND4 g_331 (.B(w741), .C(w742), .A(w740), .D(w744), .Z(w570) );
	io_NOT g_332 (.A(w745), .nZ(w740) );
	io_NAND4 g_333 (.B(w746), .C(w741), .A(w745), .D(w743) );
	io_NOT g_334 (.A(w743), .nZ(w744) );
	io_NOR3 g_335 (.Z(w710), .C(w16), .B(w172), .A(w747) );
	io_NOT g_336 (.A(w746), .nZ(w742) );
	io_NOT g_337 (.A(w32), .nZ(w747) );
	io_AND g_338 (.Z(w208), .B(w240), .A(w192) );
	io_MUX g_339 (.C(w240), .Z(w207), .A(w609), .B(w193) );
	io_DFFRPOS g_340 (.Q(w609), .nRES(w127), .D(w199), .C(w608) );
	io_OR g_341 (.B(w9), .Z(w608), .A(w6) );
	io_OR g_342 (.A(w230), .Z(w729), .B(1'b0) );
	io_AON22 g_343 (.Z(w606), .B2(w733), .A2(w721), .B1(1'b0), .A1(w730) );
	io_DFFRPOS g_344 (.Q(w732), .nRES(w50), .D(w606), .C(w729) );
	io_TFF g_345 (.Q(w722), .T(w610), .C(w611) );
	io_TFF g_346 (.Q(w611), .T(w610), .C(w612) );
	io_TFF g_347 (.Q(w612), .T(w610), .C(w616) );
	io_NOT g_348 (.A(w590), .nZ(w614) );
	io_NOT g_349 (.A(w230), .nZ(w613) );
	io_NOT g_350 (.A(w680), .nZ(w620) );
	io_AND g_351 (.Z(w615), .B(w507), .A(w618) );
	io_NOT g_352 (.A(w619), .nZ(w618) );
	io_DFFRPOS g_353 (.Q(w619), .nRES(w261), .D(w621), .C(w602) );
	io_cell_47 g_354 (.i2(w613), .i3(1'b0), .i4(w614), .i11(w629), .i18(w534), .o20(w626), .o21(w622) );
	io_DFFRPOS g_355 (.Q(w628), .nRES(w261), .D(w627), .C(w602) );
	io_AON22 g_356 (.Z(w621), .B2(w625), .A2(w630), .B1(w628), .A1(w598) );
	io_AON22 g_357 (.Z(w627), .B2(w625), .A2(w598), .B1(w631), .A1(w632) );
	io_DFFRPOS g_358 (.Q(w631), .nRES(w261), .D(w641), .C(w602) );
	io_AON22 g_359 (.Z(w642), .B2(w625), .A2(w643), .B1(w634), .A1(w598) );
	io_DFFRPOS g_360 (.Q(w640), .nRES(w261), .D(w642), .C(w602) );
	io_AON22 g_361 (.Z(w641), .B1(w625), .A2(w598), .B2(w640), .A1(w639) );
	io_SLATCH g_362 (.nQ(w635), .C(w644), .Q(w720), .D(w186) );
	io_NOT g_363 (.A(w570), .nZ(w644) );
	io_SLATCH g_364 (.nQ(w646), .C(w644), .Q(w731), .D(w130) );
	io_SLATCH g_365 (.nQ(w645), .C(w644), .Q(w736), .D(w165) );
	io_SLATCH g_366 (.nQ(w639), .C(w644), .Q(w651), .D(w336) );
	io_SLATCH g_367 (.nQ(w643), .C(w644), .Q(w248), .D(w156) );
	io_SLATCH g_368 (.nQ(w630), .C(w644), .Q(w253), .D(w143) );
	io_SLATCH g_369 (.nQ(w632), .C(w644), .Q(w159), .D(w337) );
	io_SLATCH g_370 (.nQ(w650), .C(w644), .Q(w734), .D(w138) );
	io_DFFSPOS g_371 (.C(w346), .D(w652), .nSET(w184), .Q(w737) );
	io_AND g_372 (.Z(w652), .B(w388), .A(w687) );
	io_SLATCH g_373 (.nQ(w569), .C(w568), .Q(w748), .D(w130) );
	io_NOT g_374 (.A(w684), .nZ(w687) );
	io_SLATCH g_375 (.nQ(w681), .C(w568), .Q(w749), .D(w336) );
	io_BUF g_376 (.Z(w432), .A(w127) );
	io_DFFRPOS g_377 (.Q(w684), .nRES(w184), .D(w683), .C(w539) );
	io_SLATCH g_378 (.nQ(w935), .C(w568), .Q(w682), .D(w186) );
	io_DFFRPOS g_379 (.Q(w679), .nRES(w112), .D(w165), .C(w431) );
	io_NOT g_380 (.A(w679), .nZ(w675) );
	io_DFFSPOS g_381 (.C(w427), .D(w318), .nSET(w271), .nQ(w678), .Q(w680) );
	io_OR g_382 (.A(w675), .Z(w319), .B(w271) );
	io_SLATCH g_383 (.nQ(w690), .C(w568), .Q(w719), .D(w337) );
	io_SLATCH g_384 (.nQ(w561), .C(w568), .Q(w677), .D(w156) );
	io_SLATCH g_385 (.nQ(w676), .C(w568), .Q(w669), .D(w143) );
	io_NOT g_386 (.A(w667), .nZ(w568) );
	io_MUX8TO1 g_387 (.S0(w250), .S2(w247), .S1(w251), .G(w661), .H(w666), .F(w669), .E(w626), .Z(w671), .C(w673), .D(w672), .B(w567), .A(w670) );
	io_NOT g_388 (.A(w629), .nZ(w674) );
	io_DFFRPOS g_389 (.Q(w670), .nRES(1'b1), .D(w738), .C(w437) );
	io_DFFRPOS g_390 (.Q(w715), .nRES(1'b1), .D(w691), .C(w714) );
	io_DFFRPOS g_391 (.Q(w718), .nRES(1'b1), .D(w693), .C(w714) );
	io_SIPO_4BIT g_392 (.i1(w363), .i2(w695), .i9(w178), .o12(w694), .o13(w751), .o26(w692), .o27(w753) );
	io_BUF g_393 (.Z(w436), .A(w432) );
	io_AND g_394 (.Z(w695), .B(w846), .A(1'b1) );
	io_BUF g_395 (.Z(w462), .A(w432) );
	io_NAND4 g_396 (.B(w713), .C(w709), .A(w710), .D(w711), .Z(w667) );
	io_NAND4 g_397 (.B(w711), .C(w707), .A(w710), .D(w709), .Z(w86) );
	io_NOT g_398 (.A(w713), .nZ(w707) );
	io_NAND4 g_399 (.B(w710), .C(w711), .A(w712), .D(w707) );
	io_NAND4 g_400 (.B(w713), .C(w710), .A(w712), .D(w711), .Z(w137) );
	io_NOT g_401 (.A(w708), .nZ(w711) );
	io_NAND4 g_402 (.B(w713), .C(w708), .A(w712), .D(w710) );
	io_NAND4 g_403 (.B(w713), .C(w708), .A(w710), .D(w709), .Z(w176) );
	io_NAND4 g_404 (.B(w712), .C(w707), .A(w710), .D(w708), .Z(w629) );
	io_NAND4 g_405 (.B(w707), .C(w708), .A(w710), .D(w709) );
	io_NOT g_406 (.A(w712), .nZ(w709) );
	io_NOT g_407 (.A(w9), .nZ(w708) );
	io_DFFSPOS g_408 (.C(w363), .D(w364), .nSET(w436), .Q(w706) );
	io_OR g_409 (.B(w363), .Z(w714), .A(w706) );
	io_DFFSPOS g_410 (.C(w624), .D(w700), .nSET(w462), .nQ(w363), .Q(w701) );
	io_DFFRPOS g_411 (.nQ(w581), .Q(w575), .nRES(w589), .D(w585), .C(w230) );
	io_NAND6 g_412 (.C(w588), .D(w583), .B(w587), .E(w582), .A(1'b1), .F(w581), .Z(w590) );
	io_NAND3 g_413 (.A(w583), .B(w582), .C(w581), .Z(w573) );
	io_DFFRPOS g_414 (.nQ(w587), .Q(w572), .nRES(w589), .D(w578), .C(w230) );
	io_NAND4 g_415 (.B(w575), .C(w582), .A(w587), .D(w584), .Z(w571) );
	io_DFFRPOS g_416 (.nQ(w588), .Q(w584), .nRES(w589), .D(w579), .C(w230) );
	io_NAND4 g_417 (.B(w587), .C(w575), .A(w588), .D(w582), .Z(w591) );
	io_DFFRPOS g_418 (.nQ(w582), .Q(w576), .nRES(w589), .D(w580), .C(w230) );
	io_DFFSPOS g_419 (.C(w230), .D(w591), .nSET(w589), .Q(w596) );
	io_BUF g_420 (.Z(w589), .A(w432) );
	io_NOT g_421 (.A(w595), .nZ(w594) );
	io_NOR3 g_422 (.Z(w592), .C(w594), .B(w680), .A(w597) );
	io_OR g_423 (.A(w592), .Z(w600), .B(w597) );
	io_NAND g_424 (.A(w600), .B(w593), .Z(w599) );
	io_DFFRPOS g_425 (.nQ(w597), .nRES(w501), .D(w599), .C(w427) );
	io_DFFSRPOS g_426 (.C(w596), .D(1'b0), .nRES(w534), .nSET(w622), .Q(w623) );
	io_AND g_427 (.Z(w595), .B(w389), .A(w378) );
	io_NAND4 g_428 (.B(w597), .C(w378), .A(w620), .D(w389), .Z(w379) );
	io_DFFPOS g_429 (.Q(w583), .D(w623), .C(w624) );
	io_NOT g_430 (.A(w598), .nZ(w625) );
	io_BUF g_431 (.Z(w375), .A(w432) );
	io_BUF g_432 (.Z(w534), .A(w127) );
	io_OR g_433 (.B(1'b0), .Z(w602), .A(w413) );
	io_DFFRPOS g_434 (.Q(w634), .nRES(w261), .D(w633), .C(w602) );
	io_AON22 g_435 (.Z(w633), .B2(w625), .A2(w598), .B1(w636), .A1(w635) );
	io_DFFSPOS g_436 (.C(w380), .D(w299), .nSET(w375), .Q(w637) );
	io_OR g_437 (.A(w380), .Z(w638), .B(w637) );
	io_DFFRPOS g_438 (.Q(w636), .nRES(w261), .D(w686), .C(w602) );
	io_AON22 g_439 (.Z(w686), .B2(w625), .A2(w645), .B1(w647), .A1(w598) );
	io_AON22 g_440 (.Z(w648), .B2(w625), .A2(w650), .B1(1'b0), .A1(w598) );
	io_AON22 g_441 (.Z(w603), .B2(w625), .A2(w646), .B1(w649), .A1(w598) );
	io_DFFRPOS g_442 (.Q(w649), .nRES(w261), .D(w648), .C(w602) );
	io_DFFRPOS g_443 (.Q(w647), .nRES(w261), .D(w603), .C(w602) );
	io_NOT g_444 (.A(w388), .nZ(w549) );
	io_NOT g_445 (.A(w388), .nZ(w564) );
	io_DFFRPOS g_446 (.Q(w604), .nRES(w184), .D(w601), .C(w539) );
	io_AON22 g_447 (.Z(w601), .B2(w548), .A2(w681), .B1(w685), .A1(w549) );
	io_DFFRPOS g_448 (.Q(w685), .nRES(w184), .D(w566), .C(w539) );
	io_AON22 g_449 (.Z(w566), .B2(w548), .A2(w549), .B1(w559), .A1(w561) );
	io_AON22 g_450 (.Z(w562), .B2(w548), .A2(w935), .B1(w550), .A1(w549) );
	io_DFFRPOS g_451 (.Q(w559), .nRES(w184), .D(w562), .C(w539) );
	io_DFFRPOS g_452 (.Q(w560), .nRES(w184), .D(w689), .C(w539) );
	io_AON22 g_453 (.Z(w689), .B2(w548), .A2(w690), .B1(w604), .A1(w549) );
	io_AON22 g_454 (.Z(w683), .B2(w548), .A2(w549), .B1(w560), .A1(w676) );
	io_NOT g_455 (.A(w346), .nZ(w688) );
	io_cell_47 g_456 (.i2(w688), .i3(1'b0), .i4(w564), .i11(w667), .i18(w534), .o20(w666), .o21(w665) );
	io_DFFSRPOS g_457 (.C(w514), .D(1'b0), .nRES(w534), .nSET(w665), .Q(w556) );
	io_AND g_458 (.Z(w659), .B(1'b1), .A(w664) );
	io_DFFRPOS g_459 (.Q(w661), .nRES(1'b1), .D(w660), .C(w638) );
	io_SIPO_4BIT g_460 (.i1(w380), .i2(w659), .i9(w271), .o12(w657), .o13(w658), .o26(w662), .o27(w656) );
	io_DFFRPOS g_461 (.Q(w654), .nRES(1'b1), .D(w655), .C(w638) );
	io_DFFRPOS g_462 (.Q(w463), .nRES(1'b1), .D(w653), .C(w638) );
	io_DFFSPOS g_463 (.C(w624), .D(w452), .nSET(w462), .nQ(w457), .Q(w454) );
	io_DFFSPOS g_464 (.C(w624), .D(w460), .nSET(w462), .nQ(w446), .Q(w458) );
	io_NAND4 g_465 (.B(w446), .C(w457), .A(w363), .D(w456), .Z(w464) );
	io_DFFRPOS g_466 (.nQ(w739), .Q(w434), .nRES(w436), .D(w444), .C(w363) );
	io_DFFRPOS g_467 (.Q(w704), .nRES(1'b1), .D(w705), .C(w638) );
	io_DFFRPOS g_468 (.nQ(w455), .Q(w456), .nRES(w462), .D(w703), .C(w624) );
	io_NOR g_469 (.Z(w703), .B(w456), .A(w702) );
	io_NOT g_470 (.A(w702), .nZ(w453) );
	io_NAND6 g_471 (.C(w698), .D(w466), .B(w697), .E(w464), .A(1'b1), .F(w453), .Z(w700) );
	io_NAND g_472 (.A(w701), .B(w458), .Z(w466) );
	io_NAND g_473 (.A(w701), .B(w454), .Z(w698) );
	io_NAND g_474 (.A(w455), .B(w701), .Z(w697) );
	io_NAND3 g_475 (.A(w486), .B(w571), .C(w573), .Z(w578) );
	io_NAND4 g_476 (.B(w577), .C(w487), .A(w571), .D(w486), .Z(w585) );
	io_NAND g_477 (.A(w576), .B(w575), .Z(w487) );
	io_NAND g_478 (.A(w572), .B(w575), .Z(w577) );
	io_NAND g_479 (.A(w576), .B(w572), .Z(w486) );
	io_NAND3 g_480 (.A(w576), .B(w572), .C(w581), .Z(w489) );
	io_NAND g_481 (.A(w582), .B(w575), .Z(w488) );
	io_NAND3 g_482 (.A(w488), .B(w573), .C(w489), .Z(w580) );
	io_NAND4 g_483 (.B(w573), .C(w489), .A(w574), .D(w490), .Z(w579) );
	io_NAND3 g_484 (.A(w584), .B(w576), .C(w575), .Z(w490) );
	io_NAND3 g_485 (.A(w575), .B(w584), .C(w572), .Z(w574) );
	io_NAND4 g_486 (.B(w493), .C(w492), .A(w380), .D(w502), .Z(w520) );
	io_NOT g_487 (.A(w592), .nZ(w499) );
	io_NOR g_488 (.Z(w509), .B(w502), .A(w592) );
	io_DFFRPOS g_489 (.nQ(w508), .Q(w502), .nRES(w501), .D(w509), .C(w427) );
	io_BUF g_490 (.Z(w501), .A(w432) );
	io_BUF g_491 (.Z(w411), .A(w432) );
	io_DFFSPOS g_492 (.C(w427), .D(w510), .nSET(w501), .nQ(w380), .Q(w515) );
	io_NAND g_493 (.A(w508), .B(w515), .Z(w516) );
	io_NAND6 g_494 (.C(1'b1), .D(w517), .B(w521), .E(w516), .A(w520), .F(w499), .Z(w510) );
	io_NAND g_495 (.A(w515), .B(w496), .Z(w521) );
	io_NAND g_496 (.A(w515), .B(w491), .Z(w517) );
	io_OR g_497 (.A(w515), .Z(w593), .B(w592) );
	io_DFFSPOS g_498 (.C(w413), .D(w506), .nSET(w411), .Q(w512) );
	io_NOT g_499 (.A(w507), .nZ(w598) );
	io_NOT g_500 (.A(w507), .nZ(w513) );
	io_BUF g_501 (.Z(w402), .A(w432) );
	io_DFFSPOS g_502 (.C(w346), .D(w511), .nSET(w402), .Q(w514) );
	io_NAND4 g_503 (.B(w387), .C(w384), .A(w394), .D(w383), .Z(w511) );
	io_DFFSRPOS g_504 (.C(w512), .D(1'b0), .nRES(w534), .nSET(w527), .Q(w518) );
	io_cell_47 g_505 (.i2(w535), .i3(1'b0), .i4(w513), .i11(w570), .i18(w534), .o20(w567), .o21(w527) );
	io_NOT g_506 (.A(w413), .nZ(w535) );
	io_DFFPOS g_507 (.Q(w528), .D(w556), .C(w427) );
	io_AND g_508 (.Z(w605), .B(w427), .A(w324) );
	io_DFFRPOS g_509 (.Q(w529), .nRES(w184), .D(w530), .C(w539) );
	io_BUF g_510 (.Z(w366), .A(w432) );
	io_AON22 g_511 (.Z(w530), .B2(w537), .A2(w569), .B1(w548), .A1(w549) );
	io_NOT g_512 (.A(w549), .nZ(w548) );
	io_DFFRPOS g_513 (.Q(w537), .nRES(w184), .D(w540), .C(w539) );
	io_AON22 g_514 (.Z(w540), .B2(w548), .A2(w549), .B1(1'b0), .A1(w541) );
	io_OR g_515 (.B(w346), .Z(w539), .A(1'b0) );
	io_AON22 g_516 (.Z(w547), .B2(w548), .A2(w483), .B1(w529), .A1(w549) );
	io_DFFRPOS g_517 (.Q(w550), .nRES(w184), .D(w547), .C(w539) );
	io_SLATCH g_518 (.nQ(w541), .C(w568), .Q(w565), .D(w138) );
	io_SLATCH g_519 (.nQ(w483), .C(w568), .Q(w558), .D(w165) );
	io_NOT g_520 (.A(w475), .nZ(w482) );
	io_NOR3 g_521 (.Z(w374), .C(w479), .B(w557), .A(w482) );
	io_DFFRPOS g_522 (.nQ(w479), .nRES(w366), .D(w480), .C(w367) );
	io_OR g_523 (.B(w481), .Z(w484), .A(w374) );
	io_NAND g_524 (.A(w485), .B(w484), .Z(w480) );
	io_OR g_525 (.B(w479), .Z(w485), .A(w374) );
	io_DFFRPOS g_526 (.Q(w478), .nRES(w112), .D(w336), .C(w431) );
	io_NOT g_527 (.A(w478), .nZ(w331) );
	io_DFFRPOS g_528 (.Q(w255), .nRES(w112), .D(w156), .C(w431) );
	io_NOT g_529 (.A(w557), .nZ(w555) );
	io_AND g_530 (.Z(w475), .B(w355), .A(w467) );
	io_NAND4 g_531 (.B(w479), .C(w467), .A(w555), .D(w355), .Z(w477) );
	io_NOT g_532 (.A(w255), .nZ(w313) );
	io_NAND4 g_533 (.B(w554), .C(w474), .A(w477), .D(w473), .Z(w433) );
	io_NAND g_534 (.A(w470), .B(w354), .Z(w474) );
	io_DFFRPOS g_535 (.nQ(w467), .Q(w470), .nRES(w358), .D(w476), .C(w356) );
	io_NAND4 g_536 (.B(w554), .C(w473), .A(w477), .D(w357), .Z(w476) );
	io_NAND3 g_537 (.A(w471), .B(w467), .C(w354), .Z(w473) );
	io_DFFRPOS g_538 (.nQ(w552), .Q(w471), .nRES(w358), .D(w430), .C(w356) );
	io_NAND4 g_539 (.B(w554), .C(w472), .A(w477), .D(w357), .Z(w430) );
	io_NAND3 g_540 (.A(w470), .B(w471), .C(w354), .Z(w472) );
	io_NAND4 g_541 (.B(w552), .C(w467), .A(w551), .D(w354), .Z(w554) );
	io_NAND4 g_542 (.B(w552), .C(w467), .A(w553), .D(w354), .Z(w357) );
	io_DFFRPOS g_543 (.nQ(w553), .Q(w551), .nRES(w358), .D(w468), .C(w356) );
	io_NAND4 g_544 (.B(w461), .C(w469), .A(w477), .D(w357), .Z(w468) );
	io_NAND3 g_545 (.A(w354), .B(w551), .C(w471), .Z(w469) );
	io_NAND3 g_546 (.A(w470), .B(w551), .C(w354), .Z(w461) );
	io_NAND4 g_547 (.A(w459), .D(w451), .B(w453), .C(w449), .Z(w460) );
	io_NAND g_548 (.A(w454), .B(w458), .Z(w459) );
	io_NAND g_549 (.A(w455), .B(w458), .Z(w451) );
	io_NAND3 g_550 (.A(w456), .B(w457), .C(w446), .Z(w449) );
	io_NAND g_551 (.A(w456), .B(w457), .Z(w450) );
	io_NAND g_552 (.A(w455), .B(w454), .Z(w448) );
	io_NAND3 g_553 (.A(w450), .B(w448), .C(w453), .Z(w452) );
	io_NAND4 g_554 (.B(w447), .C(w360), .A(w434), .D(w441), .Z(w364) );
	io_NAND4 g_555 (.B(w447), .C(w361), .A(w434), .D(w441), .Z(w443) );
	io_NAND3 g_556 (.A(w434), .B(w435), .C(w447), .Z(w439) );
	io_DFFRPOS g_557 (.nQ(w447), .Q(w429), .nRES(w436), .D(w445), .C(w363) );
	io_NAND4 g_558 (.B(w443), .C(w439), .A(w364), .D(w365), .Z(w445) );
	io_DFFRPOS g_559 (.nQ(w441), .Q(w435), .nRES(w436), .D(w442), .C(w363) );
	io_NAND4 g_560 (.B(w443), .C(w440), .A(w364), .D(w365), .Z(w442) );
	io_NAND4 g_561 (.B(w365), .C(w438), .A(w443), .D(w439), .Z(w444) );
	io_NAND3 g_562 (.A(w434), .B(w429), .C(w435), .Z(w440) );
	io_NAND g_563 (.A(w429), .B(w434), .Z(w438) );
	io_NAND g_564 (.A(w508), .B(w496), .Z(w494) );
	io_NAND g_565 (.A(w508), .B(w491), .Z(w495) );
	io_NAND g_566 (.A(w491), .B(w496), .Z(w422) );
	io_NAND4 g_567 (.B(w494), .C(w422), .A(w499), .D(w423), .Z(w500) );
	io_NAND3 g_568 (.A(w495), .B(w499), .C(w498), .Z(w497) );
	io_NAND g_569 (.A(w502), .B(w492), .Z(w498) );
	io_NAND3 g_570 (.A(w493), .B(w502), .C(w492), .Z(w423) );
	io_DFFSPOS g_571 (.C(w427), .D(w497), .nSET(w501), .nQ(w492), .Q(w491) );
	io_DFFSPOS g_572 (.C(w427), .D(w500), .nSET(w501), .nQ(w493), .Q(w496) );
	io_NAND3 g_573 (.A(w504), .B(w419), .C(w416), .Z(w421) );
	io_NAND4 g_574 (.A(w503), .D(w410), .B(w296), .C(w419), .Z(w506) );
	io_NAND6 g_575 (.C(w504), .D(w410), .B(w503), .E(w416), .A(1'b1), .F(w419), .Z(w507) );
	io_DFFRPOS g_576 (.nQ(w503), .Q(w329), .nRES(w411), .D(w426), .C(w413) );
	io_DFFPOS g_577 (.Q(w504), .D(w518), .C(w367) );
	io_NAND g_578 (.A(w405), .B(w394), .Z(w409) );
	io_NAND g_579 (.A(w398), .B(w394), .Z(w519) );
	io_NAND4 g_580 (.A(w409), .D(w404), .B(w519), .C(w403), .Z(w408) );
	io_DFFRPOS g_581 (.nQ(w385), .Q(w394), .nRES(w402), .D(w408), .C(w346) );
	io_NAND4 g_582 (.B(w406), .C(w384), .A(w394), .D(w383), .Z(w404) );
	io_NAND3 g_583 (.A(w398), .B(w405), .C(w385), .Z(w399) );
	io_NAND3 g_584 (.A(w394), .B(w406), .C(w398), .Z(w407) );
	io_NAND3 g_585 (.A(w405), .B(w406), .C(w523), .Z(w525) );
	io_NAND4 g_586 (.B(w407), .C(w396), .A(w525), .D(w399), .Z(w523) );
	io_DFFRPOS g_587 (.nQ(w387), .Q(w406), .nRES(w402), .D(w523), .C(w346) );
	io_NAND3 g_588 (.A(w384), .B(w385), .C(w528), .Z(w396) );
	io_NAND6 g_589 (.C(w387), .D(w383), .B(1'b1), .E(w384), .A(w528), .F(w385), .Z(w388) );
	io_DFFRPOS g_590 (.nQ(w389), .Q(w372), .nRES(w375), .D(w532), .C(w380) );
	io_NAND g_591 (.A(w373), .B(w372), .Z(w533) );
	io_NAND4 g_592 (.B(w533), .C(w376), .A(w379), .D(w377), .Z(w532) );
	io_NAND4 g_593 (.B(w379), .C(w376), .A(w299), .D(w377), .Z(w531) );
	io_DFFRPOS g_594 (.nQ(w378), .Q(w373), .nRES(w375), .D(w531), .C(w380) );
	io_DFFPOS g_595 (.nQ(w300), .Q(w127), .D(w292), .C(w115) );
	io_NOT g_596 (.A(w374), .nZ(w339) );
	io_NOR g_597 (.Z(w542), .B(w342), .A(w374) );
	io_DFFRPOS g_598 (.nQ(w345), .Q(w342), .nRES(w366), .D(w542), .C(w367) );
	io_NAND4 g_599 (.B(w368), .C(w342), .A(w356), .D(w343), .Z(w348) );
	io_DFFRPOS g_600 (.Q(w369), .nRES(1'b1), .D(w138), .C(w333) );
	io_NAND g_601 (.A(w345), .B(w481), .Z(w543) );
	io_DFFRPOS g_602 (.Q(w252), .nRES(w112), .D(w143), .C(w431) );
	io_NAND g_603 (.A(w344), .B(w481), .Z(w544) );
	io_NAND6 g_604 (.C(w544), .D(w348), .B(w543), .E(w339), .A(w545), .F(1'b1), .Z(w546) );
	io_NAND g_605 (.A(w481), .B(w350), .Z(w545) );
	io_DFFSPOS g_606 (.C(w367), .D(w546), .nSET(w366), .nQ(w356), .Q(w481) );
	io_DFFRPOS g_607 (.Q(w351), .nRES(1'b1), .D(w186), .C(w333) );
	io_NOT g_608 (.A(w352), .nZ(w310) );
	io_DFFRPOS g_609 (.Q(w352), .nRES(w112), .D(w337), .C(w431) );
	io_DFFRPOS g_610 (.Q(w353), .nRES(w112), .D(w130), .C(w431) );
	io_NOT g_611 (.A(w353), .nZ(w322) );
	io_BUF g_612 (.Z(w358), .A(w432) );
	io_DFFRPOS g_613 (.nQ(w355), .Q(w354), .nRES(w358), .D(w433), .C(w356) );
	io_DFFSPOS g_614 (.C(w356), .D(w357), .nSET(w358), .Q(w359) );
	io_OR g_615 (.A(w359), .Z(w437), .B(w356) );
	io_DFFRPOS g_616 (.nQ(w360), .Q(w361), .nRES(w436), .D(w362), .C(w363) );
	io_NAND4 g_617 (.B(w365), .C(w334), .A(w364), .D(w335), .Z(w362) );
	io_NAND3 g_618 (.A(w434), .B(w435), .C(w361), .Z(w335) );
	io_NAND3 g_619 (.A(w429), .B(w361), .C(w434), .Z(w334) );
	io_OR g_620 (.A(w325), .Z(w16), .B(w266) );
	io_DFFRPOS g_621 (.nQ(w410), .Q(w412), .nRES(w411), .D(w415), .C(w413) );
	io_DFFRPOS g_622 (.nQ(w416), .Q(w296), .nRES(w411), .D(w414), .C(w413) );
	io_NAND g_623 (.A(w412), .B(w296), .Z(w295) );
	io_NAND4 g_624 (.B(w418), .C(w294), .A(w417), .D(w295), .Z(w414) );
	io_NAND3 g_625 (.A(w421), .B(w418), .C(w294), .Z(w415) );
	io_NAND g_626 (.A(w420), .B(w412), .Z(w418) );
	io_NAND g_627 (.A(w420), .B(w296), .Z(w417) );
	io_NAND4 g_628 (.B(w419), .C(w329), .A(w410), .D(w296), .Z(w294) );
	io_DFFRPOS g_629 (.nQ(w419), .Q(w420), .nRES(w411), .D(w425), .C(w413) );
	io_NAND3 g_630 (.A(w416), .B(w412), .C(w420), .Z(w424) );
	io_NAND g_631 (.A(w419), .B(w296), .Z(w428) );
	io_NAND3 g_632 (.A(w424), .B(w421), .C(w428), .Z(w425) );
	io_NAND3 g_633 (.A(w420), .B(w329), .C(w296), .Z(w297) );
	io_NAND4 g_634 (.B(w424), .C(w298), .A(w421), .D(w297), .Z(w426) );
	io_NAND3 g_635 (.A(w412), .B(w329), .C(w296), .Z(w298) );
	io_DFFRPOS g_636 (.nQ(w383), .Q(w405), .nRES(w402), .D(w401), .C(w346) );
	io_NAND g_637 (.A(w398), .B(w405), .Z(w403) );
	io_NAND3 g_638 (.A(w403), .B(w404), .C(w396), .Z(w401) );
	io_DFFRPOS g_639 (.nQ(w384), .Q(w398), .nRES(w402), .D(w397), .C(w346) );
	io_NAND3 g_640 (.A(w393), .B(w399), .C(w396), .Z(w397) );
	io_NAND g_641 (.A(w384), .B(w394), .Z(w393) );
	io_AND g_642 (.Z(w400), .B(w391), .A(w395) );
	io_NOR g_643 (.Z(w392), .B(w300), .A(w400) );
	io_BUF g_644 (.Z(w119), .A(w392) );
	io_AND g_645 (.Z(w391), .B(1'b1), .A(w524) );
	io_DFFRPOS g_646 (.nQ(w326), .Q(w390), .nRES(w375), .D(w381), .C(w380) );
	io_DFFRPOS g_647 (.nQ(w328), .Q(w327), .nRES(w375), .D(w382), .C(w380) );
	io_NAND3 g_648 (.A(w373), .B(w390), .C(w372), .Z(w301) );
	io_NAND4 g_649 (.B(w377), .C(w301), .A(w379), .D(w299), .Z(w381) );
	io_NAND4 g_650 (.B(w372), .C(w326), .A(w378), .D(w327), .Z(w377) );
	io_NAND4 g_651 (.B(w299), .C(w302), .A(w379), .D(w303), .Z(w382) );
	io_NAND4 g_652 (.B(w378), .C(w326), .A(w372), .D(w328), .Z(w299) );
	io_NAND3 g_653 (.A(w378), .B(w390), .C(w372), .Z(w376) );
	io_NAND3 g_654 (.A(w372), .B(w327), .C(w390), .Z(w303) );
	io_NAND3 g_655 (.A(w373), .B(w327), .C(w372), .Z(w302) );
	io_NAND g_656 (.A(w344), .B(w350), .Z(w304) );
	io_NAND g_657 (.A(w350), .B(w345), .Z(w371) );
	io_NAND4 g_658 (.B(w371), .C(w304), .A(w339), .D(w305), .Z(w370) );
	io_DFFSPOS g_659 (.C(w367), .D(w370), .nSET(w366), .nQ(w368), .Q(w350) );
	io_NAND3 g_660 (.A(w343), .B(w342), .C(w368), .Z(w305) );
	io_DFFSPOS g_661 (.C(w367), .D(w340), .nSET(w366), .nQ(w343), .Q(w344) );
	io_NAND g_662 (.A(w342), .B(w343), .Z(w341) );
	io_NAND3 g_663 (.A(w338), .B(w339), .C(w341), .Z(w340) );
	io_NAND g_664 (.A(w345), .B(w344), .Z(w338) );
	io_MUX g_665 (.C(w324), .Z(w347), .A(w306), .B(w346) );
	io_NOT g_666 (.A(w293), .nZ(w121) );
	io_NOT g_667 (.A(w252), .nZ(w308) );
	io_DFFRPOS g_668 (.Q(w330), .nRES(1'b1), .D(w143), .C(w333) );
	io_DFFRPOS g_669 (.Q(w309), .nRES(1'b1), .D(w337), .C(w333) );
	io_DFFRPOS g_670 (.Q(w323), .nRES(1'b1), .D(w130), .C(w333) );
	io_DFFRPOS g_671 (.Q(w311), .nRES(1'b1), .D(w336), .C(w333) );
	io_DFFRPOS g_672 (.Q(w320), .nRES(1'b1), .D(w165), .C(w333) );
	io_DFFRPOS g_673 (.Q(w312), .nRES(1'b1), .D(w156), .C(w333) );
	io_DFFSPOS g_674 (.C(w12), .D(w186), .nSET(w122), .Q(w132) );
	io_RCDELAY g_675 (.A(w658), .Z(w655) );
	io_RCDELAY g_676 (.A(w692), .Z(w693) );
	io_RCDELAY g_677 (.A(w694), .Z(w691) );
	io_RCDELAY g_678 (.A(w657), .Z(w653) );
	io_RCDELAY g_679 (.A(w662), .Z(w705) );
	io_RCDELAY g_680 (.A(w750), .Z(w738) );
	io_RCDELAY g_681 (.A(w753), .Z(w752) );
	io_RCDELAY g_682 (.A(w844), .Z(w843) );
	io_RCDELAY g_683 (.A(w842), .Z(w848) );
	io_RCDELAY g_684 (.A(w751), .Z(w839) );
	io_RCDELAY g_685 (.A(w656), .Z(w845) );
	io_RCDELAY g_686 (.A(w836), .Z(w849) );
	io_RCDELAY g_687 (.A(w875), .Z(w866) );
	io_RCDELAY g_688 (.A(w852), .Z(w864) );
	io_RCDELAY g_689 (.A(w854), .Z(w853) );
	io_RCDELAY g_690 (.A(w274), .Z(w919) );
	io_RCDELAY g_691 (.A(w918), .Z(w917) );
	io_RCDELAY g_692 (.A(w916), .Z(w922) );
	io_RCDELAY g_693 (.A(w923), .Z(w910) );
	io_RCDELAY g_694 (.A(w924), .Z(w863) );
	io_RCDELAY g_695 (.A(w867), .Z(w929) );
	io_RCDELAY g_696 (.A(w911), .Z(w273) );
	io_RCDELAY g_697 (.A(w926), .Z(w902) );
	io_RCDELAY g_698 (.A(w668), .Z(w660) );
endmodule // IO

// Module Definitions [It is possible to wrap here on your primitives]

module io_AND (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // io_AND

module io_OR (  A, Z, B);

	input wire A;
	output wire Z;
	input wire B;

endmodule // io_OR

module io_NOR (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // io_NOR

module io_NOT (  A, nZ);

	input wire A;
	output wire nZ;

endmodule // io_NOT

module io_OR4 (  Z, D, C, B, A);

	output wire Z;
	input wire D;
	input wire C;
	input wire B;
	input wire A;

endmodule // io_OR4

module io_OR3 (  Z, C, B, A);

	output wire Z;
	input wire C;
	input wire B;
	input wire A;

endmodule // io_OR3

module io_NAND (  A, B, Z);

	input wire A;
	input wire B;
	output wire Z;

endmodule // io_NAND

module io_NAND8 (  Z, D, C, B, A, E, F, G, H);

	output wire Z;
	input wire D;
	input wire C;
	input wire B;
	input wire A;
	input wire E;
	input wire F;
	input wire G;
	input wire H;

endmodule // io_NAND8

module io_AND3 (  Z, C, B, A);

	output wire Z;
	input wire C;
	input wire B;
	input wire A;

endmodule // io_AND3

module io_NOR3 (  Z, C, B, A);

	output wire Z;
	input wire C;
	input wire B;
	input wire A;

endmodule // io_NOR3

module io_DFFRPOS (  nQ, Q, nRES, D, C);

	output wire nQ;
	output wire Q;
	input wire nRES;
	input wire D;
	input wire C;

endmodule // io_DFFRPOS

module io_MUX4BIT (  C, Z0, B0, A0, B1, A1, Z1, Z2, A2, B2, B3, A3, Z3);

	input wire C;
	output wire Z0;
	input wire B0;
	input wire A0;
	input wire B1;
	input wire A1;
	output wire Z1;
	output wire Z2;
	input wire A2;
	input wire B2;
	input wire B3;
	input wire A3;
	output wire Z3;

endmodule // io_MUX4BIT

module io_DFFSPOS (  C, D, nSET, nQ, Q);

	input wire C;
	input wire D;
	input wire nSET;
	output wire nQ;
	output wire Q;

endmodule // io_DFFSPOS

module io_NOR4 (  Z, D, C, B, A);

	output wire Z;
	input wire D;
	input wire C;
	input wire B;
	input wire A;

endmodule // io_NOR4

module io_NAND4 (  B, C, A, D, Z);

	input wire B;
	input wire C;
	input wire A;
	input wire D;
	output wire Z;

endmodule // io_NAND4

module io_CNT_BIT (  Q, nQ, C, RES, D, nLD, CO, CI);

	output wire Q;
	output wire nQ;
	input wire C;
	input wire RES;
	input wire D;
	input wire nLD;
	output wire CO;
	input wire CI;

endmodule // io_CNT_BIT

module io_MUX8TO1 (  S0, S2, S1, G, H, F, E, Z, C, D, B, A);

	input wire S0;
	input wire S2;
	input wire S1;
	input wire G;
	input wire H;
	input wire F;
	input wire E;
	output wire Z;
	input wire C;
	input wire D;
	input wire B;
	input wire A;

endmodule // io_MUX8TO1

module io_SIPO_4BIT (  i1, D, i9, o12, o13, o26, Q3);

	input wire i1;
	input wire D;
	input wire i9;
	output wire o12;
	output wire o13;
	output wire o26;
	output wire Q3;

endmodule // io_SIPO_4BIT

module io_BUF (  Z, A);

	output wire Z;
	input wire A;

endmodule // io_BUF

module io_AON22 (  Z, B2, A2, B1, A1);

	output wire Z;
	input wire B2;
	input wire A2;
	input wire B1;
	input wire A1;

endmodule // io_AON22

module io_NOR6 (  Z, F, E, D, C, B, A);

	output wire Z;
	input wire F;
	input wire E;
	input wire D;
	input wire C;
	input wire B;
	input wire A;

endmodule // io_NOR6

module io_TFF (  nQ, Q, T, C);

	output wire nQ;
	output wire Q;
	input wire T;
	input wire C;

endmodule // io_TFF

module io_MUX (  C, Z, A, B);

	input wire C;
	output wire Z;
	input wire A;
	input wire B;

endmodule // io_MUX

module io_SLATCH (  nQ, C, Q, D);

	output wire nQ;
	input wire C;
	output wire Q;
	input wire D;

endmodule // io_SLATCH

module io_MUX2BIT4TO1 (  i2, i3, o5, i8, i9, i12, i13, o15, i18, i19, i21, i23);

	input wire i2;
	input wire i3;
	output wire o5;
	input wire i8;
	input wire i9;
	input wire i12;
	input wire i13;
	output wire o15;
	input wire i18;
	input wire i19;
	input wire i21;
	input wire i23;

endmodule // io_MUX2BIT4TO1

module io_XNOR (  A, B, Z);

	input wire A;
	input wire B;
	output wire Z;

endmodule // io_XNOR

module io_cell_47 (  i2, i3, i4, i11, i18, o20, o21);

	input wire i2;
	input wire i3;
	input wire i4;
	input wire i11;
	input wire i18;
	output wire o20;
	output wire o21;

endmodule // io_cell_47

module io_NAND6 (  C, D, B, E, A, F, Z);

	input wire C;
	input wire D;
	input wire B;
	input wire E;
	input wire A;
	input wire F;
	output wire Z;

endmodule // io_NAND6

module io_NAND3 (  A, B, C, Z);

	input wire A;
	input wire B;
	input wire C;
	output wire Z;

endmodule // io_NAND3

module io_DFFSRPOS (  C, D, nRES, nQ, nSET, Q);

	input wire C;
	input wire D;
	input wire nRES;
	output wire nQ;
	input wire nSET;
	output wire Q;

endmodule // io_DFFSRPOS

module io_DFFPOS (  nQ, Q, D, C);

	output wire nQ;
	output wire Q;
	input wire D;
	input wire C;

endmodule // io_DFFPOS

module io_RCDELAY (  A, Z);

	input wire A;
	output wire Z;

endmodule // io_RCDELAY



// ERROR: floating wire w19
// ERROR: floating wire w34
// ERROR: floating wire w78
// ERROR: floating wire w87
// ERROR: floating wire w89
// ERROR: floating wire w114
// ERROR: floating wire w177
// ERROR: floating wire w185
// ERROR: floating wire w187
// ERROR: floating wire w220
// ERROR: floating wire w332
// ERROR: floating wire w336
// ERROR: floating wire w349
// ERROR: floating wire w386
// ERROR: floating wire w465
// ERROR: floating wire w505
// ERROR: floating wire w522
// ERROR: floating wire w526
// ERROR: floating wire w536
// ERROR: floating wire w538
// ERROR: floating wire w563
// ERROR: floating wire w586
// ERROR: floating wire w607
// ERROR: floating wire w617
// ERROR: floating wire w663
// ERROR: floating wire w664
// ERROR: floating wire w696
// ERROR: floating wire w699
// ERROR: floating wire w716
// ERROR: floating wire w717
// ERROR: floating wire w800
// ERROR: floating wire w801
// ERROR: floating wire w925
// WARNING: Cell io_DFFRPOS:g_17 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_18 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_20 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_21 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_26 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_27 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_29 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_30 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_36 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_38 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_39 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_40 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_42 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_42 port Q not connected.
// WARNING: Cell io_MUX4BIT:g_43 port Z0 not connected.
// WARNING: Cell io_DFFRPOS:g_44 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_44 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_47 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_48 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_49 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_49 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_50 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_50 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_51 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_51 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_52 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_52 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_53 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_53 port Q not connected.
// WARNING: Cell io_NAND4:g_54 port Z not connected.
// WARNING: Cell io_NAND4:g_57 port Z not connected.
// WARNING: Cell io_NAND4:g_59 port Z not connected.
// WARNING: Cell io_NAND4:g_61 port Z not connected.
// WARNING: Cell io_NAND4:g_63 port Z not connected.
// WARNING: Cell io_CNT_BIT:g_78 port Q not connected.
// WARNING: Cell io_CNT_BIT:g_78 port CO not connected.
// WARNING: Cell io_CNT_BIT:g_80 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_82 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_83 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_84 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_85 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_87 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_93 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_95 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_98 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_99 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_100 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_105 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_106 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_113 port nQ not connected.
// WARNING: Cell io_CNT_BIT:g_129 port Q not connected.
// WARNING: Cell io_CNT_BIT:g_130 port Q not connected.
// WARNING: Cell io_CNT_BIT:g_133 port Q not connected.
// WARNING: Cell io_CNT_BIT:g_134 port Q not connected.
// WARNING: Cell io_CNT_BIT:g_134 port CO not connected.
// WARNING: Cell io_DFFSPOS:g_139 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_140 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_142 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_143 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_145 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_146 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_150 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_151 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_152 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_153 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_154 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_154 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_155 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_156 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_159 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_160 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_164 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_164 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_165 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_166 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_177 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_179 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_182 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_183 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_184 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_185 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_186 port nQ not connected.
// WARNING: Cell io_CNT_BIT:g_188 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_189 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_190 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_191 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_192 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_193 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_194 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_195 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_197 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_200 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_202 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_208 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_210 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_211 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_213 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_214 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_215 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_216 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_220 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_229 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_231 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_234 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_236 port nQ not connected.
// WARNING: Cell io_TFF:g_238 port nQ not connected.
// WARNING: Cell io_TFF:g_239 port nQ not connected.
// WARNING: Cell io_TFF:g_240 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_241 port nQ not connected.
// WARNING: Cell io_TFF:g_243 port nQ not connected.
// WARNING: Cell io_TFF:g_244 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_261 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_272 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_273 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_274 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_277 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_278 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_280 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_281 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_302 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_312 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_314 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_315 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_316 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_318 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_320 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_321 port nQ not connected.
// WARNING: Cell io_NAND4:g_333 port Z not connected.
// WARNING: Cell io_DFFRPOS:g_340 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_344 port nQ not connected.
// WARNING: Cell io_TFF:g_345 port nQ not connected.
// WARNING: Cell io_TFF:g_346 port nQ not connected.
// WARNING: Cell io_TFF:g_347 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_353 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_355 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_358 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_360 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_371 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_377 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_379 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_389 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_390 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_391 port nQ not connected.
// WARNING: Cell io_NAND4:g_399 port Z not connected.
// WARNING: Cell io_NAND4:g_402 port Z not connected.
// WARNING: Cell io_NAND4:g_405 port Z not connected.
// WARNING: Cell io_DFFSPOS:g_408 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_419 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_425 port Q not connected.
// WARNING: Cell io_DFFSRPOS:g_426 port nQ not connected.
// WARNING: Cell io_DFFPOS:g_429 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_434 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_436 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_438 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_442 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_443 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_446 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_448 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_451 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_452 port nQ not connected.
// WARNING: Cell io_DFFSRPOS:g_457 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_459 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_461 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_462 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_467 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_498 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_502 port nQ not connected.
// WARNING: Cell io_DFFSRPOS:g_504 port nQ not connected.
// WARNING: Cell io_DFFPOS:g_507 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_509 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_513 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_517 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_522 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_526 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_528 port nQ not connected.
// WARNING: Cell io_DFFPOS:g_577 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_600 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_602 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_607 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_609 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_610 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_614 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_668 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_669 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_670 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_671 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_672 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_673 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_674 port nQ not connected.
