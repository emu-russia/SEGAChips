module VDP (  CH0_EN, CH0VOL[0], CH0VOL[1], CH1_EN, CH1VOL[0], CH1VOL[1], CH2_EN, CH2VOL[0], CH2VOL[1], CH3_EN, CH3VOL[0], CH3VOL[1], PSGDAC0[0], PSGDAC0[1], PSGDAC0[2], PSGDAC0[3], PSGDAC0[4], PSGDAC0[5], PSGDAC0[6], PSGDAC0[7], PSGDAC1[0], PSGDAC1[1], PSGDAC1[2], PSGDAC1[3], PSGDAC1[4], PSGDAC1[5], PSGDAC1[6], PSGDAC1[7], PSGDAC2[0], PSGDAC2[1], PSGDAC2[2], PSGDAC2[3], PSGDAC2[4], PSGDAC2[5], PSGDAC2[6], PSGDAC2[7], PSGDAC3[0], PSGDAC3[1], PSGDAC3[2], PSGDAC3[3], PSGDAC3[4], PSGDAC3[5], PSGDAC3[6], PSGDAC3[7], CAi[22], CAo[22], CA[19], DTACK_OUT, Z80_INT, RA[7], RA[6], RA[5], RA[4], RA[2], RA[1], RA[0], nRAS0, RA[3], nCAS0, nOE0, nLWR, nUWR, DTACK_IN, RnW, nLDS, nUDS, nAS, nM1, nWR, nRD, nIORQ, nILP2, nILP1, nINTAK, nMREQ, nBG, BGACK_OUT, BGACK_IN, nBR, VSYNC, nCSYNC, nCSYNC_IN, nHSYNC, nHSYNC_IN, DB[15], DB[14], DB[13], DB[12], DB[11], DB[10], DB[9], DB[8], DB[7], DB[6], DB[5], DB[4], DB[3], DB[2], DB[1], DB[0], CA[0], CA[1], CA[2], CA[3], CA[4], CA[5], CA[6], CA[7], CA[8], CA[9], CA[10], CA[11], CA[12], CA[13], CA[14], CA[15], CA[16], CA[17], CA[18], CA[20], CA[21], R_DAC[0], R_DAC[1], R_DAC[2], R_DAC[3], R_DAC[4], R_DAC[5], R_DAC[6], R_DAC[7], R_DAC[8], G_DAC[0], G_DAC[1], G_DAC[2], G_DAC[3], G_DAC[4], G_DAC[5], G_DAC[6], G_DAC[7], G_DAC[8], R_DAC[9], R_DAC[10], R_DAC[11], R_DAC[12], R_DAC[13], R_DAC[14], R_DAC[15], R_DAC[16], B_DAC[0], B_DAC[1], B_DAC[2], B_DAC[3], B_DAC[4], B_DAC[5], B_DAC[6], B_DAC[7], B_DAC[8], G_DAC[9], G_DAC[10], G_DAC[11], G_DAC[12], G_DAC[13], G_DAC[14], G_DAC[15], G_DAC[16], B_DAC[9], B_DAC[10], B_DAC[11], B_DAC[12], B_DAC[13], B_DAC[14], B_DAC[15], B_DAC[16], nOE1, nWE0, nWE1, nCAS1, nRAS1, AD_RD_DIR, nYS, nSC, nSE0_1, ADo[7], ADo[6], ADo[5], ADo[4], ADo[3], ADo[2], ADo[1], ADo[0], RDo[6], RDo[5], RDo[4], RDo[3], RDo[2], RDo[1], RDo[0], RDi[6], RDi[7], RDi[4], RDi[5], RDi[2], RDi[3], RDi[0], RDi[1], ADi[6], ADi[7], ADi[4], ADi[5], ADi[2], ADi[3], ADi[0], ADi[1], RDo[7], SD[7], SD[6], SD[5], SD[4], SD[3], SD[2], SD[1], SD[0], CLK1, CLK0, EDCLKi, EDCLKo, MCLK, SUB_CLK, nRES_PAD, 68kCLKi, EDCLKd, CA_PAD_DIR, DB_PAD_DIR, SEL0_M3, nPAL, nHL, SPA/Bo, SPA/Bi);

	output wire CH0_EN;
	output wire CH0VOL[0];
	output wire CH0VOL[1];
	output wire CH1_EN;
	output wire CH1VOL[0];
	output wire CH1VOL[1];
	output wire CH2_EN;
	output wire CH2VOL[0];
	output wire CH2VOL[1];
	output wire CH3_EN;
	output wire CH3VOL[0];
	output wire CH3VOL[1];
	output wire PSGDAC0[0];
	output wire PSGDAC0[1];
	output wire PSGDAC0[2];
	output wire PSGDAC0[3];
	output wire PSGDAC0[4];
	output wire PSGDAC0[5];
	output wire PSGDAC0[6];
	output wire PSGDAC0[7];
	output wire PSGDAC1[0];
	output wire PSGDAC1[1];
	output wire PSGDAC1[2];
	output wire PSGDAC1[3];
	output wire PSGDAC1[4];
	output wire PSGDAC1[5];
	output wire PSGDAC1[6];
	output wire PSGDAC1[7];
	output wire PSGDAC2[0];
	output wire PSGDAC2[1];
	output wire PSGDAC2[2];
	output wire PSGDAC2[3];
	output wire PSGDAC2[4];
	output wire PSGDAC2[5];
	output wire PSGDAC2[6];
	output wire PSGDAC2[7];
	output wire PSGDAC3[0];
	output wire PSGDAC3[1];
	output wire PSGDAC3[2];
	output wire PSGDAC3[3];
	output wire PSGDAC3[4];
	output wire PSGDAC3[5];
	output wire PSGDAC3[6];
	output wire PSGDAC3[7];
	input wire CAi[22];
	output wire CAo[22];
	output wire CA[19];
	output wire DTACK_OUT;
	output wire Z80_INT;
	output wire RA[7];
	output wire RA[6];
	output wire RA[5];
	output wire RA[4];
	output wire RA[2];
	output wire RA[1];
	output wire RA[0];
	output wire nRAS0;
	output wire RA[3];
	output wire nCAS0;
	output wire nOE0;
	output wire nLWR;
	output wire nUWR;
	input wire DTACK_IN;
	input wire RnW;
	input wire nLDS;
	input wire nUDS;
	input wire nAS;
	input wire nM1;
	input wire nWR;
	input wire nRD;
	input wire nIORQ;
	output wire nILP2;
	output wire nILP1;
	input wire nINTAK;
	input wire nMREQ;
	input wire nBG;
	output wire BGACK_OUT;
	input wire BGACK_IN;
	output wire nBR;
	output wire VSYNC;
	output wire nCSYNC;
	input wire nCSYNC_IN;
	output wire nHSYNC;
	input wire nHSYNC_IN;
	inout wire DB[15];
	inout wire DB[14];
	inout wire DB[13];
	inout wire DB[12];
	inout wire DB[11];
	inout wire DB[10];
	inout wire DB[9];
	inout wire DB[8];
	inout wire DB[7];
	inout wire DB[6];
	inout wire DB[5];
	inout wire DB[4];
	inout wire DB[3];
	inout wire DB[2];
	inout wire DB[1];
	inout wire DB[0];
	inout wire CA[0];
	inout wire CA[1];
	inout wire CA[2];
	inout wire CA[3];
	inout wire CA[4];
	inout wire CA[5];
	inout wire CA[6];
	inout wire CA[7];
	inout wire CA[8];
	inout wire CA[9];
	inout wire CA[10];
	inout wire CA[11];
	inout wire CA[12];
	inout wire CA[13];
	inout wire CA[14];
	inout wire CA[15];
	inout wire CA[16];
	inout wire CA[17];
	output wire CA[18];
	inout wire CA[20];
	inout wire CA[21];
	output wire R_DAC[0];
	output wire R_DAC[1];
	output wire R_DAC[2];
	output wire R_DAC[3];
	output wire R_DAC[4];
	output wire R_DAC[5];
	output wire R_DAC[6];
	output wire R_DAC[7];
	output wire R_DAC[8];
	output wire G_DAC[0];
	output wire G_DAC[1];
	output wire G_DAC[2];
	output wire G_DAC[3];
	output wire G_DAC[4];
	output wire G_DAC[5];
	output wire G_DAC[6];
	output wire G_DAC[7];
	output wire G_DAC[8];
	output wire R_DAC[9];
	output wire R_DAC[10];
	output wire R_DAC[11];
	output wire R_DAC[12];
	output wire R_DAC[13];
	output wire R_DAC[14];
	output wire R_DAC[15];
	output wire R_DAC[16];
	output wire B_DAC[0];
	output wire B_DAC[1];
	output wire B_DAC[2];
	output wire B_DAC[3];
	output wire B_DAC[4];
	output wire B_DAC[5];
	output wire B_DAC[6];
	output wire B_DAC[7];
	output wire B_DAC[8];
	output wire G_DAC[9];
	output wire G_DAC[10];
	output wire G_DAC[11];
	output wire G_DAC[12];
	output wire G_DAC[13];
	output wire G_DAC[14];
	output wire G_DAC[15];
	output wire G_DAC[16];
	output wire B_DAC[9];
	output wire B_DAC[10];
	output wire B_DAC[11];
	output wire B_DAC[12];
	output wire B_DAC[13];
	output wire B_DAC[14];
	output wire B_DAC[15];
	output wire B_DAC[16];
	output wire nOE1;
	output wire nWE0;
	output wire nWE1;
	output wire nCAS1;
	output wire nRAS1;
	output wire AD_RD_DIR;
	output wire nYS;
	output wire nSC;
	output wire nSE0_1;
	output wire ADo[7];
	output wire ADo[6];
	output wire ADo[5];
	output wire ADo[4];
	output wire ADo[3];
	output wire ADo[2];
	output wire ADo[1];
	output wire ADo[0];
	output wire RDo[6];
	output wire RDo[5];
	output wire RDo[4];
	output wire RDo[3];
	output wire RDo[2];
	output wire RDo[1];
	output wire RDo[0];
	input wire RDi[6];
	input wire RDi[7];
	input wire RDi[4];
	input wire RDi[5];
	input wire RDi[2];
	input wire RDi[3];
	input wire RDi[0];
	input wire RDi[1];
	input wire ADi[6];
	input wire ADi[7];
	input wire ADi[4];
	input wire ADi[5];
	input wire ADi[2];
	input wire ADi[3];
	input wire ADi[0];
	input wire ADi[1];
	output wire RDo[7];
	input wire SD[7];
	input wire SD[6];
	input wire SD[5];
	input wire SD[4];
	input wire SD[3];
	input wire SD[2];
	input wire SD[1];
	input wire SD[0];
	output wire CLK1;
	output wire CLK0;
	input wire EDCLKi;
	output wire EDCLKo;
	input wire MCLK;
	output wire SUB_CLK;
	input wire nRES_PAD;
	input wire 68kCLKi;
	output wire EDCLKd;
	output wire CA_PAD_DIR;
	output wire DB_PAD_DIR;
	input wire SEL0_M3;
	input wire nPAL;
	input wire nHL;
	output wire SPA/Bo;
	input wire SPA/Bi;

	// Wires

	wire w1;
	wire H40;
	wire w3;
	wire w4;
	wire w5;
	wire w6;
	wire w7;
	wire w8;
	wire w9;
	wire w10;
	wire w11;
	wire w12;
	wire w13;
	wire w14;
	wire w15;
	wire w16;
	wire w17;
	wire w18;
	wire w19;
	wire w20;
	wire w21;
	wire w22;
	wire w23;
	wire w24;
	wire w25;
	wire w26;
	wire w27;
	wire w28;
	wire w29;
	wire w30;
	wire w31;
	wire w32;
	wire w33;
	wire w34;
	wire w35;
	wire w36;
	wire w37;
	wire w38;
	wire w39;
	wire w40;
	wire w41;
	wire w42;
	wire w43;
	wire w44;
	wire w45;
	wire w46;
	wire w47;
	wire w48;
	wire ODD/EVEN;
	wire w50;
	wire w51;
	wire w52;
	wire w53;
	wire w54;
	wire w55;
	wire w56;
	wire w57;
	wire w58;
	wire w59;
	wire FIFOo[7];
	wire FIFOo[6];
	wire FIFOo[5];
	wire FIFOo[4];
	wire FIFOo[3];
	wire FIFOo[2];
	wire FIFOo[1];
	wire FIFOo[0];
	wire w68;
	wire w69;
	wire w70;
	wire w71;
	wire w72;
	wire w73;
	wire w74;
	wire w75;
	wire w76;
	wire w77;
	wire w78;
	wire w79;
	wire w80;
	wire w81;
	wire w82;
	wire w83;
	wire VRAMA[8];
	wire w85;
	wire w86;
	wire w87;
	wire w88;
	wire w89;
	wire w90;
	wire w91;
	wire w92;
	wire w93;
	wire w94;
	wire w95;
	wire w96;
	wire w97;
	wire w98;
	wire w99;
	wire w100;
	wire w101;
	wire VPOS[9];
	wire w103;
	wire w104;
	wire w105;
	wire w106;
	wire HPOS[0];
	wire w108;
	wire w109;
	wire w110;
	wire w111;
	wire w112;
	wire w113;
	wire w114;
	wire w115;
	wire w116;
	wire VPOS[8];
	wire w118;
	wire w119;
	wire w120;
	wire w121;
	wire w122;
	wire w123;
	wire w124;
	wire w125;
	wire w126;
	wire w127;
	wire w128;
	wire w129;
	wire w130;
	wire w131;
	wire w132;
	wire w133;
	wire w134;
	wire AD_DATA[7];
	wire AD_DATA[6];
	wire AD_DATA[4];
	wire RD_DATA[2];
	wire RD_DATA[1];
	wire RD_DATA[0];
	wire AD_DATA[5];
	wire w142;
	wire w143;
	wire DCLK1;
	wire DCLK2;
	wire nDCLK1;
	wire nDCLK2;
	wire HCLK1;
	wire HCLK2;
	wire nHCLK1;
	wire nHCLK2;
	wire SYSRES;
	wire DB[0];
	wire DB[1];
	wire DB[2];
	wire w156;
	wire DB[4];
	wire DB[5];
	wire DB[6];
	wire w160;
	wire DB[8];
	wire DB[9];
	wire AD_DATA[3];
	wire AD_DATA[2];
	wire AD_DATA[1];
	wire AD_DATA[0];
	wire DB[14];
	wire DB[13];
	wire DB[12];
	wire w170;
	wire DB[10];
	wire w172;
	wire M5;
	wire w174;
	wire w175;
	wire w176;
	wire HPOS[1];
	wire w178;
	wire w179;
	wire w180;
	wire w181;
	wire w182;
	wire w183;
	wire w184;
	wire w185;
	wire w186;
	wire w187;
	wire w188;
	wire w189;
	wire w190;
	wire VPOS[2];
	wire HPOS[3];
	wire w193;
	wire w194;
	wire w195;
	wire w196;
	wire w197;
	wire w198;
	wire w199;
	wire w200;
	wire w201;
	wire w202;
	wire w203;
	wire w204;
	wire w205;
	wire VPOS[4];
	wire HPOS[5];
	wire w208;
	wire RD_DATA[4];
	wire w210;
	wire w211;
	wire w212;
	wire w213;
	wire w214;
	wire w215;
	wire w216;
	wire w217;
	wire w218;
	wire w219;
	wire w220;
	wire w221;
	wire HPOS[7];
	wire w223;
	wire RD_DATA[6];
	wire w225;
	wire w226;
	wire w227;
	wire w228;
	wire w229;
	wire w230;
	wire w231;
	wire w232;
	wire w233;
	wire w234;
	wire w235;
	wire w236;
	wire w237;
	wire w238;
	wire w239;
	wire w240;
	wire w241;
	wire w242;
	wire w243;
	wire w244;
	wire w245;
	wire w246;
	wire w247;
	wire w248;
	wire w249;
	wire w250;
	wire w251;
	wire w252;
	wire w253;
	wire w254;
	wire w255;
	wire w256;
	wire w257;
	wire w258;
	wire w259;
	wire w260;
	wire w261;
	wire w262;
	wire w263;
	wire w264;
	wire w265;
	wire w266;
	wire w267;
	wire w268;
	wire w269;
	wire w270;
	wire w271;
	wire w272;
	wire w273;
	wire w274;
	wire w275;
	wire w276;
	wire w277;
	wire w278;
	wire w279;
	wire w280;
	wire w281;
	wire w282;
	wire w283;
	wire w284;
	wire w285;
	wire w286;
	wire w287;
	wire w288;
	wire w289;
	wire w290;
	wire w291;
	wire w292;
	wire w293;
	wire w294;
	wire w295;
	wire w296;
	wire w297;
	wire w298;
	wire w299;
	wire w300;
	wire w301;
	wire w302;
	wire w303;
	wire w304;
	wire w305;
	wire w306;
	wire w307;
	wire w308;
	wire w309;
	wire HPOS[2];
	wire VPOS[1];
	wire w312;
	wire w313;
	wire w314;
	wire w315;
	wire w316;
	wire w317;
	wire w318;
	wire w319;
	wire w320;
	wire w321;
	wire w322;
	wire VPOS[3];
	wire w324;
	wire w325;
	wire HPOS[4];
	wire w327;
	wire w328;
	wire w329;
	wire w330;
	wire w331;
	wire w332;
	wire w333;
	wire w334;
	wire w335;
	wire w336;
	wire w337;
	wire w338;
	wire w339;
	wire HPOS[6];
	wire VPOS[5];
	wire RD_DATA[5];
	wire w343;
	wire w344;
	wire w345;
	wire w346;
	wire w347;
	wire w348;
	wire w349;
	wire w350;
	wire w351;
	wire w352;
	wire w353;
	wire w354;
	wire w355;
	wire HPOS[8];
	wire VPOS[7];
	wire w358;
	wire w359;
	wire w360;
	wire w361;
	wire w362;
	wire w363;
	wire w364;
	wire w365;
	wire w366;
	wire w367;
	wire w368;
	wire w369;
	wire w370;
	wire w371;
	wire w372;
	wire w373;
	wire w374;
	wire w375;
	wire w376;
	wire w377;
	wire w378;
	wire w379;
	wire w380;
	wire w381;
	wire w382;
	wire w383;
	wire w384;
	wire w385;
	wire w386;
	wire w387;
	wire w388;
	wire w389;
	wire w390;
	wire w391;
	wire w392;
	wire w393;
	wire w394;
	wire w395;
	wire w396;
	wire w397;
	wire w398;
	wire w399;
	wire w400;
	wire w401;
	wire w402;
	wire w403;
	wire w404;
	wire w405;
	wire w406;
	wire w407;
	wire w408;
	wire w409;
	wire w410;
	wire w411;
	wire w412;
	wire w413;
	wire w414;
	wire w415;
	wire w416;
	wire w417;
	wire w418;
	wire w419;
	wire w420;
	wire w421;
	wire w422;
	wire w423;
	wire w424;
	wire w425;
	wire w426;
	wire w427;
	wire w428;
	wire w429;
	wire w430;
	wire w431;
	wire w432;
	wire w433;
	wire w434;
	wire w435;
	wire w436;
	wire w437;
	wire 128k;
	wire w439;
	wire w440;
	wire w441;
	wire w442;
	wire w443;
	wire w444;
	wire w445;
	wire w446;
	wire w447;
	wire w448;
	wire w449;
	wire w450;
	wire w451;
	wire w452;
	wire w453;
	wire w454;
	wire w455;
	wire w456;
	wire w457;
	wire w458;
	wire w459;
	wire w460;
	wire w461;
	wire w462;
	wire w463;
	wire w464;
	wire w465;
	wire w466;
	wire w467;
	wire w468;
	wire w469;
	wire w470;
	wire w471;
	wire w472;
	wire w473;
	wire w474;
	wire CA[0];
	wire w476;
	wire w477;
	wire w478;
	wire w479;
	wire w480;
	wire w481;
	wire w482;
	wire w483;
	wire w484;
	wire w485;
	wire w486;
	wire w487;
	wire w488;
	wire w489;
	wire w490;
	wire w491;
	wire w492;
	wire w493;
	wire w494;
	wire w495;
	wire w496;
	wire w497;
	wire w498;
	wire w499;
	wire w500;
	wire w501;
	wire w502;
	wire w503;
	wire w504;
	wire w505;
	wire w506;
	wire w507;
	wire w508;
	wire w509;
	wire w510;
	wire w511;
	wire w512;
	wire w513;
	wire w514;
	wire w515;
	wire w516;
	wire w517;
	wire w518;
	wire w519;
	wire w520;
	wire w521;
	wire w522;
	wire w523;
	wire w524;
	wire w525;
	wire w526;
	wire w527;
	wire w528;
	wire w529;
	wire w530;
	wire w531;
	wire w532;
	wire w533;
	wire w534;
	wire w535;
	wire w536;
	wire w537;
	wire w538;
	wire w539;
	wire w540;
	wire w541;
	wire w542;
	wire w543;
	wire w544;
	wire w545;
	wire w546;
	wire w547;
	wire w548;
	wire w549;
	wire w550;
	wire w551;
	wire w552;
	wire w553;
	wire w554;
	wire w555;
	wire w556;
	wire w557;
	wire w558;
	wire w559;
	wire w560;
	wire w561;
	wire w562;
	wire w563;
	wire w564;
	wire w565;
	wire w566;
	wire VRAMA[0];
	wire w568;
	wire w569;
	wire w570;
	wire w571;
	wire w572;
	wire w573;
	wire w574;
	wire w575;
	wire w576;
	wire w577;
	wire w578;
	wire w579;
	wire w580;
	wire w581;
	wire w582;
	wire w583;
	wire w584;
	wire w585;
	wire w586;
	wire w587;
	wire w588;
	wire w589;
	wire w590;
	wire w591;
	wire w592;
	wire w593;
	wire w594;
	wire w595;
	wire w596;
	wire w597;
	wire w598;
	wire w599;
	wire w600;
	wire w601;
	wire w602;
	wire w603;
	wire DMA_BUSY;
	wire w605;
	wire w606;
	wire w607;
	wire w608;
	wire w609;
	wire w610;
	wire w611;
	wire w612;
	wire w613;
	wire w614;
	wire w615;
	wire w616;
	wire w617;
	wire w618;
	wire w619;
	wire w620;
	wire w621;
	wire w622;
	wire w623;
	wire w624;
	wire w625;
	wire w626;
	wire w627;
	wire w628;
	wire w629;
	wire w630;
	wire w631;
	wire w632;
	wire w633;
	wire w634;
	wire w635;
	wire w636;
	wire w637;
	wire w638;
	wire w639;
	wire w640;
	wire w641;
	wire CA[8];
	wire CA[7];
	wire w644;
	wire w645;
	wire w646;
	wire w647;
	wire w648;
	wire w649;
	wire w650;
	wire w651;
	wire w652;
	wire w653;
	wire w654;
	wire w655;
	wire w656;
	wire CA[9];
	wire w658;
	wire VRAMA[7];
	wire w660;
	wire w661;
	wire VRAMA[9];
	wire w663;
	wire CA[6];
	wire w665;
	wire w666;
	wire w667;
	wire w668;
	wire w669;
	wire w670;
	wire w671;
	wire w672;
	wire w673;
	wire w674;
	wire w675;
	wire w676;
	wire w677;
	wire w678;
	wire w679;
	wire w680;
	wire w681;
	wire VRAMA[10];
	wire VRAMA[6];
	wire w684;
	wire w685;
	wire w686;
	wire w687;
	wire w688;
	wire w689;
	wire CA[10];
	wire w691;
	wire w692;
	wire w693;
	wire w694;
	wire w695;
	wire w696;
	wire w697;
	wire w698;
	wire w699;
	wire CA[11];
	wire w701;
	wire w702;
	wire w703;
	wire w704;
	wire w705;
	wire w706;
	wire w707;
	wire w708;
	wire w709;
	wire w710;
	wire VRAMA[5];
	wire w712;
	wire w713;
	wire VRAMA[11];
	wire CA[5];
	wire w716;
	wire w717;
	wire w718;
	wire w719;
	wire VRAMA[12];
	wire VRAMA[4];
	wire w722;
	wire w723;
	wire w724;
	wire w725;
	wire w726;
	wire CA[12];
	wire w728;
	wire w729;
	wire CA[4];
	wire w731;
	wire w732;
	wire w733;
	wire w734;
	wire CA[19];
	wire w736;
	wire w737;
	wire w738;
	wire w739;
	wire w740;
	wire VRAMA[13];
	wire w742;
	wire w743;
	wire w744;
	wire VRAMA[3];
	wire CA[3];
	wire w747;
	wire w748;
	wire CA[13];
	wire CA[20];
	wire w751;
	wire w752;
	wire w753;
	wire w754;
	wire w755;
	wire w756;
	wire VRAMA[14];
	wire VRAMA[2];
	wire w759;
	wire w760;
	wire w761;
	wire w762;
	wire w763;
	wire CA[2];
	wire w765;
	wire w766;
	wire w767;
	wire CA[21];
	wire w769;
	wire w770;
	wire w771;
	wire w772;
	wire w773;
	wire CA[14];
	wire w775;
	wire w776;
	wire VRAMA[15];
	wire CA[15];
	wire VRAMA[1];
	wire w780;
	wire w781;
	wire w782;
	wire w783;
	wire w784;
	wire w785;
	wire w786;
	wire w787;
	wire w788;
	wire w789;
	wire w790;
	wire CA[17];
	wire CA[1];
	wire VRAMA[16];
	wire w794;
	wire w795;
	wire CA[16];
	wire w797;
	wire w798;
	wire w799;
	wire w800;
	wire w801;
	wire w802;
	wire w803;
	wire w804;
	wire w805;
	wire w806;
	wire w807;
	wire w808;
	wire w809;
	wire w810;
	wire w811;
	wire w812;
	wire w813;
	wire w814;
	wire w815;
	wire w816;
	wire w817;
	wire w818;
	wire w819;
	wire w820;
	wire w821;
	wire w822;
	wire w823;
	wire w824;
	wire w825;
	wire w826;
	wire w827;
	wire w828;
	wire w829;
	wire w830;
	wire w831;
	wire w832;
	wire w833;
	wire w834;
	wire w835;
	wire w836;
	wire w837;
	wire w838;
	wire w839;
	wire w840;
	wire w841;
	wire w842;
	wire w843;
	wire w844;
	wire w845;
	wire w846;
	wire w847;
	wire w848;
	wire w849;
	wire w850;
	wire w851;
	wire w852;
	wire w853;
	wire w854;
	wire w855;
	wire w856;
	wire w857;
	wire w858;
	wire w859;
	wire w860;
	wire w861;
	wire w862;
	wire w863;
	wire w864;
	wire w865;
	wire w866;
	wire w867;
	wire w868;
	wire w869;
	wire w870;
	wire w871;
	wire w872;
	wire w873;
	wire w874;
	wire w875;
	wire w876;
	wire w877;
	wire w878;
	wire w879;
	wire w880;
	wire w881;
	wire w882;
	wire w883;
	wire w884;
	wire w885;
	wire w886;
	wire w887;
	wire w888;
	wire w889;
	wire w890;
	wire w891;
	wire w892;
	wire w893;
	wire w894;
	wire w895;
	wire w896;
	wire w897;
	wire w898;
	wire w899;
	wire w900;
	wire w901;
	wire w902;
	wire w903;
	wire w904;
	wire w905;
	wire w906;
	wire w907;
	wire w908;
	wire w909;
	wire w910;
	wire w911;
	wire w912;
	wire w913;
	wire w914;
	wire w915;
	wire w916;
	wire w917;
	wire w918;
	wire w919;
	wire w920;
	wire w921;
	wire w922;
	wire w923;
	wire w924;
	wire w925;
	wire w926;
	wire w927;
	wire w928;
	wire w929;
	wire w930;
	wire w931;
	wire w932;
	wire w933;
	wire w934;
	wire w935;
	wire w936;
	wire w937;
	wire w938;
	wire w939;
	wire w940;
	wire w941;
	wire w942;
	wire w943;
	wire w944;
	wire w945;
	wire w946;
	wire w947;
	wire w948;
	wire w949;
	wire w950;
	wire w951;
	wire w952;
	wire w953;
	wire w954;
	wire w955;
	wire w956;
	wire w957;
	wire w958;
	wire w959;
	wire w960;
	wire w961;
	wire w962;
	wire w963;
	wire w964;
	wire w965;
	wire w966;
	wire w967;
	wire w968;
	wire w969;
	wire w970;
	wire w971;
	wire w972;
	wire w973;
	wire w974;
	wire w975;
	wire w976;
	wire w977;
	wire w978;
	wire w979;
	wire w980;
	wire w981;
	wire w982;
	wire w983;
	wire w984;
	wire w985;
	wire w986;
	wire w987;
	wire w988;
	wire w989;
	wire w990;
	wire w991;
	wire w992;
	wire w993;
	wire w994;
	wire w995;
	wire w996;
	wire w997;
	wire w998;
	wire w999;
	wire w1000;
	wire w1001;
	wire w1002;
	wire w1003;
	wire w1004;
	wire w1005;
	wire w1006;
	wire w1007;
	wire w1008;
	wire w1009;
	wire w1010;
	wire w1011;
	wire w1012;
	wire w1013;
	wire w1014;
	wire w1015;
	wire w1016;
	wire w1017;
	wire w1018;
	wire w1019;
	wire w1020;
	wire w1021;
	wire w1022;
	wire w1023;
	wire w1024;
	wire w1025;
	wire w1026;
	wire w1027;
	wire w1028;
	wire w1029;
	wire w1030;
	wire w1031;
	wire w1032;
	wire w1033;
	wire w1034;
	wire w1035;
	wire w1036;
	wire w1037;
	wire w1038;
	wire w1039;
	wire w1040;
	wire w1041;
	wire w1042;
	wire w1043;
	wire w1044;
	wire w1045;
	wire w1046;
	wire w1047;
	wire w1048;
	wire w1049;
	wire w1050;
	wire w1051;
	wire w1052;
	wire w1053;
	wire w1054;
	wire w1055;
	wire w1056;
	wire w1057;
	wire w1058;
	wire w1059;
	wire w1060;
	wire w1061;
	wire w1062;
	wire w1063;
	wire VPOS[0];
	wire w1065;
	wire w1066;
	wire w1067;
	wire w1068;
	wire w1069;
	wire w1070;
	wire w1071;
	wire w1072;
	wire w1073;
	wire w1074;
	wire w1075;
	wire w1076;
	wire w1077;
	wire w1078;
	wire w1079;
	wire w1080;
	wire w1081;
	wire w1082;
	wire w1083;
	wire w1084;
	wire w1085;
	wire w1086;
	wire COL[0];
	wire COL[1];
	wire COL[2];
	wire COL[3];
	wire COL[4];
	wire COL[5];
	wire COL[6];
	wire w1094;
	wire w1095;
	wire w1096;
	wire w1097;
	wire w1098;
	wire w1099;
	wire w1100;
	wire w1101;
	wire w1102;
	wire w1103;
	wire w1104;
	wire w1105;
	wire w1106;
	wire w1107;
	wire w1108;
	wire w1109;
	wire w1110;
	wire w1111;
	wire w1112;
	wire w1113;
	wire w1114;
	wire w1115;
	wire w1116;
	wire w1117;
	wire w1118;
	wire w1119;
	wire w1120;
	wire w1121;
	wire w1122;
	wire w1123;
	wire w1124;
	wire w1125;
	wire w1126;
	wire w1127;
	wire w1128;
	wire w1129;
	wire w1130;
	wire w1131;
	wire w1132;
	wire w1133;
	wire w1134;
	wire w1135;
	wire w1136;
	wire w1137;
	wire w1138;
	wire w1139;
	wire w1140;
	wire w1141;
	wire w1142;
	wire w1143;
	wire w1144;
	wire w1145;
	wire w1146;
	wire w1147;
	wire w1148;
	wire w1149;
	wire w1150;
	wire w1151;
	wire w1152;
	wire w1153;
	wire w1154;
	wire w1155;
	wire w1156;
	wire w1157;
	wire w1158;
	wire w1159;
	wire w1160;
	wire w1161;
	wire w1162;
	wire w1163;
	wire w1164;
	wire w1165;
	wire w1166;
	wire w1167;
	wire w1168;
	wire w1169;
	wire w1170;
	wire w1171;
	wire w1172;
	wire w1173;
	wire w1174;
	wire w1175;
	wire w1176;
	wire w1177;
	wire w1178;
	wire w1179;
	wire w1180;
	wire w1181;
	wire w1182;
	wire w1183;
	wire w1184;
	wire w1185;
	wire w1186;
	wire w1187;
	wire w1188;
	wire w1189;
	wire w1190;
	wire w1191;
	wire w1192;
	wire w1193;
	wire w1194;
	wire w1195;
	wire w1196;
	wire w1197;
	wire w1198;
	wire w1199;
	wire w1200;
	wire w1201;
	wire w1202;
	wire w1203;
	wire w1204;
	wire w1205;
	wire w1206;
	wire w1207;
	wire w1208;
	wire w1209;
	wire w1210;
	wire w1211;
	wire w1212;
	wire w1213;
	wire w1214;
	wire w1215;
	wire w1216;
	wire w1217;
	wire w1218;
	wire w1219;
	wire w1220;
	wire w1221;
	wire w1222;
	wire w1223;
	wire w1224;
	wire w1225;
	wire w1226;
	wire w1227;
	wire w1228;
	wire w1229;
	wire w1230;
	wire w1231;
	wire w1232;
	wire w1233;
	wire w1234;
	wire w1235;
	wire w1236;
	wire w1237;
	wire w1238;
	wire w1239;
	wire w1240;
	wire w1241;
	wire w1242;
	wire w1243;
	wire w1244;
	wire w1245;
	wire w1246;
	wire w1247;
	wire w1248;
	wire w1249;
	wire w1250;
	wire w1251;
	wire w1252;
	wire w1253;
	wire w1254;
	wire w1255;
	wire w1256;
	wire w1257;
	wire w1258;
	wire w1259;
	wire w1260;
	wire w1261;
	wire w1262;
	wire w1263;
	wire w1264;
	wire w1265;
	wire w1266;
	wire w1267;
	wire w1268;
	wire w1269;
	wire w1270;
	wire w1271;
	wire w1272;
	wire w1273;
	wire w1274;
	wire w1275;
	wire w1276;
	wire w1277;
	wire w1278;
	wire w1279;
	wire w1280;
	wire w1281;
	wire w1282;
	wire w1283;
	wire w1284;
	wire w1285;
	wire w1286;
	wire w1287;
	wire w1288;
	wire w1289;
	wire w1290;
	wire w1291;
	wire w1292;
	wire w1293;
	wire w1294;
	wire w1295;
	wire w1296;
	wire w1297;
	wire w1298;
	wire w1299;
	wire w1300;
	wire w1301;
	wire w1302;
	wire w1303;
	wire w1304;
	wire w1305;
	wire w1306;
	wire w1307;
	wire w1308;
	wire w1309;
	wire w1310;
	wire w1311;
	wire w1312;
	wire w1313;
	wire w1314;
	wire w1315;
	wire w1316;
	wire w1317;
	wire w1318;
	wire w1319;
	wire w1320;
	wire w1321;
	wire w1322;
	wire w1323;
	wire w1324;
	wire w1325;
	wire w1326;
	wire w1327;
	wire w1328;
	wire w1329;
	wire w1330;
	wire w1331;
	wire w1332;
	wire w1333;
	wire w1334;
	wire w1335;
	wire w1336;
	wire w1337;
	wire w1338;
	wire w1339;
	wire w1340;
	wire w1341;
	wire w1342;
	wire w1343;
	wire w1344;
	wire w1345;
	wire w1346;
	wire w1347;
	wire w1348;
	wire w1349;
	wire w1350;
	wire w1351;
	wire w1352;
	wire w1353;
	wire w1354;
	wire w1355;
	wire w1356;
	wire w1357;
	wire w1358;
	wire w1359;
	wire w1360;
	wire w1361;
	wire w1362;
	wire w1363;
	wire w1364;
	wire w1365;
	wire w1366;
	wire w1367;
	wire w1368;
	wire w1369;
	wire w1370;
	wire w1371;
	wire w1372;
	wire w1373;
	wire w1374;
	wire w1375;
	wire w1376;
	wire w1377;
	wire w1378;
	wire w1379;
	wire w1380;
	wire w1381;
	wire w1382;
	wire w1383;
	wire w1384;
	wire w1385;
	wire w1386;
	wire w1387;
	wire w1388;
	wire w1389;
	wire w1390;
	wire w1391;
	wire w1392;
	wire w1393;
	wire w1394;
	wire w1395;
	wire w1396;
	wire w1397;
	wire w1398;
	wire VRAM_REFRESH;
	wire w1400;
	wire w1401;
	wire w1402;
	wire w1403;
	wire w1404;
	wire w1405;
	wire w1406;
	wire w1407;
	wire w1408;
	wire w1409;
	wire w1410;
	wire w1411;
	wire w1412;
	wire w1413;
	wire w1414;
	wire w1415;
	wire w1416;
	wire w1417;
	wire w1418;
	wire w1419;
	wire w1420;
	wire w1421;
	wire w1422;
	wire w1423;
	wire w1424;
	wire w1425;
	wire w1426;
	wire w1427;
	wire w1428;
	wire w1429;
	wire w1430;
	wire w1431;
	wire w1432;
	wire w1433;
	wire w1434;
	wire w1435;
	wire w1436;
	wire w1437;
	wire w1438;
	wire w1439;
	wire w1440;
	wire w1441;
	wire w1442;
	wire w1443;
	wire w1444;
	wire w1445;
	wire w1446;
	wire w1447;
	wire w1448;
	wire w1449;
	wire w1450;
	wire w1451;
	wire w1452;
	wire w1453;
	wire w1454;
	wire w1455;
	wire w1456;
	wire w1457;
	wire w1458;
	wire w1459;
	wire w1460;
	wire w1461;
	wire w1462;
	wire w1463;
	wire w1464;
	wire w1465;
	wire w1466;
	wire w1467;
	wire w1468;
	wire w1469;
	wire w1470;
	wire w1471;
	wire w1472;
	wire w1473;
	wire w1474;
	wire w1475;
	wire w1476;
	wire w1477;
	wire w1478;
	wire w1479;
	wire w1480;
	wire w1481;
	wire w1482;
	wire w1483;
	wire w1484;
	wire w1485;
	wire w1486;
	wire w1487;
	wire w1488;
	wire w1489;
	wire w1490;
	wire w1491;
	wire w1492;
	wire w1493;
	wire w1494;
	wire w1495;
	wire w1496;
	wire w1497;
	wire w1498;
	wire w1499;
	wire w1500;
	wire w1501;
	wire w1502;
	wire w1503;
	wire w1504;
	wire w1505;
	wire w1506;
	wire w1507;
	wire w1508;
	wire w1509;
	wire w1510;
	wire w1511;
	wire CA[18];
	wire w1513;
	wire w1514;
	wire w1515;
	wire w1516;
	wire w1517;
	wire w1518;
	wire w1519;
	wire w1520;
	wire w1521;
	wire w1522;
	wire w1523;
	wire w1524;
	wire w1525;
	wire w1526;
	wire w1527;
	wire w1528;
	wire w1529;
	wire w1530;
	wire w1531;
	wire w1532;
	wire w1533;
	wire w1534;
	wire w1535;
	wire w1536;
	wire w1537;
	wire w1538;
	wire w1539;
	wire w1540;
	wire w1541;
	wire w1542;
	wire w1543;
	wire w1544;
	wire w1545;
	wire w1546;
	wire w1547;
	wire w1548;
	wire w1549;
	wire w1550;
	wire w1551;
	wire w1552;
	wire w1553;
	wire w1554;
	wire w1555;
	wire w1556;
	wire w1557;
	wire w1558;
	wire w1559;
	wire w1560;
	wire w1561;
	wire w1562;
	wire w1563;
	wire w1564;
	wire w1565;
	wire w1566;
	wire w1567;
	wire w1568;
	wire w1569;
	wire w1570;
	wire w1571;
	wire w1572;
	wire w1573;
	wire VPOS[6];
	wire w1575;
	wire w1576;
	wire w1577;
	wire w1578;
	wire w1579;
	wire w1580;
	wire w1581;
	wire w1582;
	wire w1583;
	wire w1584;
	wire w1585;
	wire w1586;
	wire w1587;
	wire w1588;
	wire w1589;
	wire w1590;
	wire w1591;
	wire w1592;
	wire w1593;
	wire w1594;
	wire w1595;
	wire w1596;
	wire w1597;
	wire w1598;
	wire w1599;
	wire w1600;
	wire w1601;
	wire w1602;
	wire w1603;
	wire w1604;
	wire w1605;
	wire w1606;
	wire w1607;
	wire w1608;
	wire w1609;
	wire w1610;
	wire w1611;
	wire w1612;
	wire w1613;
	wire w1614;
	wire w1615;
	wire w1616;
	wire w1617;
	wire w1618;
	wire w1619;
	wire w1620;
	wire w1621;
	wire w1622;
	wire w1623;
	wire w1624;
	wire w1625;
	wire w1626;
	wire w1627;
	wire w1628;
	wire w1629;
	wire w1630;
	wire w1631;
	wire w1632;
	wire w1633;
	wire w1634;
	wire w1635;
	wire w1636;
	wire w1637;
	wire w1638;
	wire w1639;
	wire w1640;
	wire w1641;
	wire w1642;
	wire w1643;
	wire w1644;
	wire w1645;
	wire w1646;
	wire w1647;
	wire w1648;
	wire w1649;
	wire w1650;
	wire w1651;
	wire w1652;
	wire w1653;
	wire w1654;
	wire w1655;
	wire w1656;
	wire w1657;
	wire w1658;
	wire w1659;
	wire w1660;
	wire w1661;
	wire w1662;
	wire w1663;
	wire w1664;
	wire w1665;
	wire w1666;
	wire w1667;
	wire w1668;
	wire w1669;
	wire w1670;
	wire w1671;
	wire w1672;
	wire w1673;
	wire w1674;
	wire w1675;
	wire w1676;
	wire w1677;
	wire w1678;
	wire w1679;
	wire w1680;
	wire w1681;
	wire w1682;
	wire w1683;
	wire w1684;
	wire w1685;
	wire w1686;
	wire w1687;
	wire w1688;
	wire w1689;
	wire w1690;
	wire w1691;
	wire w1692;
	wire w1693;
	wire w1694;
	wire w1695;
	wire w1696;
	wire w1697;
	wire w1698;
	wire w1699;
	wire w1700;
	wire w1701;
	wire w1702;
	wire w1703;
	wire w1704;
	wire w1705;
	wire w1706;
	wire w1707;
	wire w1708;
	wire w1709;
	wire w1710;
	wire w1711;
	wire w1712;
	wire w1713;
	wire w1714;
	wire w1715;
	wire w1716;
	wire w1717;
	wire w1718;
	wire w1719;
	wire w1720;
	wire w1721;
	wire w1722;
	wire w1723;
	wire w1724;
	wire w1725;
	wire w1726;
	wire w1727;
	wire w1728;
	wire w1729;
	wire w1730;
	wire w1731;
	wire w1732;
	wire w1733;
	wire w1734;
	wire w1735;
	wire w1736;
	wire w1737;
	wire w1738;
	wire w1739;
	wire w1740;
	wire w1741;
	wire w1742;
	wire w1743;
	wire w1744;
	wire w1745;
	wire w1746;
	wire w1747;
	wire w1748;
	wire w1749;
	wire w1750;
	wire w1751;
	wire w1752;
	wire w1753;
	wire w1754;
	wire w1755;
	wire w1756;
	wire w1757;
	wire w1758;
	wire w1759;
	wire w1760;
	wire w1761;
	wire w1762;
	wire w1763;
	wire w1764;
	wire w1765;
	wire w1766;
	wire w1767;
	wire w1768;
	wire w1769;
	wire w1770;
	wire w1771;
	wire w1772;
	wire w1773;
	wire w1774;
	wire w1775;
	wire w1776;
	wire w1777;
	wire w1778;
	wire w1779;
	wire w1780;
	wire w1781;
	wire w1782;
	wire w1783;
	wire w1784;
	wire w1785;
	wire w1786;
	wire w1787;
	wire w1788;
	wire w1789;
	wire w1790;
	wire w1791;
	wire w1792;
	wire w1793;
	wire w1794;
	wire w1795;
	wire w1796;
	wire w1797;
	wire w1798;
	wire w1799;
	wire w1800;
	wire w1801;
	wire w1802;
	wire w1803;
	wire w1804;
	wire w1805;
	wire w1806;
	wire w1807;
	wire w1808;
	wire w1809;
	wire w1810;
	wire w1811;
	wire w1812;
	wire w1813;
	wire w1814;
	wire w1815;
	wire w1816;
	wire w1817;
	wire w1818;
	wire w1819;
	wire w1820;
	wire w1821;
	wire w1822;
	wire w1823;
	wire w1824;
	wire w1825;
	wire w1826;
	wire w1827;
	wire w1828;
	wire w1829;
	wire w1830;
	wire w1831;
	wire w1832;
	wire w1833;
	wire w1834;
	wire w1835;
	wire w1836;
	wire w1837;
	wire w1838;
	wire w1839;
	wire w1840;
	wire w1841;
	wire w1842;
	wire w1843;
	wire w1844;
	wire w1845;
	wire w1846;
	wire w1847;
	wire w1848;
	wire w1849;
	wire w1850;
	wire w1851;
	wire w1852;
	wire w1853;
	wire w1854;
	wire w1855;
	wire w1856;
	wire w1857;
	wire w1858;
	wire w1859;
	wire w1860;
	wire w1861;
	wire w1862;
	wire w1863;
	wire w1864;
	wire w1865;
	wire w1866;
	wire w1867;
	wire w1868;
	wire w1869;
	wire w1870;
	wire w1871;
	wire w1872;
	wire w1873;
	wire w1874;
	wire w1875;
	wire w1876;
	wire w1877;
	wire w1878;
	wire w1879;
	wire w1880;
	wire w1881;
	wire w1882;
	wire w1883;
	wire w1884;
	wire w1885;
	wire w1886;
	wire w1887;
	wire w1888;
	wire w1889;
	wire w1890;
	wire w1891;
	wire w1892;
	wire w1893;
	wire w1894;
	wire w1895;
	wire w1896;
	wire w1897;
	wire w1898;
	wire w1899;
	wire w1900;
	wire w1901;
	wire w1902;
	wire w1903;
	wire w1904;
	wire w1905;
	wire w1906;
	wire w1907;
	wire w1908;
	wire w1909;
	wire w1910;
	wire w1911;
	wire w1912;
	wire w1913;
	wire w1914;
	wire w1915;
	wire w1916;
	wire w1917;
	wire w1918;
	wire w1919;
	wire w1920;
	wire w1921;
	wire w1922;
	wire w1923;
	wire w1924;
	wire w1925;
	wire w1926;
	wire w1927;
	wire w1928;
	wire w1929;
	wire w1930;
	wire w1931;
	wire w1932;
	wire w1933;
	wire w1934;
	wire w1935;
	wire w1936;
	wire w1937;
	wire w1938;
	wire w1939;
	wire w1940;
	wire w1941;
	wire w1942;
	wire w1943;
	wire w1944;
	wire w1945;
	wire w1946;
	wire w1947;
	wire w1948;
	wire w1949;
	wire w1950;
	wire w1951;
	wire w1952;
	wire w1953;
	wire w1954;
	wire w1955;
	wire w1956;
	wire w1957;
	wire w1958;
	wire w1959;
	wire w1960;
	wire w1961;
	wire w1962;
	wire w1963;
	wire w1964;
	wire w1965;
	wire w1966;
	wire w1967;
	wire w1968;
	wire w1969;
	wire w1970;
	wire w1971;
	wire w1972;
	wire w1973;
	wire w1974;
	wire w1975;
	wire w1976;
	wire w1977;
	wire w1978;
	wire w1979;
	wire w1980;
	wire w1981;
	wire w1982;
	wire w1983;
	wire w1984;
	wire w1985;
	wire w1986;
	wire w1987;
	wire w1988;
	wire w1989;
	wire w1990;
	wire w1991;
	wire w1992;
	wire w1993;
	wire w1994;
	wire w1995;
	wire w1996;
	wire w1997;
	wire w1998;
	wire w1999;
	wire w2000;
	wire w2001;
	wire w2002;
	wire w2003;
	wire w2004;
	wire w2005;
	wire w2006;
	wire w2007;
	wire w2008;
	wire w2009;
	wire w2010;
	wire w2011;
	wire w2012;
	wire w2013;
	wire w2014;
	wire w2015;
	wire w2016;
	wire w2017;
	wire w2018;
	wire w2019;
	wire w2020;
	wire w2021;
	wire w2022;
	wire w2023;
	wire w2024;
	wire w2025;
	wire w2026;
	wire w2027;
	wire w2028;
	wire w2029;
	wire w2030;
	wire w2031;
	wire w2032;
	wire w2033;
	wire w2034;
	wire w2035;
	wire w2036;
	wire w2037;
	wire w2038;
	wire w2039;
	wire w2040;
	wire w2041;
	wire w2042;
	wire w2043;
	wire w2044;
	wire w2045;
	wire w2046;
	wire w2047;
	wire w2048;
	wire w2049;
	wire w2050;
	wire w2051;
	wire w2052;
	wire w2053;
	wire w2054;
	wire w2055;
	wire w2056;
	wire w2057;
	wire w2058;
	wire w2059;
	wire w2060;
	wire w2061;
	wire w2062;
	wire w2063;
	wire w2064;
	wire w2065;
	wire w2066;
	wire w2067;
	wire w2068;
	wire w2069;
	wire w2070;
	wire w2071;
	wire w2072;
	wire w2073;
	wire w2074;
	wire w2075;
	wire w2076;
	wire w2077;
	wire w2078;
	wire w2079;
	wire w2080;
	wire w2081;
	wire w2082;
	wire w2083;
	wire w2084;
	wire w2085;
	wire w2086;
	wire w2087;
	wire w2088;
	wire w2089;
	wire w2090;
	wire w2091;
	wire w2092;
	wire w2093;
	wire w2094;
	wire w2095;
	wire w2096;
	wire w2097;
	wire w2098;
	wire w2099;
	wire w2100;
	wire w2101;
	wire w2102;
	wire w2103;
	wire w2104;
	wire w2105;
	wire w2106;
	wire w2107;
	wire w2108;
	wire w2109;
	wire w2110;
	wire w2111;
	wire w2112;
	wire w2113;
	wire w2114;
	wire w2115;
	wire w2116;
	wire w2117;
	wire w2118;
	wire w2119;
	wire w2120;
	wire w2121;
	wire w2122;
	wire w2123;
	wire w2124;
	wire w2125;
	wire w2126;
	wire w2127;
	wire w2128;
	wire w2129;
	wire w2130;
	wire w2131;
	wire w2132;
	wire w2133;
	wire w2134;
	wire w2135;
	wire w2136;
	wire w2137;
	wire w2138;
	wire w2139;
	wire w2140;
	wire w2141;
	wire w2142;
	wire w2143;
	wire w2144;
	wire w2145;
	wire w2146;
	wire w2147;
	wire w2148;
	wire w2149;
	wire w2150;
	wire w2151;
	wire w2152;
	wire w2153;
	wire w2154;
	wire w2155;
	wire w2156;
	wire w2157;
	wire w2158;
	wire w2159;
	wire w2160;
	wire w2161;
	wire w2162;
	wire w2163;
	wire w2164;
	wire w2165;
	wire w2166;
	wire w2167;
	wire w2168;
	wire w2169;
	wire w2170;
	wire w2171;
	wire w2172;
	wire w2173;
	wire w2174;
	wire w2175;
	wire w2176;
	wire w2177;
	wire w2178;
	wire w2179;
	wire w2180;
	wire w2181;
	wire w2182;
	wire w2183;
	wire w2184;
	wire w2185;
	wire w2186;
	wire w2187;
	wire w2188;
	wire w2189;
	wire w2190;
	wire w2191;
	wire w2192;
	wire w2193;
	wire w2194;
	wire w2195;
	wire w2196;
	wire w2197;
	wire w2198;
	wire w2199;
	wire w2200;
	wire w2201;
	wire w2202;
	wire w2203;
	wire w2204;
	wire w2205;
	wire w2206;
	wire w2207;
	wire w2208;
	wire w2209;
	wire w2210;
	wire w2211;
	wire w2212;
	wire w2213;
	wire w2214;
	wire w2215;
	wire w2216;
	wire w2217;
	wire w2218;
	wire w2219;
	wire w2220;
	wire w2221;
	wire w2222;
	wire w2223;
	wire w2224;
	wire w2225;
	wire w2226;
	wire w2227;
	wire w2228;
	wire w2229;
	wire w2230;
	wire w2231;
	wire w2232;
	wire w2233;
	wire w2234;
	wire w2235;
	wire w2236;
	wire w2237;
	wire w2238;
	wire w2239;
	wire w2240;
	wire w2241;
	wire w2242;
	wire w2243;
	wire w2244;
	wire w2245;
	wire w2246;
	wire w2247;
	wire w2248;
	wire w2249;
	wire w2250;
	wire w2251;
	wire w2252;
	wire w2253;
	wire w2254;
	wire w2255;
	wire w2256;
	wire w2257;
	wire w2258;
	wire w2259;
	wire w2260;
	wire w2261;
	wire w2262;
	wire w2263;
	wire w2264;
	wire w2265;
	wire w2266;
	wire w2267;
	wire w2268;
	wire w2269;
	wire w2270;
	wire w2271;
	wire w2272;
	wire w2273;
	wire w2274;
	wire w2275;
	wire w2276;
	wire w2277;
	wire w2278;
	wire w2279;
	wire w2280;
	wire w2281;
	wire w2282;
	wire w2283;
	wire w2284;
	wire w2285;
	wire w2286;
	wire w2287;
	wire w2288;
	wire w2289;
	wire w2290;
	wire w2291;
	wire w2292;
	wire w2293;
	wire w2294;
	wire w2295;
	wire w2296;
	wire w2297;
	wire w2298;
	wire w2299;
	wire w2300;
	wire w2301;
	wire w2302;
	wire w2303;
	wire w2304;
	wire w2305;
	wire w2306;
	wire w2307;
	wire w2308;
	wire w2309;
	wire w2310;
	wire w2311;
	wire w2312;
	wire w2313;
	wire w2314;
	wire w2315;
	wire w2316;
	wire w2317;
	wire w2318;
	wire w2319;
	wire w2320;
	wire w2321;
	wire w2322;
	wire w2323;
	wire w2324;
	wire w2325;
	wire w2326;
	wire w2327;
	wire w2328;
	wire w2329;
	wire w2330;
	wire w2331;
	wire w2332;
	wire w2333;
	wire w2334;
	wire w2335;
	wire w2336;
	wire w2337;
	wire w2338;
	wire w2339;
	wire w2340;
	wire w2341;
	wire w2342;
	wire w2343;
	wire w2344;
	wire w2345;
	wire w2346;
	wire w2347;
	wire w2348;
	wire w2349;
	wire w2350;
	wire w2351;
	wire w2352;
	wire w2353;
	wire w2354;
	wire w2355;
	wire w2356;
	wire w2357;
	wire w2358;
	wire w2359;
	wire w2360;
	wire w2361;
	wire w2362;
	wire w2363;
	wire w2364;
	wire w2365;
	wire w2366;
	wire w2367;
	wire w2368;
	wire w2369;
	wire w2370;
	wire w2371;
	wire w2372;
	wire w2373;
	wire w2374;
	wire w2375;
	wire w2376;
	wire w2377;
	wire w2378;
	wire w2379;
	wire w2380;
	wire w2381;
	wire w2382;
	wire w2383;
	wire w2384;
	wire w2385;
	wire w2386;
	wire w2387;
	wire w2388;
	wire w2389;
	wire w2390;
	wire w2391;
	wire w2392;
	wire w2393;
	wire w2394;
	wire w2395;
	wire w2396;
	wire w2397;
	wire w2398;
	wire w2399;
	wire w2400;
	wire w2401;
	wire w2402;
	wire w2403;
	wire w2404;
	wire w2405;
	wire w2406;
	wire w2407;
	wire w2408;
	wire w2409;
	wire w2410;
	wire w2411;
	wire w2412;
	wire w2413;
	wire w2414;
	wire w2415;
	wire w2416;
	wire w2417;
	wire w2418;
	wire w2419;
	wire w2420;
	wire w2421;
	wire w2422;
	wire w2423;
	wire w2424;
	wire w2425;
	wire w2426;
	wire w2427;
	wire w2428;
	wire w2429;
	wire w2430;
	wire w2431;
	wire w2432;
	wire w2433;
	wire w2434;
	wire w2435;
	wire w2436;
	wire w2437;
	wire w2438;
	wire w2439;
	wire w2440;
	wire w2441;
	wire w2442;
	wire w2443;
	wire w2444;
	wire w2445;
	wire w2446;
	wire w2447;
	wire w2448;
	wire w2449;
	wire w2450;
	wire w2451;
	wire w2452;
	wire w2453;
	wire w2454;
	wire w2455;
	wire w2456;
	wire w2457;
	wire w2458;
	wire w2459;
	wire w2460;
	wire w2461;
	wire w2462;
	wire w2463;
	wire w2464;
	wire w2465;
	wire w2466;
	wire w2467;
	wire w2468;
	wire w2469;
	wire w2470;
	wire w2471;
	wire w2472;
	wire w2473;
	wire w2474;
	wire w2475;
	wire w2476;
	wire w2477;
	wire w2478;
	wire w2479;
	wire w2480;
	wire w2481;
	wire w2482;
	wire w2483;
	wire w2484;
	wire w2485;
	wire w2486;
	wire w2487;
	wire w2488;
	wire w2489;
	wire w2490;
	wire w2491;
	wire w2492;
	wire w2493;
	wire w2494;
	wire w2495;
	wire w2496;
	wire w2497;
	wire w2498;
	wire w2499;
	wire w2500;
	wire w2501;
	wire w2502;
	wire w2503;
	wire w2504;
	wire w2505;
	wire w2506;
	wire w2507;
	wire w2508;
	wire w2509;
	wire w2510;
	wire w2511;
	wire w2512;
	wire w2513;
	wire w2514;
	wire w2515;
	wire w2516;
	wire w2517;
	wire w2518;
	wire w2519;
	wire w2520;
	wire w2521;
	wire w2522;
	wire w2523;
	wire w2524;
	wire w2525;
	wire w2526;
	wire w2527;
	wire w2528;
	wire w2529;
	wire w2530;
	wire w2531;
	wire w2532;
	wire w2533;
	wire w2534;
	wire w2535;
	wire w2536;
	wire w2537;
	wire w2538;
	wire w2539;
	wire w2540;
	wire w2541;
	wire w2542;
	wire w2543;
	wire w2544;
	wire w2545;
	wire w2546;
	wire w2547;
	wire w2548;
	wire w2549;
	wire w2550;
	wire w2551;
	wire w2552;
	wire w2553;
	wire w2554;
	wire w2555;
	wire w2556;
	wire w2557;
	wire w2558;
	wire w2559;
	wire w2560;
	wire w2561;
	wire w2562;
	wire w2563;
	wire w2564;
	wire w2565;
	wire w2566;
	wire w2567;
	wire w2568;
	wire w2569;
	wire w2570;
	wire w2571;
	wire w2572;
	wire w2573;
	wire w2574;
	wire w2575;
	wire w2576;
	wire w2577;
	wire w2578;
	wire w2579;
	wire w2580;
	wire w2581;
	wire w2582;
	wire w2583;
	wire w2584;
	wire w2585;
	wire w2586;
	wire w2587;
	wire w2588;
	wire w2589;
	wire w2590;
	wire w2591;
	wire w2592;
	wire w2593;
	wire w2594;
	wire w2595;
	wire w2596;
	wire w2597;
	wire w2598;
	wire w2599;
	wire w2600;
	wire w2601;
	wire w2602;
	wire w2603;
	wire w2604;
	wire w2605;
	wire w2606;
	wire w2607;
	wire w2608;
	wire w2609;
	wire w2610;
	wire w2611;
	wire w2612;
	wire w2613;
	wire w2614;
	wire w2615;
	wire w2616;
	wire w2617;
	wire w2618;
	wire w2619;
	wire w2620;
	wire w2621;
	wire w2622;
	wire w2623;
	wire w2624;
	wire w2625;
	wire w2626;
	wire w2627;
	wire w2628;
	wire w2629;
	wire w2630;
	wire w2631;
	wire w2632;
	wire w2633;
	wire w2634;
	wire w2635;
	wire w2636;
	wire w2637;
	wire w2638;
	wire w2639;
	wire w2640;
	wire w2641;
	wire w2642;
	wire w2643;
	wire w2644;
	wire w2645;
	wire w2646;
	wire w2647;
	wire RES;
	wire w2649;
	wire w2650;
	wire w2651;
	wire w2652;
	wire EDCLK_O;
	wire nYS;
	wire w2655;
	wire w2656;
	wire w2657;
	wire w2658;
	wire w2659;
	wire w2660;
	wire w2661;
	wire w2662;
	wire w2663;
	wire w2664;
	wire w2665;
	wire w2666;
	wire w2667;
	wire w2668;
	wire w2669;
	wire w2670;
	wire w2671;
	wire w2672;
	wire w2673;
	wire w2674;
	wire w2675;
	wire w2676;
	wire w2677;
	wire w2678;
	wire w2679;
	wire w2680;
	wire w2681;
	wire w2682;
	wire w2683;
	wire w2684;
	wire w2685;
	wire w2686;
	wire w2687;
	wire w2688;
	wire w2689;
	wire w2690;
	wire w2691;
	wire w2692;
	wire w2693;
	wire w2694;
	wire w2695;
	wire w2696;
	wire w2697;
	wire w2698;
	wire w2699;
	wire w2700;
	wire w2701;
	wire w2702;
	wire w2703;
	wire w2704;
	wire w2705;
	wire w2706;
	wire w2707;
	wire w2708;
	wire w2709;
	wire w2710;
	wire w2711;
	wire w2712;
	wire w2713;
	wire w2714;
	wire w2715;
	wire w2716;
	wire w2717;
	wire w2718;
	wire w2719;
	wire w2720;
	wire w2721;
	wire w2722;
	wire SPR_PRIO;
	wire w2724;
	wire w2725;
	wire w2726;
	wire w2727;
	wire w2728;
	wire w2729;
	wire w2730;
	wire w2731;
	wire w2732;
	wire w2733;
	wire w2734;
	wire w2735;
	wire w2736;
	wire w2737;
	wire w2738;
	wire w2739;
	wire w2740;
	wire w2741;
	wire w2742;
	wire w2743;
	wire w2744;
	wire w2745;
	wire w2746;
	wire w2747;
	wire w2748;
	wire w2749;
	wire w2750;
	wire w2751;
	wire w2752;
	wire w2753;
	wire w2754;
	wire w2755;
	wire w2756;
	wire w2757;
	wire w2758;
	wire w2759;
	wire w2760;
	wire w2761;
	wire w2762;
	wire w2763;
	wire w2764;
	wire w2765;
	wire w2766;
	wire w2767;
	wire w2768;
	wire w2769;
	wire w2770;
	wire w2771;
	wire w2772;
	wire w2773;
	wire w2774;
	wire w2775;
	wire w2776;
	wire w2777;
	wire w2778;
	wire w2779;
	wire w2780;
	wire w2781;
	wire w2782;
	wire w2783;
	wire w2784;
	wire w2785;
	wire w2786;
	wire w2787;
	wire w2788;
	wire w2789;
	wire w2790;
	wire w2791;
	wire w2792;
	wire w2793;
	wire PLANE_A_PRIO;
	wire PLANE_B_PRIO;
	wire w2796;
	wire w2797;
	wire w2798;
	wire w2799;
	wire w2800;
	wire w2801;
	wire w2802;
	wire w2803;
	wire w2804;
	wire w2805;
	wire w2806;
	wire w2807;
	wire w2808;
	wire w2809;
	wire w2810;
	wire w2811;
	wire w2812;
	wire w2813;
	wire w2814;
	wire w2815;
	wire w2816;
	wire w2817;
	wire w2818;
	wire w2819;
	wire w2820;
	wire w2821;
	wire w2822;
	wire w2823;
	wire w2824;
	wire w2825;
	wire w2826;
	wire w2827;
	wire w2828;
	wire w2829;
	wire w2830;
	wire w2831;
	wire w2832;
	wire w2833;
	wire w2834;
	wire w2835;
	wire w2836;
	wire w2837;
	wire w2838;
	wire w2839;
	wire w2840;
	wire w2841;
	wire w2842;
	wire w2843;
	wire w2844;
	wire w2845;
	wire w2846;
	wire w2847;
	wire w2848;
	wire w2849;
	wire w2850;
	wire w2851;
	wire w2852;
	wire w2853;
	wire w2854;
	wire w2855;
	wire w2856;
	wire w2857;
	wire w2858;
	wire w2859;
	wire w2860;
	wire w2861;
	wire w2862;
	wire w2863;
	wire w2864;
	wire w2865;
	wire w2866;
	wire w2867;
	wire w2868;
	wire w2869;
	wire w2870;
	wire w2871;
	wire w2872;
	wire w2873;
	wire w2874;
	wire w2875;
	wire w2876;
	wire w2877;
	wire w2878;
	wire w2879;
	wire w2880;
	wire w2881;
	wire w2882;
	wire w2883;
	wire w2884;
	wire w2885;
	wire w2886;
	wire w2887;
	wire w2888;
	wire w2889;
	wire w2890;
	wire w2891;
	wire w2892;
	wire w2893;
	wire w2894;
	wire w2895;
	wire w2896;
	wire w2897;
	wire w2898;
	wire w2899;
	wire w2900;
	wire w2901;
	wire w2902;
	wire w2903;
	wire w2904;
	wire w2905;
	wire w2906;
	wire w2907;
	wire w2908;
	wire w2909;
	wire w2910;
	wire w2911;
	wire w2912;
	wire w2913;
	wire w2914;
	wire w2915;
	wire w2916;
	wire w2917;
	wire w2918;
	wire w2919;
	wire w2920;
	wire w2921;
	wire w2922;
	wire w2923;
	wire w2924;
	wire w2925;
	wire w2926;
	wire w2927;
	wire w2928;
	wire w2929;
	wire w2930;
	wire w2931;
	wire w2932;
	wire w2933;
	wire w2934;
	wire w2935;
	wire w2936;
	wire w2937;
	wire w2938;
	wire w2939;
	wire w2940;
	wire w2941;
	wire w2942;
	wire w2943;
	wire w2944;
	wire w2945;
	wire w2946;
	wire w2947;
	wire w2948;
	wire w2949;
	wire w2950;
	wire w2951;
	wire w2952;
	wire w2953;
	wire w2954;
	wire w2955;
	wire w2956;
	wire w2957;
	wire w2958;
	wire w2959;
	wire w2960;
	wire w2961;
	wire w2962;
	wire w2963;
	wire w2964;
	wire w2965;
	wire w2966;
	wire w2967;
	wire w2968;
	wire w2969;
	wire w2970;
	wire w2971;
	wire w2972;
	wire w2973;
	wire w2974;
	wire w2975;
	wire w2976;
	wire w2977;
	wire w2978;
	wire w2979;
	wire w2980;
	wire w2981;
	wire w2982;
	wire w2983;
	wire w2984;
	wire w2985;
	wire w2986;
	wire w2987;
	wire w2988;
	wire w2989;
	wire w2990;
	wire w2991;
	wire w2992;
	wire w2993;
	wire w2994;
	wire w2995;
	wire w2996;
	wire w2997;
	wire w2998;
	wire w2999;
	wire w3000;
	wire w3001;
	wire w3002;
	wire w3003;
	wire w3004;
	wire w3005;
	wire w3006;
	wire w3007;
	wire w3008;
	wire w3009;
	wire w3010;
	wire w3011;
	wire w3012;
	wire w3013;
	wire w3014;
	wire w3015;
	wire w3016;
	wire w3017;
	wire w3018;
	wire w3019;
	wire w3020;
	wire w3021;
	wire w3022;
	wire w3023;
	wire w3024;
	wire w3025;
	wire w3026;
	wire w3027;
	wire w3028;
	wire w3029;
	wire w3030;
	wire w3031;
	wire w3032;
	wire w3033;
	wire w3034;
	wire w3035;
	wire w3036;
	wire w3037;
	wire w3038;
	wire w3039;
	wire w3040;
	wire w3041;
	wire w3042;
	wire w3043;
	wire w3044;
	wire w3045;
	wire w3046;
	wire w3047;
	wire w3048;
	wire w3049;
	wire w3050;
	wire w3051;
	wire w3052;
	wire w3053;
	wire w3054;
	wire w3055;
	wire w3056;
	wire w3057;
	wire w3058;
	wire w3059;
	wire w3060;
	wire w3061;
	wire w3062;
	wire w3063;
	wire w3064;
	wire w3065;
	wire w3066;
	wire w3067;
	wire w3068;
	wire w3069;
	wire w3070;
	wire w3071;
	wire w3072;
	wire w3073;
	wire w3074;
	wire w3075;
	wire w3076;
	wire w3077;
	wire S[3];
	wire w3079;
	wire w3080;
	wire S[7];
	wire S[2];
	wire w3083;
	wire w3084;
	wire w3085;
	wire w3086;
	wire w3087;
	wire w3088;
	wire S[6];
	wire S[1];
	wire S[5];
	wire S[0];
	wire S[4];
	wire w3094;
	wire w3095;
	wire w3096;
	wire w3097;
	wire w3098;
	wire w3099;
	wire w3100;
	wire w3101;
	wire w3102;
	wire w3103;
	wire w3104;
	wire w3105;
	wire w3106;
	wire w3107;
	wire w3108;
	wire w3109;
	wire w3110;
	wire w3111;
	wire w3112;
	wire w3113;
	wire w3114;
	wire w3115;
	wire w3116;
	wire w3117;
	wire w3118;
	wire w3119;
	wire w3120;
	wire w3121;
	wire w3122;
	wire w3123;
	wire w3124;
	wire w3125;
	wire w3126;
	wire w3127;
	wire w3128;
	wire w3129;
	wire w3130;
	wire w3131;
	wire w3132;
	wire w3133;
	wire w3134;
	wire w3135;
	wire w3136;
	wire w3137;
	wire w3138;
	wire w3139;
	wire w3140;
	wire w3141;
	wire w3142;
	wire w3143;
	wire w3144;
	wire w3145;
	wire w3146;
	wire w3147;
	wire w3148;
	wire w3149;
	wire w3150;
	wire w3151;
	wire w3152;
	wire w3153;
	wire w3154;
	wire w3155;
	wire w3156;
	wire w3157;
	wire w3158;
	wire w3159;
	wire w3160;
	wire w3161;
	wire w3162;
	wire w3163;
	wire w3164;
	wire w3165;
	wire w3166;
	wire w3167;
	wire w3168;
	wire w3169;
	wire w3170;
	wire w3171;
	wire w3172;
	wire w3173;
	wire w3174;
	wire w3175;
	wire w3176;
	wire w3177;
	wire w3178;
	wire w3179;
	wire w3180;
	wire w3181;
	wire w3182;
	wire w3183;
	wire w3184;
	wire w3185;
	wire w3186;
	wire w3187;
	wire w3188;
	wire w3189;
	wire w3190;
	wire w3191;
	wire w3192;
	wire w3193;
	wire w3194;
	wire w3195;
	wire w3196;
	wire w3197;
	wire w3198;
	wire w3199;
	wire w3200;
	wire w3201;
	wire w3202;
	wire w3203;
	wire w3204;
	wire w3205;
	wire w3206;
	wire w3207;
	wire w3208;
	wire w3209;
	wire w3210;
	wire w3211;
	wire w3212;
	wire w3213;
	wire w3214;
	wire w3215;
	wire w3216;
	wire w3217;
	wire w3218;
	wire w3219;
	wire w3220;
	wire w3221;
	wire w3222;
	wire w3223;
	wire w3224;
	wire w3225;
	wire w3226;
	wire w3227;
	wire w3228;
	wire w3229;
	wire w3230;
	wire w3231;
	wire w3232;
	wire w3233;
	wire w3234;
	wire w3235;
	wire w3236;
	wire w3237;
	wire w3238;
	wire w3239;
	wire w3240;
	wire w3241;
	wire w3242;
	wire w3243;
	wire w3244;
	wire w3245;
	wire w3246;
	wire w3247;
	wire w3248;
	wire w3249;
	wire w3250;
	wire w3251;
	wire w3252;
	wire w3253;
	wire w3254;
	wire w3255;
	wire w3256;
	wire w3257;
	wire w3258;
	wire w3259;
	wire w3260;
	wire w3261;
	wire w3262;
	wire w3263;
	wire w3264;
	wire w3265;
	wire w3266;
	wire w3267;
	wire w3268;
	wire w3269;
	wire w3270;
	wire w3271;
	wire w3272;
	wire w3273;
	wire w3274;
	wire w3275;
	wire w3276;
	wire w3277;
	wire w3278;
	wire w3279;
	wire w3280;
	wire w3281;
	wire w3282;
	wire w3283;
	wire w3284;
	wire w3285;
	wire w3286;
	wire w3287;
	wire w3288;
	wire w3289;
	wire w3290;
	wire w3291;
	wire w3292;
	wire w3293;
	wire w3294;
	wire w3295;
	wire w3296;
	wire w3297;
	wire w3298;
	wire w3299;
	wire w3300;
	wire w3301;
	wire w3302;
	wire w3303;
	wire w3304;
	wire w3305;
	wire w3306;
	wire w3307;
	wire w3308;
	wire w3309;
	wire w3310;
	wire w3311;
	wire w3312;
	wire w3313;
	wire w3314;
	wire w3315;
	wire w3316;
	wire w3317;
	wire w3318;
	wire w3319;
	wire w3320;
	wire w3321;
	wire w3322;
	wire w3323;
	wire w3324;
	wire w3325;
	wire w3326;
	wire w3327;
	wire w3328;
	wire w3329;
	wire w3330;
	wire w3331;
	wire w3332;
	wire w3333;
	wire w3334;
	wire w3335;
	wire w3336;
	wire w3337;
	wire w3338;
	wire w3339;
	wire w3340;
	wire w3341;
	wire w3342;
	wire w3343;
	wire w3344;
	wire w3345;
	wire w3346;
	wire w3347;
	wire w3348;
	wire w3349;
	wire w3350;
	wire w3351;
	wire w3352;
	wire w3353;
	wire w3354;
	wire w3355;
	wire w3356;
	wire w3357;
	wire w3358;
	wire w3359;
	wire w3360;
	wire w3361;
	wire w3362;
	wire w3363;
	wire w3364;
	wire w3365;
	wire w3366;
	wire w3367;
	wire w3368;
	wire w3369;
	wire w3370;
	wire w3371;
	wire w3372;
	wire w3373;
	wire w3374;
	wire w3375;
	wire w3376;
	wire w3377;
	wire w3378;
	wire w3379;
	wire w3380;
	wire w3381;
	wire w3382;
	wire w3383;
	wire w3384;
	wire w3385;
	wire w3386;
	wire w3387;
	wire w3388;
	wire w3389;
	wire w3390;
	wire w3391;
	wire w3392;
	wire w3393;
	wire w3394;
	wire w3395;
	wire w3396;
	wire w3397;
	wire w3398;
	wire w3399;
	wire w3400;
	wire w3401;
	wire w3402;
	wire w3403;
	wire w3404;
	wire w3405;
	wire w3406;
	wire w3407;
	wire w3408;
	wire w3409;
	wire w3410;
	wire w3411;
	wire w3412;
	wire w3413;
	wire w3414;
	wire w3415;
	wire w3416;
	wire w3417;
	wire w3418;
	wire w3419;
	wire w3420;
	wire w3421;
	wire w3422;
	wire w3423;
	wire w3424;
	wire w3425;
	wire w3426;
	wire w3427;
	wire w3428;
	wire w3429;
	wire w3430;
	wire w3431;
	wire w3432;
	wire w3433;
	wire w3434;
	wire w3435;
	wire w3436;
	wire w3437;
	wire w3438;
	wire w3439;
	wire w3440;
	wire w3441;
	wire w3442;
	wire w3443;
	wire w3444;
	wire w3445;
	wire w3446;
	wire w3447;
	wire w3448;
	wire w3449;
	wire w3450;
	wire w3451;
	wire w3452;
	wire w3453;
	wire w3454;
	wire w3455;
	wire w3456;
	wire w3457;
	wire w3458;
	wire w3459;
	wire w3460;
	wire w3461;
	wire w3462;
	wire w3463;
	wire w3464;
	wire w3465;
	wire w3466;
	wire w3467;
	wire w3468;
	wire w3469;
	wire w3470;
	wire w3471;
	wire w3472;
	wire w3473;
	wire w3474;
	wire w3475;
	wire w3476;
	wire w3477;
	wire w3478;
	wire w3479;
	wire w3480;
	wire w3481;
	wire w3482;
	wire w3483;
	wire w3484;
	wire w3485;
	wire w3486;
	wire w3487;
	wire w3488;
	wire w3489;
	wire w3490;
	wire w3491;
	wire w3492;
	wire w3493;
	wire w3494;
	wire w3495;
	wire w3496;
	wire w3497;
	wire w3498;
	wire w3499;
	wire w3500;
	wire w3501;
	wire w3502;
	wire w3503;
	wire w3504;
	wire w3505;
	wire w3506;
	wire w3507;
	wire w3508;
	wire w3509;
	wire w3510;
	wire w3511;
	wire w3512;
	wire w3513;
	wire w3514;
	wire w3515;
	wire w3516;
	wire w3517;
	wire w3518;
	wire w3519;
	wire w3520;
	wire w3521;
	wire w3522;
	wire w3523;
	wire w3524;
	wire w3525;
	wire w3526;
	wire w3527;
	wire w3528;
	wire w3529;
	wire w3530;
	wire w3531;
	wire w3532;
	wire w3533;
	wire w3534;
	wire w3535;
	wire w3536;
	wire w3537;
	wire w3538;
	wire w3539;
	wire w3540;
	wire w3541;
	wire w3542;
	wire w3543;
	wire w3544;
	wire w3545;
	wire w3546;
	wire w3547;
	wire w3548;
	wire w3549;
	wire w3550;
	wire w3551;
	wire w3552;
	wire w3553;
	wire w3554;
	wire w3555;
	wire w3556;
	wire w3557;
	wire w3558;
	wire w3559;
	wire w3560;
	wire w3561;
	wire w3562;
	wire w3563;
	wire w3564;
	wire w3565;
	wire w3566;
	wire w3567;
	wire w3568;
	wire w3569;
	wire w3570;
	wire w3571;
	wire w3572;
	wire w3573;
	wire w3574;
	wire w3575;
	wire w3576;
	wire w3577;
	wire w3578;
	wire w3579;
	wire w3580;
	wire w3581;
	wire w3582;
	wire w3583;
	wire w3584;
	wire w3585;
	wire w3586;
	wire w3587;
	wire w3588;
	wire w3589;
	wire w3590;
	wire w3591;
	wire w3592;
	wire w3593;
	wire w3594;
	wire w3595;
	wire w3596;
	wire w3597;
	wire w3598;
	wire w3599;
	wire w3600;
	wire w3601;
	wire w3602;
	wire w3603;
	wire w3604;
	wire w3605;
	wire w3606;
	wire w3607;
	wire w3608;
	wire w3609;
	wire w3610;
	wire w3611;
	wire w3612;
	wire w3613;
	wire w3614;
	wire w3615;
	wire w3616;
	wire w3617;
	wire w3618;
	wire w3619;
	wire w3620;
	wire w3621;
	wire w3622;
	wire w3623;
	wire w3624;
	wire w3625;
	wire w3626;
	wire w3627;
	wire w3628;
	wire w3629;
	wire w3630;
	wire w3631;
	wire w3632;
	wire w3633;
	wire w3634;
	wire w3635;
	wire w3636;
	wire w3637;
	wire w3638;
	wire w3639;
	wire w3640;
	wire w3641;
	wire w3642;
	wire w3643;
	wire w3644;
	wire w3645;
	wire w3646;
	wire w3647;
	wire w3648;
	wire w3649;
	wire w3650;
	wire w3651;
	wire w3652;
	wire w3653;
	wire w3654;
	wire w3655;
	wire w3656;
	wire w3657;
	wire w3658;
	wire w3659;
	wire w3660;
	wire w3661;
	wire w3662;
	wire w3663;
	wire w3664;
	wire w3665;
	wire w3666;
	wire w3667;
	wire w3668;
	wire w3669;
	wire w3670;
	wire w3671;
	wire w3672;
	wire w3673;
	wire w3674;
	wire w3675;
	wire w3676;
	wire w3677;
	wire w3678;
	wire w3679;
	wire w3680;
	wire w3681;
	wire w3682;
	wire w3683;
	wire w3684;
	wire w3685;
	wire w3686;
	wire w3687;
	wire w3688;
	wire w3689;
	wire w3690;
	wire w3691;
	wire w3692;
	wire w3693;
	wire w3694;
	wire w3695;
	wire w3696;
	wire w3697;
	wire w3698;
	wire w3699;
	wire w3700;
	wire w3701;
	wire w3702;
	wire w3703;
	wire w3704;
	wire w3705;
	wire w3706;
	wire w3707;
	wire w3708;
	wire w3709;
	wire w3710;
	wire w3711;
	wire w3712;
	wire w3713;
	wire w3714;
	wire w3715;
	wire w3716;
	wire w3717;
	wire w3718;
	wire w3719;
	wire w3720;
	wire w3721;
	wire w3722;
	wire w3723;
	wire w3724;
	wire w3725;
	wire w3726;
	wire w3727;
	wire w3728;
	wire w3729;
	wire w3730;
	wire w3731;
	wire w3732;
	wire w3733;
	wire w3734;
	wire w3735;
	wire w3736;
	wire w3737;
	wire w3738;
	wire w3739;
	wire w3740;
	wire w3741;
	wire w3742;
	wire w3743;
	wire w3744;
	wire w3745;
	wire w3746;
	wire w3747;
	wire w3748;
	wire w3749;
	wire w3750;
	wire w3751;
	wire w3752;
	wire w3753;
	wire w3754;
	wire w3755;
	wire w3756;
	wire w3757;
	wire w3758;
	wire w3759;
	wire w3760;
	wire w3761;
	wire w3762;
	wire w3763;
	wire w3764;
	wire w3765;
	wire w3766;
	wire w3767;
	wire w3768;
	wire w3769;
	wire w3770;
	wire w3771;
	wire w3772;
	wire w3773;
	wire w3774;
	wire w3775;
	wire w3776;
	wire w3777;
	wire w3778;
	wire w3779;
	wire w3780;
	wire w3781;
	wire w3782;
	wire w3783;
	wire w3784;
	wire w3785;
	wire w3786;
	wire w3787;
	wire w3788;
	wire w3789;
	wire w3790;
	wire w3791;
	wire w3792;
	wire w3793;
	wire w3794;
	wire w3795;
	wire w3796;
	wire w3797;
	wire w3798;
	wire w3799;
	wire w3800;
	wire w3801;
	wire w3802;
	wire w3803;
	wire w3804;
	wire w3805;
	wire w3806;
	wire w3807;
	wire w3808;
	wire w3809;
	wire w3810;
	wire w3811;
	wire w3812;
	wire w3813;
	wire w3814;
	wire w3815;
	wire w3816;
	wire w3817;
	wire w3818;
	wire w3819;
	wire w3820;
	wire w3821;
	wire w3822;
	wire w3823;
	wire w3824;
	wire w3825;
	wire w3826;
	wire w3827;
	wire w3828;
	wire w3829;
	wire w3830;
	wire w3831;
	wire w3832;
	wire w3833;
	wire w3834;
	wire w3835;
	wire w3836;
	wire w3837;
	wire w3838;
	wire w3839;
	wire w3840;
	wire w3841;
	wire w3842;
	wire w3843;
	wire w3844;
	wire w3845;
	wire w3846;
	wire w3847;
	wire w3848;
	wire w3849;
	wire w3850;
	wire w3851;
	wire w3852;
	wire w3853;
	wire w3854;
	wire w3855;
	wire w3856;
	wire w3857;
	wire w3858;
	wire w3859;
	wire w3860;
	wire w3861;
	wire w3862;
	wire w3863;
	wire w3864;
	wire w3865;
	wire w3866;
	wire w3867;
	wire w3868;
	wire w3869;
	wire w3870;
	wire w3871;
	wire w3872;
	wire w3873;
	wire w3874;
	wire w3875;
	wire w3876;
	wire w3877;
	wire w3878;
	wire w3879;
	wire w3880;
	wire w3881;
	wire w3882;
	wire w3883;
	wire w3884;
	wire w3885;
	wire w3886;
	wire w3887;
	wire w3888;
	wire w3889;
	wire w3890;
	wire w3891;
	wire w3892;
	wire w3893;
	wire w3894;
	wire w3895;
	wire w3896;
	wire w3897;
	wire w3898;
	wire w3899;
	wire w3900;
	wire w3901;
	wire w3902;
	wire w3903;
	wire w3904;
	wire w3905;
	wire w3906;
	wire w3907;
	wire w3908;
	wire w3909;
	wire w3910;
	wire w3911;
	wire w3912;
	wire w3913;
	wire w3914;
	wire w3915;
	wire w3916;
	wire w3917;
	wire w3918;
	wire w3919;
	wire w3920;
	wire w3921;
	wire w3922;
	wire w3923;
	wire w3924;
	wire w3925;
	wire w3926;
	wire w3927;
	wire w3928;
	wire w3929;
	wire w3930;
	wire w3931;
	wire w3932;
	wire w3933;
	wire w3934;
	wire w3935;
	wire w3936;
	wire w3937;
	wire w3938;
	wire w3939;
	wire w3940;
	wire w3941;
	wire w3942;
	wire w3943;
	wire w3944;
	wire w3945;
	wire w3946;
	wire w3947;
	wire w3948;
	wire w3949;
	wire w3950;
	wire w3951;
	wire w3952;
	wire w3953;
	wire w3954;
	wire w3955;
	wire w3956;
	wire w3957;
	wire w3958;
	wire w3959;
	wire w3960;
	wire w3961;
	wire w3962;
	wire w3963;
	wire w3964;
	wire w3965;
	wire w3966;
	wire w3967;
	wire w3968;
	wire w3969;
	wire w3970;
	wire w3971;
	wire w3972;
	wire w3973;
	wire w3974;
	wire w3975;
	wire w3976;
	wire w3977;
	wire w3978;
	wire w3979;
	wire w3980;
	wire w3981;
	wire w3982;
	wire w3983;
	wire w3984;
	wire w3985;
	wire w3986;
	wire w3987;
	wire w3988;
	wire w3989;
	wire w3990;
	wire w3991;
	wire w3992;
	wire w3993;
	wire w3994;
	wire w3995;
	wire w3996;
	wire w3997;
	wire w3998;
	wire w3999;
	wire w4000;
	wire w4001;
	wire w4002;
	wire w4003;
	wire w4004;
	wire w4005;
	wire w4006;
	wire w4007;
	wire w4008;
	wire w4009;
	wire w4010;
	wire w4011;
	wire w4012;
	wire w4013;
	wire w4014;
	wire w4015;
	wire w4016;
	wire w4017;
	wire w4018;
	wire w4019;
	wire w4020;
	wire w4021;
	wire w4022;
	wire w4023;
	wire w4024;
	wire w4025;
	wire w4026;
	wire w4027;
	wire w4028;
	wire w4029;
	wire w4030;
	wire w4031;
	wire w4032;
	wire w4033;
	wire w4034;
	wire w4035;
	wire w4036;
	wire w4037;
	wire w4038;
	wire w4039;
	wire w4040;
	wire w4041;
	wire w4042;
	wire w4043;
	wire w4044;
	wire w4045;
	wire w4046;
	wire w4047;
	wire w4048;
	wire w4049;
	wire w4050;
	wire w4051;
	wire w4052;
	wire w4053;
	wire w4054;
	wire w4055;
	wire w4056;
	wire w4057;
	wire w4058;
	wire w4059;
	wire w4060;
	wire w4061;
	wire w4062;
	wire w4063;
	wire w4064;
	wire w4065;
	wire w4066;
	wire w4067;
	wire w4068;
	wire w4069;
	wire w4070;
	wire w4071;
	wire w4072;
	wire w4073;
	wire w4074;
	wire w4075;
	wire w4076;
	wire w4077;
	wire w4078;
	wire w4079;
	wire w4080;
	wire w4081;
	wire w4082;
	wire w4083;
	wire w4084;
	wire w4085;
	wire w4086;
	wire w4087;
	wire w4088;
	wire w4089;
	wire w4090;
	wire w4091;
	wire w4092;
	wire w4093;
	wire w4094;
	wire w4095;
	wire w4096;
	wire w4097;
	wire w4098;
	wire w4099;
	wire w4100;
	wire w4101;
	wire w4102;
	wire w4103;
	wire w4104;
	wire w4105;
	wire w4106;
	wire w4107;
	wire w4108;
	wire w4109;
	wire w4110;
	wire w4111;
	wire w4112;
	wire w4113;
	wire w4114;
	wire w4115;
	wire w4116;
	wire w4117;
	wire w4118;
	wire w4119;
	wire w4120;
	wire w4121;
	wire w4122;
	wire w4123;
	wire w4124;
	wire w4125;
	wire w4126;
	wire w4127;
	wire w4128;
	wire w4129;
	wire w4130;
	wire w4131;
	wire w4132;
	wire w4133;
	wire w4134;
	wire w4135;
	wire w4136;
	wire w4137;
	wire w4138;
	wire w4139;
	wire w4140;
	wire w4141;
	wire w4142;
	wire w4143;
	wire w4144;
	wire w4145;
	wire w4146;
	wire w4147;
	wire w4148;
	wire w4149;
	wire w4150;
	wire w4151;
	wire w4152;
	wire w4153;
	wire w4154;
	wire w4155;
	wire w4156;
	wire w4157;
	wire w4158;
	wire w4159;
	wire w4160;
	wire w4161;
	wire w4162;
	wire w4163;
	wire w4164;
	wire w4165;
	wire w4166;
	wire w4167;
	wire w4168;
	wire w4169;
	wire w4170;
	wire w4171;
	wire w4172;
	wire w4173;
	wire w4174;
	wire w4175;
	wire w4176;
	wire w4177;
	wire w4178;
	wire w4179;
	wire w4180;
	wire w4181;
	wire w4182;
	wire w4183;
	wire w4184;
	wire w4185;
	wire w4186;
	wire w4187;
	wire w4188;
	wire w4189;
	wire w4190;
	wire w4191;
	wire w4192;
	wire w4193;
	wire w4194;
	wire w4195;
	wire w4196;
	wire w4197;
	wire w4198;
	wire w4199;
	wire w4200;
	wire w4201;
	wire w4202;
	wire w4203;
	wire w4204;
	wire w4205;
	wire w4206;
	wire w4207;
	wire w4208;
	wire w4209;
	wire w4210;
	wire w4211;
	wire w4212;
	wire w4213;
	wire w4214;
	wire w4215;
	wire w4216;
	wire w4217;
	wire w4218;
	wire w4219;
	wire w4220;
	wire w4221;
	wire w4222;
	wire w4223;
	wire w4224;
	wire w4225;
	wire w4226;
	wire w4227;
	wire w4228;
	wire w4229;
	wire w4230;
	wire w4231;
	wire w4232;
	wire w4233;
	wire w4234;
	wire w4235;
	wire w4236;
	wire w4237;
	wire w4238;
	wire w4239;
	wire w4240;
	wire w4241;
	wire w4242;
	wire w4243;
	wire w4244;
	wire w4245;
	wire w4246;
	wire w4247;
	wire w4248;
	wire w4249;
	wire w4250;
	wire w4251;
	wire w4252;
	wire w4253;
	wire w4254;
	wire w4255;
	wire w4256;
	wire w4257;
	wire w4258;
	wire w4259;
	wire w4260;
	wire w4261;
	wire w4262;
	wire w4263;
	wire w4264;
	wire w4265;
	wire w4266;
	wire w4267;
	wire w4268;
	wire w4269;
	wire w4270;
	wire w4271;
	wire w4272;
	wire w4273;
	wire w4274;
	wire w4275;
	wire w4276;
	wire w4277;
	wire w4278;
	wire w4279;
	wire w4280;
	wire w4281;
	wire w4282;
	wire w4283;
	wire w4284;
	wire w4285;
	wire w4286;
	wire w4287;
	wire w4288;
	wire w4289;
	wire w4290;
	wire w4291;
	wire w4292;
	wire w4293;
	wire w4294;
	wire w4295;
	wire w4296;
	wire w4297;
	wire w4298;
	wire w4299;
	wire w4300;
	wire w4301;
	wire w4302;
	wire w4303;
	wire w4304;
	wire w4305;
	wire w4306;
	wire w4307;
	wire w4308;
	wire w4309;
	wire w4310;
	wire w4311;
	wire w4312;
	wire w4313;
	wire w4314;
	wire w4315;
	wire w4316;
	wire w4317;
	wire w4318;
	wire w4319;
	wire w4320;
	wire w4321;
	wire w4322;
	wire w4323;
	wire w4324;
	wire w4325;
	wire w4326;
	wire w4327;
	wire w4328;
	wire w4329;
	wire w4330;
	wire w4331;
	wire w4332;
	wire w4333;
	wire w4334;
	wire w4335;
	wire w4336;
	wire w4337;
	wire w4338;
	wire w4339;
	wire w4340;
	wire w4341;
	wire w4342;
	wire w4343;
	wire w4344;
	wire w4345;
	wire w4346;
	wire w4347;
	wire w4348;
	wire w4349;
	wire w4350;
	wire w4351;
	wire w4352;
	wire w4353;
	wire w4354;
	wire w4355;
	wire w4356;
	wire w4357;
	wire w4358;
	wire w4359;
	wire w4360;
	wire w4361;
	wire w4362;
	wire w4363;
	wire w4364;
	wire w4365;
	wire w4366;
	wire w4367;
	wire w4368;
	wire w4369;
	wire w4370;
	wire w4371;
	wire w4372;
	wire w4373;
	wire w4374;
	wire w4375;
	wire w4376;
	wire w4377;
	wire w4378;
	wire w4379;
	wire w4380;
	wire w4381;
	wire w4382;
	wire w4383;
	wire w4384;
	wire w4385;
	wire w4386;
	wire w4387;
	wire w4388;
	wire w4389;
	wire w4390;
	wire w4391;
	wire w4392;
	wire w4393;
	wire w4394;
	wire w4395;
	wire w4396;
	wire w4397;
	wire w4398;
	wire w4399;
	wire w4400;
	wire w4401;
	wire w4402;
	wire w4403;
	wire w4404;
	wire w4405;
	wire w4406;
	wire w4407;
	wire w4408;
	wire w4409;
	wire w4410;
	wire w4411;
	wire w4412;
	wire w4413;
	wire w4414;
	wire w4415;
	wire w4416;
	wire w4417;
	wire w4418;
	wire w4419;
	wire w4420;
	wire w4421;
	wire w4422;
	wire w4423;
	wire w4424;
	wire w4425;
	wire w4426;
	wire w4427;
	wire w4428;
	wire w4429;
	wire w4430;
	wire w4431;
	wire w4432;
	wire w4433;
	wire w4434;
	wire w4435;
	wire w4436;
	wire w4437;
	wire w4438;
	wire w4439;
	wire w4440;
	wire w4441;
	wire w4442;
	wire w4443;
	wire w4444;
	wire w4445;
	wire w4446;
	wire w4447;
	wire w4448;
	wire w4449;
	wire w4450;
	wire w4451;
	wire w4452;
	wire w4453;
	wire w4454;
	wire w4455;
	wire w4456;
	wire w4457;
	wire w4458;
	wire w4459;
	wire w4460;
	wire w4461;
	wire w4462;
	wire w4463;
	wire w4464;
	wire w4465;
	wire w4466;
	wire w4467;
	wire w4468;
	wire w4469;
	wire w4470;
	wire w4471;
	wire w4472;
	wire w4473;
	wire w4474;
	wire 68K CPU CLOCK;
	wire w4476;
	wire w4477;
	wire w4478;
	wire w4479;
	wire w4480;
	wire w4481;
	wire w4482;
	wire w4483;
	wire w4484;
	wire w4485;
	wire w4486;
	wire w4487;
	wire w4488;
	wire w4489;
	wire w4490;
	wire w4491;
	wire w4492;
	wire w4493;
	wire w4494;
	wire w4495;
	wire w4496;
	wire w4497;
	wire w4498;
	wire w4499;
	wire w4500;
	wire w4501;
	wire w4502;
	wire w4503;
	wire w4504;
	wire w4505;
	wire w4506;
	wire w4507;
	wire w4508;
	wire w4509;
	wire w4510;
	wire w4511;
	wire w4512;
	wire w4513;
	wire w4514;
	wire w4515;
	wire w4516;
	wire w4517;
	wire w4518;
	wire w4519;
	wire nRAS1;
	wire nCAS1;
	wire nWE1;
	wire nWE0;
	wire nOE1;
	wire AD_RD_DIR;
	wire w4526;
	wire w4527;
	wire w4528;
	wire w4529;
	wire w4530;
	wire w4531;
	wire w4532;
	wire w4533;
	wire w4534;
	wire w4535;
	wire w4536;
	wire w4537;
	wire w4538;
	wire w4539;
	wire w4540;
	wire w4541;
	wire w4542;
	wire w4543;
	wire w4544;
	wire w4545;
	wire w4546;
	wire w4547;
	wire w4548;
	wire w4549;
	wire w4550;
	wire w4551;
	wire w4552;
	wire w4553;
	wire w4554;
	wire w4555;
	wire w4556;
	wire w4557;
	wire w4558;
	wire w4559;
	wire w4560;
	wire w4561;
	wire w4562;
	wire w4563;
	wire w4564;
	wire w4565;
	wire w4566;
	wire w4567;
	wire w4568;
	wire w4569;
	wire w4570;
	wire w4571;
	wire w4572;
	wire w4573;
	wire w4574;
	wire w4575;
	wire w4576;
	wire w4577;
	wire w4578;
	wire w4579;
	wire w4580;
	wire w4581;
	wire w4582;
	wire w4583;
	wire w4584;
	wire w4585;
	wire w4586;
	wire w4587;
	wire w4588;
	wire w4589;
	wire w4590;
	wire w4591;
	wire w4592;
	wire w4593;
	wire w4594;
	wire w4595;
	wire w4596;
	wire w4597;
	wire w4598;
	wire w4599;
	wire w4600;
	wire w4601;
	wire w4602;
	wire w4603;
	wire w4604;
	wire w4605;
	wire w4606;
	wire w4607;
	wire w4608;
	wire w4609;
	wire w4610;
	wire w4611;
	wire w4612;
	wire w4613;
	wire w4614;
	wire w4615;
	wire w4616;
	wire w4617;
	wire w4618;
	wire w4619;
	wire w4620;
	wire w4621;
	wire w4622;
	wire w4623;
	wire w4624;
	wire w4625;
	wire w4626;
	wire w4627;
	wire w4628;
	wire w4629;
	wire w4630;
	wire w4631;
	wire w4632;
	wire w4633;
	wire w4634;
	wire w4635;
	wire w4636;
	wire w4637;
	wire w4638;
	wire w4639;
	wire w4640;
	wire w4641;
	wire w4642;
	wire w4643;
	wire w4644;
	wire w4645;
	wire w4646;
	wire w4647;
	wire w4648;
	wire w4649;
	wire w4650;
	wire w4651;
	wire w4652;
	wire w4653;
	wire w4654;
	wire w4655;
	wire w4656;
	wire w4657;
	wire w4658;
	wire w4659;
	wire w4660;
	wire w4661;
	wire w4662;
	wire w4663;
	wire w4664;
	wire w4665;
	wire w4666;
	wire w4667;
	wire w4668;
	wire w4669;
	wire w4670;
	wire w4671;
	wire w4672;
	wire w4673;
	wire w4674;
	wire w4675;
	wire w4676;
	wire w4677;
	wire w4678;
	wire w4679;
	wire w4680;
	wire w4681;
	wire w4682;
	wire w4683;
	wire w4684;
	wire w4685;
	wire w4686;
	wire w4687;
	wire w4688;
	wire w4689;
	wire w4690;
	wire w4691;
	wire w4692;
	wire w4693;
	wire w4694;
	wire w4695;
	wire w4696;
	wire w4697;
	wire w4698;
	wire w4699;
	wire w4700;
	wire w4701;
	wire w4702;
	wire w4703;
	wire w4704;
	wire w4705;
	wire w4706;
	wire w4707;
	wire w4708;
	wire w4709;
	wire w4710;
	wire w4711;
	wire w4712;
	wire w4713;
	wire w4714;
	wire w4715;
	wire w4716;
	wire w4717;
	wire w4718;
	wire w4719;
	wire w4720;
	wire w4721;
	wire w4722;
	wire w4723;
	wire w4724;
	wire w4725;
	wire w4726;
	wire w4727;
	wire w4728;
	wire w4729;
	wire w4730;
	wire w4731;
	wire w4732;
	wire w4733;
	wire w4734;
	wire w4735;
	wire w4736;
	wire w4737;
	wire w4738;
	wire w4739;
	wire w4740;
	wire w4741;
	wire w4742;
	wire w4743;
	wire w4744;
	wire w4745;
	wire w4746;
	wire w4747;
	wire w4748;
	wire w4749;
	wire w4750;
	wire w4751;
	wire w4752;
	wire w4753;
	wire w4754;
	wire w4755;
	wire w4756;
	wire w4757;
	wire w4758;
	wire w4759;
	wire w4760;
	wire w4761;
	wire w4762;
	wire w4763;
	wire w4764;
	wire w4765;
	wire w4766;
	wire w4767;
	wire w4768;
	wire w4769;
	wire w4770;
	wire w4771;
	wire w4772;
	wire w4773;
	wire w4774;
	wire w4775;
	wire w4776;
	wire w4777;
	wire w4778;
	wire w4779;
	wire w4780;
	wire w4781;
	wire w4782;
	wire w4783;
	wire w4784;
	wire w4785;
	wire w4786;
	wire w4787;
	wire w4788;
	wire w4789;
	wire w4790;
	wire w4791;
	wire w4792;
	wire w4793;
	wire w4794;
	wire w4795;
	wire w4796;
	wire w4797;
	wire w4798;
	wire w4799;
	wire w4800;
	wire w4801;
	wire w4802;
	wire w4803;
	wire w4804;
	wire w4805;
	wire w4806;
	wire w4807;
	wire w4808;
	wire w4809;
	wire w4810;
	wire w4811;
	wire w4812;
	wire w4813;
	wire w4814;
	wire w4815;
	wire w4816;
	wire w4817;
	wire w4818;
	wire w4819;
	wire w4820;
	wire w4821;
	wire w4822;
	wire w4823;
	wire w4824;
	wire w4825;
	wire w4826;
	wire w4827;
	wire w4828;
	wire w4829;
	wire w4830;
	wire w4831;
	wire w4832;
	wire w4833;
	wire w4834;
	wire w4835;
	wire w4836;
	wire w4837;
	wire w4838;
	wire w4839;
	wire w4840;
	wire w4841;
	wire w4842;
	wire w4843;
	wire w4844;
	wire w4845;
	wire w4846;
	wire w4847;
	wire w4848;
	wire w4849;
	wire w4850;
	wire w4851;
	wire w4852;
	wire w4853;
	wire w4854;
	wire w4855;
	wire w4856;
	wire w4857;
	wire w4858;
	wire w4859;
	wire w4860;
	wire w4861;
	wire w4862;
	wire w4863;
	wire w4864;
	wire w4865;
	wire w4866;
	wire w4867;
	wire w4868;
	wire w4869;
	wire w4870;
	wire w4871;
	wire w4872;
	wire w4873;
	wire w4874;
	wire w4875;
	wire w4876;
	wire w4877;
	wire w4878;
	wire w4879;
	wire w4880;
	wire w4881;
	wire w4882;
	wire w4883;
	wire w4884;
	wire w4885;
	wire w4886;
	wire w4887;
	wire w4888;
	wire w4889;
	wire w4890;
	wire w4891;
	wire w4892;
	wire w4893;
	wire w4894;
	wire w4895;
	wire w4896;
	wire w4897;
	wire w4898;
	wire w4899;
	wire w4900;
	wire w4901;
	wire w4902;
	wire w4903;
	wire w4904;
	wire w4905;
	wire w4906;
	wire w4907;
	wire w4908;
	wire w4909;
	wire w4910;
	wire w4911;
	wire w4912;
	wire w4913;
	wire w4914;
	wire w4915;
	wire w4916;
	wire w4917;
	wire w4918;
	wire w4919;
	wire w4920;
	wire w4921;
	wire w4922;
	wire w4923;
	wire w4924;
	wire w4925;
	wire w4926;
	wire w4927;
	wire w4928;
	wire w4929;
	wire w4930;
	wire w4931;
	wire w4932;
	wire w4933;
	wire w4934;
	wire w4935;
	wire w4936;
	wire w4937;
	wire w4938;
	wire w4939;
	wire w4940;
	wire w4941;
	wire w4942;
	wire w4943;
	wire w4944;
	wire w4945;
	wire w4946;
	wire w4947;
	wire w4948;
	wire w4949;
	wire w4950;
	wire w4951;
	wire w4952;
	wire w4953;
	wire w4954;
	wire w4955;
	wire w4956;
	wire w4957;
	wire w4958;
	wire w4959;
	wire w4960;
	wire w4961;
	wire w4962;
	wire w4963;
	wire w4964;
	wire w4965;
	wire w4966;
	wire w4967;
	wire w4968;
	wire w4969;
	wire w4970;
	wire w4971;
	wire w4972;
	wire w4973;
	wire w4974;
	wire w4975;
	wire w4976;
	wire w4977;
	wire w4978;
	wire w4979;
	wire w4980;
	wire w4981;
	wire w4982;
	wire w4983;
	wire w4984;
	wire w4985;
	wire w4986;
	wire w4987;
	wire w4988;
	wire w4989;
	wire w4990;
	wire w4991;
	wire w4992;
	wire w4993;
	wire w4994;
	wire w4995;
	wire w4996;
	wire w4997;
	wire w4998;
	wire w4999;
	wire w5000;
	wire w5001;
	wire w5002;
	wire w5003;
	wire w5004;
	wire w5005;
	wire w5006;
	wire w5007;
	wire w5008;
	wire w5009;
	wire w5010;
	wire w5011;
	wire w5012;
	wire w5013;
	wire w5014;
	wire w5015;
	wire w5016;
	wire w5017;
	wire w5018;
	wire w5019;
	wire w5020;
	wire w5021;
	wire w5022;
	wire w5023;
	wire w5024;
	wire w5025;
	wire w5026;
	wire w5027;
	wire w5028;
	wire w5029;
	wire w5030;
	wire w5031;
	wire w5032;
	wire w5033;
	wire w5034;
	wire w5035;
	wire w5036;
	wire w5037;
	wire w5038;
	wire w5039;
	wire w5040;
	wire w5041;
	wire w5042;
	wire w5043;
	wire w5044;
	wire w5045;
	wire w5046;
	wire w5047;
	wire w5048;
	wire w5049;
	wire w5050;
	wire w5051;
	wire w5052;
	wire w5053;
	wire w5054;
	wire w5055;
	wire w5056;
	wire w5057;
	wire w5058;
	wire w5059;
	wire w5060;
	wire w5061;
	wire w5062;
	wire w5063;
	wire w5064;
	wire w5065;
	wire w5066;
	wire w5067;
	wire w5068;
	wire w5069;
	wire w5070;
	wire w5071;
	wire w5072;
	wire w5073;
	wire w5074;
	wire w5075;
	wire w5076;
	wire w5077;
	wire w5078;
	wire w5079;
	wire w5080;
	wire w5081;
	wire w5082;
	wire w5083;
	wire w5084;
	wire w5085;
	wire w5086;
	wire w5087;
	wire w5088;
	wire w5089;
	wire w5090;
	wire w5091;
	wire w5092;
	wire w5093;
	wire w5094;
	wire w5095;
	wire w5096;
	wire w5097;
	wire w5098;
	wire w5099;
	wire w5100;
	wire w5101;
	wire w5102;
	wire w5103;
	wire w5104;
	wire w5105;
	wire w5106;
	wire w5107;
	wire w5108;
	wire w5109;
	wire w5110;
	wire w5111;
	wire w5112;
	wire w5113;
	wire w5114;
	wire w5115;
	wire w5116;
	wire w5117;
	wire w5118;
	wire w5119;
	wire w5120;
	wire w5121;
	wire w5122;
	wire w5123;
	wire w5124;
	wire w5125;
	wire w5126;
	wire w5127;
	wire w5128;
	wire w5129;
	wire w5130;
	wire w5131;
	wire w5132;
	wire w5133;
	wire w5134;
	wire w5135;
	wire w5136;
	wire w5137;
	wire w5138;
	wire w5139;
	wire w5140;
	wire w5141;
	wire w5142;
	wire w5143;
	wire w5144;
	wire w5145;
	wire w5146;
	wire w5147;
	wire w5148;
	wire w5149;
	wire w5150;
	wire w5151;
	wire w5152;
	wire w5153;
	wire w5154;
	wire w5155;
	wire w5156;
	wire w5157;
	wire w5158;
	wire w5159;
	wire w5160;
	wire w5161;
	wire w5162;
	wire w5163;
	wire w5164;
	wire w5165;
	wire w5166;
	wire w5167;
	wire w5168;
	wire w5169;
	wire w5170;
	wire w5171;
	wire w5172;
	wire w5173;
	wire w5174;
	wire w5175;
	wire w5176;
	wire w5177;
	wire w5178;
	wire w5179;
	wire w5180;
	wire w5181;
	wire w5182;
	wire w5183;
	wire w5184;
	wire w5185;
	wire w5186;
	wire w5187;
	wire w5188;
	wire w5189;
	wire w5190;
	wire w5191;
	wire w5192;
	wire w5193;
	wire w5194;
	wire w5195;
	wire w5196;
	wire w5197;
	wire w5198;
	wire w5199;
	wire w5200;
	wire w5201;
	wire w5202;
	wire w5203;
	wire w5204;
	wire w5205;
	wire w5206;
	wire w5207;
	wire w5208;
	wire w5209;
	wire w5210;
	wire w5211;
	wire w5212;
	wire w5213;
	wire w5214;
	wire w5215;
	wire w5216;
	wire w5217;
	wire w5218;
	wire w5219;
	wire w5220;
	wire w5221;
	wire w5222;
	wire w5223;
	wire w5224;
	wire w5225;
	wire w5226;
	wire w5227;
	wire w5228;
	wire w5229;
	wire w5230;
	wire w5231;
	wire w5232;
	wire w5233;
	wire w5234;
	wire w5235;
	wire w5236;
	wire w5237;
	wire w5238;
	wire w5239;
	wire w5240;
	wire w5241;
	wire w5242;
	wire w5243;
	wire w5244;
	wire w5245;
	wire w5246;
	wire w5247;
	wire w5248;
	wire w5249;
	wire w5250;
	wire w5251;
	wire w5252;
	wire w5253;
	wire w5254;
	wire w5255;
	wire w5256;
	wire w5257;
	wire w5258;
	wire w5259;
	wire w5260;
	wire w5261;
	wire w5262;
	wire w5263;
	wire w5264;
	wire w5265;
	wire w5266;
	wire w5267;
	wire w5268;
	wire w5269;
	wire w5270;
	wire w5271;
	wire w5272;
	wire w5273;
	wire w5274;
	wire w5275;
	wire w5276;
	wire w5277;
	wire w5278;
	wire w5279;
	wire w5280;
	wire w5281;
	wire w5282;
	wire w5283;
	wire w5284;
	wire w5285;
	wire w5286;
	wire w5287;
	wire w5288;
	wire w5289;
	wire w5290;
	wire w5291;
	wire w5292;
	wire w5293;
	wire w5294;
	wire w5295;
	wire w5296;
	wire w5297;
	wire w5298;
	wire w5299;
	wire w5300;
	wire w5301;
	wire w5302;
	wire w5303;
	wire w5304;
	wire w5305;
	wire w5306;
	wire w5307;
	wire w5308;
	wire w5309;
	wire w5310;
	wire w5311;
	wire w5312;
	wire w5313;
	wire w5314;
	wire w5315;
	wire w5316;
	wire w5317;
	wire w5318;
	wire w5319;
	wire w5320;
	wire w5321;
	wire w5322;
	wire w5323;
	wire w5324;
	wire w5325;
	wire w5326;
	wire w5327;
	wire w5328;
	wire w5329;
	wire w5330;
	wire w5331;
	wire w5332;
	wire w5333;
	wire w5334;
	wire w5335;
	wire w5336;
	wire w5337;
	wire w5338;
	wire w5339;
	wire w5340;
	wire w5341;
	wire w5342;
	wire w5343;
	wire w5344;
	wire w5345;
	wire w5346;
	wire w5347;
	wire w5348;
	wire w5349;
	wire w5350;
	wire w5351;
	wire w5352;
	wire w5353;
	wire w5354;
	wire w5355;
	wire w5356;
	wire w5357;
	wire w5358;
	wire w5359;
	wire w5360;
	wire w5361;
	wire w5362;
	wire w5363;
	wire w5364;
	wire w5365;
	wire w5366;
	wire w5367;
	wire w5368;
	wire w5369;
	wire w5370;
	wire w5371;
	wire w5372;
	wire w5373;
	wire w5374;
	wire w5375;
	wire w5376;
	wire w5377;
	wire w5378;
	wire w5379;
	wire w5380;
	wire w5381;
	wire w5382;
	wire w5383;
	wire w5384;
	wire w5385;
	wire w5386;
	wire w5387;
	wire w5388;
	wire w5389;
	wire w5390;
	wire w5391;
	wire w5392;
	wire w5393;
	wire w5394;
	wire w5395;
	wire w5396;
	wire w5397;
	wire w5398;
	wire w5399;
	wire w5400;
	wire w5401;
	wire w5402;
	wire w5403;
	wire w5404;
	wire w5405;
	wire w5406;
	wire w5407;
	wire w5408;
	wire w5409;
	wire w5410;
	wire w5411;
	wire w5412;
	wire w5413;
	wire w5414;
	wire w5415;
	wire w5416;
	wire w5417;
	wire w5418;
	wire w5419;
	wire w5420;
	wire w5421;
	wire w5422;
	wire w5423;
	wire w5424;
	wire w5425;
	wire w5426;
	wire w5427;
	wire w5428;
	wire w5429;
	wire w5430;
	wire w5431;
	wire w5432;
	wire w5433;
	wire w5434;
	wire w5435;
	wire w5436;
	wire w5437;
	wire w5438;
	wire w5439;
	wire w5440;
	wire w5441;
	wire w5442;
	wire w5443;
	wire w5444;
	wire w5445;
	wire w5446;
	wire w5447;
	wire w5448;
	wire w5449;
	wire w5450;
	wire w5451;
	wire w5452;
	wire w5453;
	wire w5454;
	wire w5455;
	wire w5456;
	wire w5457;
	wire w5458;
	wire w5459;
	wire w5460;
	wire w5461;
	wire w5462;
	wire w5463;
	wire w5464;
	wire w5465;
	wire w5466;
	wire w5467;
	wire w5468;
	wire w5469;
	wire w5470;
	wire w5471;
	wire w5472;
	wire w5473;
	wire w5474;
	wire w5475;
	wire w5476;
	wire w5477;
	wire w5478;
	wire w5479;
	wire w5480;
	wire w5481;
	wire w5482;
	wire w5483;
	wire w5484;
	wire w5485;
	wire w5486;
	wire w5487;
	wire w5488;
	wire w5489;
	wire w5490;
	wire w5491;
	wire w5492;
	wire w5493;
	wire w5494;
	wire w5495;
	wire w5496;
	wire w5497;
	wire w5498;
	wire w5499;
	wire w5500;
	wire w5501;
	wire w5502;
	wire w5503;
	wire w5504;
	wire w5505;
	wire w5506;
	wire w5507;
	wire w5508;
	wire w5509;
	wire w5510;
	wire w5511;
	wire w5512;
	wire w5513;
	wire w5514;
	wire w5515;
	wire w5516;
	wire w5517;
	wire w5518;
	wire w5519;
	wire w5520;
	wire w5521;
	wire w5522;
	wire w5523;
	wire w5524;
	wire w5525;
	wire w5526;
	wire w5527;
	wire w5528;
	wire w5529;
	wire w5530;
	wire w5531;
	wire w5532;
	wire w5533;
	wire w5534;
	wire w5535;
	wire w5536;
	wire w5537;
	wire w5538;
	wire w5539;
	wire w5540;
	wire w5541;
	wire w5542;
	wire w5543;
	wire w5544;
	wire w5545;
	wire w5546;
	wire w5547;
	wire w5548;
	wire w5549;
	wire w5550;
	wire w5551;
	wire w5552;
	wire w5553;
	wire w5554;
	wire w5555;
	wire w5556;
	wire w5557;
	wire w5558;
	wire w5559;
	wire w5560;
	wire w5561;
	wire w5562;
	wire w5563;
	wire w5564;
	wire w5565;
	wire w5566;
	wire w5567;
	wire w5568;
	wire w5569;
	wire w5570;
	wire w5571;
	wire w5572;
	wire w5573;
	wire w5574;
	wire w5575;
	wire w5576;
	wire w5577;
	wire w5578;
	wire w5579;
	wire w5580;
	wire w5581;
	wire w5582;
	wire w5583;
	wire w5584;
	wire w5585;
	wire w5586;
	wire w5587;
	wire w5588;
	wire w5589;
	wire w5590;
	wire w5591;
	wire w5592;
	wire w5593;
	wire w5594;
	wire w5595;
	wire w5596;
	wire w5597;
	wire w5598;
	wire w5599;
	wire w5600;
	wire w5601;
	wire w5602;
	wire w5603;
	wire w5604;
	wire w5605;
	wire w5606;
	wire w5607;
	wire w5608;
	wire w5609;
	wire w5610;
	wire w5611;
	wire w5612;
	wire w5613;
	wire w5614;
	wire w5615;
	wire w5616;
	wire w5617;
	wire w5618;
	wire w5619;
	wire w5620;
	wire w5621;
	wire w5622;
	wire w5623;
	wire w5624;
	wire w5625;
	wire w5626;
	wire w5627;
	wire w5628;
	wire w5629;
	wire w5630;
	wire w5631;
	wire w5632;
	wire w5633;
	wire w5634;
	wire w5635;
	wire w5636;
	wire w5637;
	wire w5638;
	wire w5639;
	wire w5640;
	wire w5641;
	wire w5642;
	wire w5643;
	wire w5644;
	wire w5645;
	wire w5646;
	wire w5647;
	wire w5648;
	wire w5649;
	wire w5650;
	wire w5651;
	wire w5652;
	wire w5653;
	wire w5654;
	wire w5655;
	wire w5656;
	wire w5657;
	wire w5658;
	wire w5659;
	wire w5660;
	wire w5661;
	wire w5662;
	wire w5663;
	wire w5664;
	wire w5665;
	wire w5666;
	wire w5667;
	wire w5668;
	wire w5669;
	wire w5670;
	wire w5671;
	wire w5672;
	wire w5673;
	wire w5674;
	wire w5675;
	wire w5676;
	wire w5677;
	wire w5678;
	wire w5679;
	wire w5680;
	wire w5681;
	wire w5682;
	wire w5683;
	wire w5684;
	wire w5685;
	wire w5686;
	wire w5687;
	wire w5688;
	wire w5689;
	wire w5690;
	wire w5691;
	wire w5692;
	wire w5693;
	wire w5694;
	wire w5695;
	wire w5696;
	wire w5697;
	wire w5698;
	wire w5699;
	wire w5700;
	wire w5701;
	wire w5702;
	wire w5703;
	wire w5704;
	wire w5705;
	wire w5706;
	wire w5707;
	wire w5708;
	wire w5709;
	wire w5710;
	wire w5711;
	wire w5712;
	wire w5713;
	wire w5714;
	wire w5715;
	wire w5716;
	wire w5717;
	wire w5718;
	wire w5719;
	wire w5720;
	wire w5721;
	wire w5722;
	wire w5723;
	wire w5724;
	wire w5725;
	wire w5726;
	wire w5727;
	wire w5728;
	wire w5729;
	wire w5730;
	wire w5731;
	wire w5732;
	wire w5733;
	wire w5734;
	wire w5735;
	wire w5736;
	wire w5737;
	wire w5738;
	wire w5739;
	wire w5740;
	wire w5741;
	wire w5742;
	wire w5743;
	wire w5744;
	wire w5745;
	wire w5746;
	wire w5747;
	wire w5748;
	wire w5749;
	wire w5750;
	wire w5751;
	wire w5752;
	wire w5753;
	wire w5754;
	wire w5755;
	wire w5756;
	wire w5757;
	wire w5758;
	wire w5759;
	wire w5760;
	wire w5761;
	wire w5762;
	wire w5763;
	wire w5764;
	wire w5765;
	wire w5766;
	wire w5767;
	wire w5768;
	wire w5769;
	wire w5770;
	wire w5771;
	wire w5772;
	wire w5773;
	wire w5774;
	wire w5775;
	wire w5776;
	wire w5777;
	wire w5778;
	wire w5779;
	wire w5780;
	wire w5781;
	wire w5782;
	wire w5783;
	wire w5784;
	wire w5785;
	wire w5786;
	wire w5787;
	wire w5788;
	wire w5789;
	wire w5790;
	wire w5791;
	wire w5792;
	wire w5793;
	wire w5794;
	wire w5795;
	wire w5796;
	wire w5797;
	wire w5798;
	wire w5799;
	wire w5800;
	wire w5801;
	wire w5802;
	wire w5803;
	wire w5804;
	wire w5805;
	wire w5806;
	wire w5807;
	wire w5808;
	wire w5809;
	wire w5810;
	wire w5811;
	wire w5812;
	wire w5813;
	wire w5814;
	wire w5815;
	wire w5816;
	wire w5817;
	wire w5818;
	wire w5819;
	wire w5820;
	wire w5821;
	wire w5822;
	wire w5823;
	wire w5824;
	wire w5825;
	wire w5826;
	wire w5827;
	wire w5828;
	wire w5829;
	wire w5830;
	wire w5831;
	wire w5832;
	wire w5833;
	wire w5834;
	wire w5835;
	wire w5836;
	wire w5837;
	wire w5838;
	wire w5839;
	wire w5840;
	wire w5841;
	wire w5842;
	wire w5843;
	wire w5844;
	wire w5845;
	wire w5846;
	wire w5847;
	wire w5848;
	wire w5849;
	wire w5850;
	wire w5851;
	wire w5852;
	wire w5853;
	wire w5854;
	wire w5855;
	wire w5856;
	wire w5857;
	wire w5858;
	wire w5859;
	wire w5860;
	wire w5861;
	wire w5862;
	wire w5863;
	wire w5864;
	wire w5865;
	wire w5866;
	wire w5867;
	wire w5868;
	wire w5869;
	wire w5870;
	wire w5871;
	wire w5872;
	wire w5873;
	wire w5874;
	wire w5875;
	wire w5876;
	wire w5877;
	wire w5878;
	wire w5879;
	wire w5880;
	wire w5881;
	wire w5882;
	wire w5883;
	wire w5884;
	wire w5885;
	wire w5886;
	wire w5887;
	wire w5888;
	wire w5889;
	wire w5890;
	wire w5891;
	wire w5892;
	wire w5893;
	wire w5894;
	wire w5895;
	wire w5896;
	wire w5897;
	wire w5898;
	wire w5899;
	wire w5900;
	wire w5901;
	wire w5902;
	wire w5903;
	wire w5904;
	wire w5905;
	wire w5906;
	wire w5907;
	wire w5908;
	wire w5909;
	wire w5910;
	wire w5911;
	wire w5912;
	wire w5913;
	wire w5914;
	wire w5915;
	wire w5916;
	wire w5917;
	wire w5918;
	wire w5919;
	wire w5920;
	wire w5921;
	wire w5922;
	wire w5923;
	wire w5924;
	wire w5925;
	wire w5926;
	wire w5927;
	wire w5928;
	wire w5929;
	wire w5930;
	wire w5931;
	wire w5932;
	wire w5933;
	wire w5934;
	wire w5935;
	wire w5936;
	wire w5937;
	wire w5938;
	wire w5939;
	wire w5940;
	wire w5941;
	wire w5942;
	wire w5943;
	wire w5944;
	wire w5945;
	wire w5946;
	wire w5947;
	wire w5948;
	wire w5949;
	wire w5950;
	wire w5951;
	wire w5952;
	wire w5953;
	wire w5954;
	wire w5955;
	wire w5956;
	wire w5957;
	wire w5958;
	wire w5959;
	wire w5960;
	wire w5961;
	wire w5962;
	wire w5963;
	wire w5964;
	wire w5965;
	wire w5966;
	wire w5967;
	wire w5968;
	wire w5969;
	wire w5970;
	wire w5971;
	wire w5972;
	wire w5973;
	wire w5974;
	wire w5975;
	wire w5976;
	wire w5977;
	wire w5978;
	wire w5979;
	wire w5980;
	wire w5981;
	wire w5982;
	wire w5983;
	wire w5984;
	wire w5985;
	wire w5986;
	wire w5987;
	wire w5988;
	wire w5989;
	wire w5990;
	wire w5991;
	wire w5992;
	wire w5993;
	wire w5994;
	wire w5995;
	wire w5996;
	wire w5997;
	wire w5998;
	wire w5999;
	wire w6000;
	wire w6001;
	wire w6002;
	wire w6003;
	wire w6004;
	wire w6005;
	wire w6006;
	wire w6007;
	wire w6008;
	wire w6009;
	wire w6010;
	wire w6011;
	wire w6012;
	wire w6013;
	wire w6014;
	wire w6015;
	wire w6016;
	wire w6017;
	wire w6018;
	wire w6019;
	wire w6020;
	wire w6021;
	wire w6022;
	wire w6023;
	wire w6024;
	wire w6025;
	wire w6026;
	wire w6027;
	wire w6028;
	wire w6029;
	wire w6030;
	wire w6031;
	wire w6032;
	wire w6033;
	wire w6034;
	wire w6035;
	wire w6036;
	wire w6037;
	wire w6038;
	wire w6039;
	wire w6040;
	wire w6041;
	wire w6042;
	wire w6043;
	wire w6044;
	wire w6045;
	wire w6046;
	wire w6047;
	wire w6048;
	wire w6049;
	wire w6050;
	wire w6051;
	wire w6052;
	wire w6053;
	wire w6054;
	wire w6055;
	wire w6056;
	wire w6057;
	wire w6058;
	wire w6059;
	wire w6060;
	wire w6061;
	wire w6062;
	wire w6063;
	wire w6064;
	wire w6065;
	wire w6066;
	wire w6067;
	wire w6068;
	wire w6069;
	wire w6070;
	wire w6071;
	wire w6072;
	wire w6073;
	wire w6074;
	wire w6075;
	wire w6076;
	wire w6077;
	wire w6078;
	wire w6079;
	wire w6080;
	wire w6081;
	wire w6082;
	wire w6083;
	wire w6084;
	wire w6085;
	wire w6086;
	wire w6087;
	wire w6088;
	wire w6089;
	wire w6090;
	wire w6091;
	wire w6092;
	wire w6093;
	wire w6094;
	wire w6095;
	wire w6096;
	wire w6097;
	wire w6098;
	wire w6099;
	wire w6100;
	wire w6101;
	wire w6102;
	wire w6103;
	wire w6104;
	wire w6105;
	wire w6106;
	wire w6107;
	wire w6108;
	wire w6109;
	wire w6110;
	wire w6111;
	wire w6112;
	wire w6113;
	wire w6114;
	wire w6115;
	wire w6116;
	wire w6117;
	wire w6118;
	wire w6119;
	wire w6120;
	wire w6121;
	wire w6122;
	wire w6123;
	wire w6124;
	wire w6125;
	wire w6126;
	wire w6127;
	wire w6128;
	wire w6129;
	wire w6130;
	wire w6131;
	wire w6132;
	wire w6133;
	wire w6134;
	wire w6135;
	wire w6136;
	wire w6137;
	wire w6138;
	wire w6139;
	wire w6140;
	wire w6141;
	wire w6142;
	wire w6143;
	wire w6144;
	wire w6145;
	wire w6146;
	wire w6147;
	wire w6148;
	wire w6149;
	wire w6150;
	wire w6151;
	wire w6152;
	wire w6153;
	wire w6154;
	wire w6155;
	wire w6156;
	wire w6157;
	wire w6158;
	wire w6159;
	wire w6160;
	wire w6161;
	wire w6162;
	wire w6163;
	wire w6164;
	wire w6165;
	wire w6166;
	wire w6167;
	wire w6168;
	wire w6169;
	wire w6170;
	wire w6171;
	wire w6172;
	wire w6173;
	wire w6174;
	wire w6175;
	wire w6176;
	wire w6177;
	wire w6178;
	wire w6179;
	wire w6180;
	wire w6181;
	wire w6182;
	wire w6183;
	wire w6184;
	wire w6185;
	wire w6186;
	wire w6187;
	wire w6188;
	wire w6189;
	wire w6190;
	wire w6191;
	wire w6192;
	wire w6193;
	wire w6194;
	wire w6195;
	wire w6196;
	wire w6197;
	wire w6198;
	wire w6199;
	wire w6200;
	wire w6201;
	wire w6202;
	wire w6203;
	wire w6204;
	wire w6205;
	wire w6206;
	wire w6207;
	wire w6208;
	wire w6209;
	wire w6210;
	wire w6211;
	wire w6212;
	wire w6213;
	wire w6214;
	wire w6215;
	wire w6216;
	wire w6217;
	wire w6218;
	wire w6219;
	wire w6220;
	wire w6221;
	wire w6222;
	wire w6223;
	wire w6224;
	wire w6225;
	wire w6226;
	wire w6227;
	wire w6228;
	wire w6229;
	wire w6230;
	wire w6231;
	wire w6232;
	wire w6233;
	wire w6234;
	wire w6235;
	wire w6236;
	wire w6237;
	wire w6238;
	wire w6239;
	wire w6240;
	wire w6241;
	wire w6242;
	wire w6243;
	wire w6244;
	wire w6245;
	wire w6246;
	wire w6247;
	wire w6248;
	wire w6249;
	wire w6250;
	wire w6251;
	wire w6252;
	wire w6253;
	wire w6254;
	wire w6255;
	wire w6256;
	wire w6257;
	wire w6258;
	wire w6259;
	wire w6260;
	wire w6261;
	wire w6262;
	wire w6263;
	wire w6264;
	wire w6265;
	wire w6266;
	wire w6267;
	wire w6268;
	wire w6269;
	wire w6270;
	wire w6271;
	wire w6272;
	wire w6273;
	wire w6274;
	wire w6275;
	wire w6276;
	wire w6277;
	wire w6278;
	wire w6279;
	wire w6280;
	wire w6281;
	wire w6282;
	wire w6283;
	wire w6284;
	wire w6285;
	wire w6286;
	wire w6287;
	wire w6288;
	wire w6289;
	wire w6290;
	wire w6291;
	wire w6292;
	wire w6293;
	wire w6294;
	wire w6295;
	wire w6296;
	wire w6297;
	wire w6298;
	wire w6299;
	wire w6300;
	wire w6301;
	wire w6302;
	wire w6303;
	wire w6304;
	wire w6305;
	wire w6306;
	wire w6307;
	wire w6308;
	wire w6309;
	wire w6310;
	wire w6311;
	wire w6312;
	wire w6313;
	wire w6314;
	wire w6315;
	wire w6316;
	wire w6317;
	wire w6318;
	wire w6319;
	wire w6320;
	wire w6321;
	wire w6322;
	wire w6323;
	wire w6324;
	wire w6325;
	wire w6326;
	wire w6327;
	wire w6328;
	wire w6329;
	wire w6330;
	wire w6331;
	wire w6332;
	wire w6333;
	wire w6334;
	wire w6335;
	wire w6336;
	wire w6337;
	wire w6338;
	wire w6339;
	wire w6340;
	wire w6341;
	wire w6342;
	wire w6343;
	wire w6344;
	wire w6345;
	wire w6346;
	wire w6347;
	wire w6348;
	wire w6349;
	wire w6350;
	wire w6351;
	wire w6352;
	wire w6353;
	wire w6354;
	wire w6355;
	wire w6356;
	wire w6357;
	wire w6358;
	wire w6359;
	wire w6360;
	wire w6361;
	wire w6362;
	wire w6363;
	wire w6364;
	wire w6365;
	wire w6366;
	wire w6367;
	wire w6368;
	wire w6369;
	wire w6370;
	wire w6371;
	wire w6372;
	wire w6373;
	wire w6374;
	wire w6375;
	wire w6376;
	wire w6377;
	wire w6378;
	wire w6379;
	wire w6380;
	wire w6381;
	wire w6382;
	wire w6383;
	wire w6384;
	wire w6385;
	wire w6386;
	wire w6387;
	wire w6388;
	wire w6389;
	wire w6390;
	wire w6391;
	wire w6392;
	wire w6393;
	wire w6394;
	wire w6395;
	wire w6396;
	wire w6397;
	wire w6398;
	wire w6399;
	wire w6400;
	wire w6401;
	wire w6402;
	wire w6403;
	wire w6404;
	wire w6405;
	wire w6406;
	wire w6407;
	wire w6408;
	wire w6409;
	wire w6410;
	wire w6411;
	wire w6412;
	wire w6413;
	wire w6414;
	wire w6415;
	wire w6416;
	wire w6417;
	wire w6418;
	wire w6419;
	wire w6420;
	wire w6421;
	wire w6422;
	wire w6423;
	wire w6424;
	wire w6425;
	wire w6426;
	wire w6427;
	wire w6428;
	wire w6429;
	wire w6430;
	wire w6431;
	wire w6432;
	wire w6433;
	wire w6434;
	wire w6435;
	wire w6436;
	wire w6437;
	wire w6438;
	wire w6439;
	wire w6440;
	wire w6441;
	wire w6442;
	wire w6443;
	wire w6444;
	wire w6445;
	wire w6446;
	wire w6447;
	wire w6448;
	wire w6449;
	wire w6450;
	wire w6451;
	wire w6452;
	wire w6453;
	wire w6454;
	wire w6455;
	wire w6456;
	wire w6457;
	wire w6458;
	wire w6459;
	wire w6460;
	wire w6461;
	wire w6462;
	wire w6463;
	wire w6464;
	wire w6465;
	wire w6466;
	wire w6467;
	wire w6468;
	wire w6469;
	wire w6470;
	wire w6471;
	wire w6472;
	wire w6473;
	wire w6474;
	wire w6475;
	wire w6476;
	wire w6477;
	wire w6478;
	wire w6479;
	wire w6480;
	wire w6481;
	wire w6482;
	wire w6483;
	wire w6484;
	wire w6485;
	wire w6486;
	wire w6487;
	wire w6488;
	wire w6489;
	wire w6490;
	wire w6491;
	wire w6492;
	wire w6493;
	wire w6494;
	wire w6495;
	wire w6496;
	wire w6497;
	wire w6498;
	wire w6499;
	wire w6500;
	wire w6501;
	wire w6502;
	wire w6503;
	wire w6504;
	wire w6505;
	wire w6506;
	wire w6507;
	wire w6508;
	wire w6509;
	wire w6510;
	wire w6511;
	wire w6512;
	wire w6513;
	wire w6514;
	wire w6515;
	wire w6516;
	wire w6517;
	wire w6518;
	wire w6519;
	wire w6520;
	wire w6521;
	wire w6522;
	wire w6523;
	wire w6524;
	wire w6525;
	wire w6526;
	wire w6527;
	wire w6528;
	wire w6529;
	wire w6530;
	wire w6531;
	wire w6532;
	wire w6533;
	wire w6534;
	wire w6535;
	wire w6536;
	wire w6537;
	wire w6538;
	wire w6539;
	wire w6540;
	wire w6541;
	wire w6542;
	wire w6543;
	wire w6544;
	wire w6545;
	wire w6546;
	wire w6547;
	wire w6548;
	wire w6549;
	wire w6550;
	wire w6551;
	wire w6552;
	wire w6553;
	wire w6554;
	wire w6555;
	wire w6556;
	wire w6557;
	wire w6558;
	wire w6559;
	wire w6560;
	wire w6561;
	wire w6562;
	wire w6563;
	wire w6564;
	wire w6565;
	wire w6566;
	wire w6567;
	wire w6568;
	wire w6569;
	wire w6570;
	wire w6571;
	wire w6572;
	wire w6573;
	wire w6574;
	wire w6575;
	wire w6576;
	wire w6577;
	wire w6578;
	wire w6579;
	wire w6580;
	wire w6581;
	wire w6582;
	wire w6583;
	wire w6584;
	wire w6585;
	wire w6586;
	wire w6587;
	wire w6588;
	wire w6589;
	wire w6590;
	wire w6591;
	wire w6592;
	wire w6593;
	wire w6594;
	wire w6595;
	wire w6596;
	wire w6597;
	wire w6598;
	wire w6599;
	wire w6600;
	wire w6601;
	wire w6602;
	wire w6603;
	wire w6604;
	wire w6605;
	wire w6606;
	wire w6607;
	wire w6608;
	wire w6609;
	wire w6610;
	wire w6611;
	wire w6612;
	wire w6613;
	wire w6614;
	wire w6615;
	wire w6616;
	wire w6617;
	wire w6618;
	wire w6619;
	wire w6620;
	wire w6621;
	wire w6622;
	wire w6623;
	wire w6624;
	wire w6625;
	wire w6626;
	wire w6627;
	wire w6628;
	wire w6629;
	wire w6630;
	wire w6631;
	wire w6632;
	wire w6633;
	wire w6634;
	wire w6635;
	wire w6636;
	wire w6637;
	wire w6638;
	wire w6639;
	wire w6640;
	wire w6641;
	wire w6642;
	wire w6643;
	wire w6644;
	wire w6645;
	wire w6646;
	wire w6647;
	wire w6648;
	wire w6649;
	wire w6650;
	wire w6651;
	wire w6652;
	wire w6653;
	wire w6654;
	wire w6655;
	wire w6656;
	wire w6657;
	wire w6658;
	wire w6659;
	wire w6660;
	wire w6661;
	wire w6662;
	wire w6663;
	wire w6664;
	wire w6665;
	wire w6666;
	wire w6667;
	wire w6668;
	wire w6669;
	wire w6670;
	wire w6671;
	wire w6672;
	wire w6673;
	wire w6674;
	wire w6675;
	wire w6676;
	wire w6677;
	wire w6678;
	wire w6679;
	wire w6680;
	wire w6681;
	wire w6682;
	wire w6683;
	wire w6684;
	wire w6685;
	wire w6686;
	wire w6687;
	wire w6688;
	wire w6689;
	wire w6690;
	wire w6691;
	wire w6692;
	wire w6693;
	wire w6694;
	wire w6695;
	wire w6696;
	wire w6697;
	wire w6698;
	wire w6699;
	wire w6700;
	wire w6701;
	wire w6702;
	wire w6703;
	wire w6704;
	wire w6705;
	wire w6706;
	wire w6707;
	wire w6708;
	wire w6709;
	wire w6710;
	wire w6711;
	wire w6712;
	wire w6713;
	wire w6714;
	wire w6715;
	wire w6716;
	wire w6717;
	wire w6718;
	wire w6719;
	wire w6720;
	wire w6721;
	wire w6722;
	wire w6723;
	wire w6724;
	wire w6725;
	wire w6726;
	wire w6727;
	wire w6728;
	wire w6729;
	wire w6730;
	wire w6731;
	wire w6732;
	wire w6733;
	wire w6734;
	wire w6735;
	wire w6736;
	wire w6737;
	wire w6738;
	wire w6739;
	wire w6740;
	wire w6741;
	wire w6742;
	wire w6743;
	wire w6744;
	wire w6745;
	wire w6746;
	wire w6747;
	wire w6748;
	wire w6749;
	wire w6750;
	wire w6751;
	wire w6752;
	wire w6753;
	wire w6754;
	wire w6755;
	wire w6756;
	wire w6757;
	wire w6758;
	wire w6759;
	wire w6760;
	wire w6761;
	wire w6762;
	wire w6763;
	wire w6764;
	wire w6765;
	wire w6766;
	wire w6767;
	wire w6768;
	wire w6769;
	wire w6770;
	wire w6771;
	wire w6772;
	wire w6773;
	wire w6774;
	wire w6775;
	wire w6776;
	wire w6777;
	wire w6778;
	wire w6779;
	wire w6780;
	wire w6781;
	wire w6782;
	wire w6783;
	wire w6784;
	wire w6785;
	wire w6786;
	wire w6787;
	wire w6788;
	wire w6789;
	wire w6790;
	wire w6791;
	wire w6792;
	wire w6793;
	wire w6794;
	wire w6795;
	wire w6796;
	wire w6797;
	wire w6798;
	wire w6799;
	wire w6800;
	wire w6801;
	wire w6802;
	wire w6803;
	wire w6804;
	wire w6805;
	wire w6806;
	wire w6807;
	wire w6808;
	wire w6809;
	wire w6810;
	wire w6811;
	wire w6812;
	wire w6813;
	wire w6814;
	wire w6815;
	wire w6816;
	wire w6817;
	wire w6818;
	wire w6819;
	wire w6820;
	wire w6821;
	wire w6822;
	wire w6823;
	wire w6824;
	wire w6825;
	wire w6826;
	wire w6827;
	wire w6828;
	wire w6829;
	wire w6830;
	wire w6831;
	wire w6832;
	wire w6833;
	wire w6834;
	wire w6835;
	wire w6836;
	wire w6837;
	wire w6838;
	wire w6839;
	wire w6840;
	wire w6841;
	wire w6842;

	assign CH0_EN = w2028;
	assign CH0VOL[0] = w2031;
	assign CH0VOL[1] = w2032;
	assign CH1_EN = w2027;
	assign CH1VOL[0] = w2091;
	assign CH1VOL[1] = w2092;
	assign CH2_EN = w2029;
	assign CH2VOL[0] = w2111;
	assign CH2VOL[1] = w2110;
	assign CH3_EN = w2026;
	assign CH3VOL[0] = w2133;
	assign CH3VOL[1] = w2132;
	assign PSGDAC0[0] = w2033;
	assign PSGDAC0[1] = w2034;
	assign PSGDAC0[2] = w2035;
	assign PSGDAC0[3] = w2036;
	assign PSGDAC0[4] = w2037;
	assign PSGDAC0[5] = w2038;
	assign PSGDAC0[6] = w2039;
	assign PSGDAC0[7] = w2040;
	assign PSGDAC1[0] = w2093;
	assign PSGDAC1[1] = w2094;
	assign PSGDAC1[2] = w2095;
	assign PSGDAC1[3] = w2096;
	assign PSGDAC1[4] = w2097;
	assign PSGDAC1[5] = w2098;
	assign PSGDAC1[6] = w2099;
	assign PSGDAC1[7] = w2100;
	assign PSGDAC2[0] = w2122;
	assign PSGDAC2[1] = w2123;
	assign PSGDAC2[2] = w2124;
	assign PSGDAC2[3] = w2125;
	assign PSGDAC2[4] = w2126;
	assign PSGDAC2[5] = w2127;
	assign PSGDAC2[6] = w2128;
	assign PSGDAC2[7] = w2129;
	assign PSGDAC3[0] = w2131;
	assign PSGDAC3[1] = w2130;
	assign PSGDAC3[2] = w2138;
	assign PSGDAC3[3] = w2137;
	assign PSGDAC3[4] = w2136;
	assign PSGDAC3[5] = w2135;
	assign PSGDAC3[6] = w2134;
	assign PSGDAC3[7] = w2139;
	assign w1210 = CAi[22];
	assign CAo[22] = w1370;
	assign CA[19] = CA[19];
	assign DTACK_OUT = w1059;
	assign Z80_INT = w1060;
	assign RA[7] = w1118;
	assign RA[6] = w1117;
	assign RA[5] = w1116;
	assign RA[4] = w1115;
	assign RA[2] = w1113;
	assign RA[1] = w1112;
	assign RA[0] = w1111;
	assign nRAS0 = w1346;
	assign RA[3] = w1114;
	assign nCAS0 = w1419;
	assign nOE0 = w1410;
	assign nLWR = w1411;
	assign nUWR = w1321;
	assign w1398 = DTACK_IN;
	assign w1006 = RnW;
	assign w1390 = nLDS;
	assign w1381 = nUDS;
	assign w1263 = nAS;
	assign w1379 = nM1;
	assign w1380 = nWR;
	assign w1377 = nRD;
	assign w1378 = nIORQ;
	assign nILP2 = w1383;
	assign nILP1 = w1382;
	assign w1244 = nINTAK;
	assign w1376 = nMREQ;
	assign w1246 = nBG;
	assign BGACK_OUT = w1261;
	assign w1397 = BGACK_IN;
	assign nBR = w1440;
	assign VSYNC = w1708;
	assign nCSYNC = w2015;
	assign w1702 = nCSYNC_IN;
	assign nHSYNC = w1768;
	assign w1986 = nHSYNC_IN;
	assign DB[15] = w358;
	assign DB[14] = DB[14];
	assign DB[13] = DB[13];
	assign DB[12] = DB[12];
	assign DB[11] = w325;
	assign DB[10] = DB[10];
	assign DB[9] = DB[9];
	assign DB[8] = DB[8];
	assign DB[7] = w160;
	assign DB[6] = DB[6];
	assign DB[5] = DB[5];
	assign DB[4] = DB[4];
	assign DB[3] = w156;
	assign DB[2] = DB[2];
	assign DB[1] = DB[1];
	assign DB[0] = DB[0];
	assign CA[0] = CA[0];
	assign CA[1] = CA[1];
	assign CA[2] = CA[2];
	assign CA[3] = CA[3];
	assign CA[4] = CA[4];
	assign CA[5] = CA[5];
	assign CA[6] = CA[6];
	assign CA[7] = CA[7];
	assign CA[8] = CA[8];
	assign CA[9] = CA[9];
	assign CA[10] = CA[10];
	assign CA[11] = CA[11];
	assign CA[12] = CA[12];
	assign CA[13] = CA[13];
	assign CA[14] = CA[14];
	assign CA[15] = CA[15];
	assign CA[17] = CA[17];
	assign CA[18] = CA[18];
	assign CA[20] = CA[20];
	assign CA[21] = CA[21];
	assign R_DAC[0] = w2973;
	assign R_DAC[1] = w2938;
	assign R_DAC[2] = w2972;
	assign R_DAC[3] = w2937;
	assign R_DAC[4] = w2971;
	assign R_DAC[5] = w2970;
	assign R_DAC[6] = w2969;
	assign R_DAC[7] = w2968;
	assign R_DAC[8] = w2934;
	assign G_DAC[0] = w2966;
	assign G_DAC[1] = w2965;
	assign G_DAC[2] = w2928;
	assign G_DAC[3] = w2927;
	assign G_DAC[4] = w2926;
	assign G_DAC[5] = w2925;
	assign G_DAC[6] = w2924;
	assign G_DAC[7] = w2923;
	assign G_DAC[8] = w2922;
	assign R_DAC[9] = w2935;
	assign R_DAC[10] = w2932;
	assign R_DAC[11] = w2936;
	assign R_DAC[12] = w2931;
	assign R_DAC[13] = w2933;
	assign R_DAC[14] = w2930;
	assign R_DAC[15] = w2929;
	assign R_DAC[16] = w2967;
	assign B_DAC[0] = w2914;
	assign B_DAC[1] = w2964;
	assign B_DAC[2] = w2960;
	assign B_DAC[3] = w2961;
	assign B_DAC[4] = w2962;
	assign B_DAC[5] = w2959;
	assign B_DAC[6] = w2963;
	assign B_DAC[7] = w3021;
	assign B_DAC[8] = w2915;
	assign G_DAC[9] = w2916;
	assign G_DAC[10] = w2921;
	assign G_DAC[11] = w2920;
	assign G_DAC[12] = w3019;
	assign G_DAC[13] = w2919;
	assign G_DAC[14] = w2918;
	assign G_DAC[15] = w2917;
	assign G_DAC[16] = w3020;
	assign B_DAC[9] = w2912;
	assign B_DAC[10] = w2913;
	assign B_DAC[11] = w2958;
	assign B_DAC[12] = w2957;
	assign B_DAC[13] = w2956;
	assign B_DAC[14] = w2955;
	assign B_DAC[15] = w2953;
	assign B_DAC[16] = w2954;
	assign nOE1 = nOE1;
	assign nWE0 = nWE0;
	assign nWE1 = nWE1;
	assign nCAS1 = nCAS1;
	assign nRAS1 = nRAS1;
	assign AD_RD_DIR = AD_RD_DIR;
	assign nYS = nYS;
	assign nSC = w2618;
	assign nSE0_1 = w2507;
	assign ADo[7] = w2466;
	assign ADo[6] = w2474;
	assign ADo[5] = w2655;
	assign ADo[4] = w2482;
	assign ADo[3] = w2596;
	assign ADo[2] = w2595;
	assign ADo[1] = w2544;
	assign ADo[0] = w2711;
	assign RDo[6] = w2656;
	assign RDo[5] = w2686;
	assign RDo[4] = w2661;
	assign RDo[3] = w2660;
	assign RDo[2] = w2688;
	assign RDo[1] = w2712;
	assign RDo[0] = w2514;
	assign w2557 = RDi[6];
	assign w2467 = RDi[7];
	assign w2481 = RDi[4];
	assign w2699 = RDi[5];
	assign w2549 = RDi[2];
	assign w2558 = RDi[3];
	assign w2689 = RDi[0];
	assign w2594 = RDi[1];
	assign w2475 = ADi[6];
	assign w2659 = ADi[7];
	assign w2500 = ADi[4];
	assign w2687 = ADi[5];
	assign w2543 = ADi[2];
	assign w2548 = ADi[3];
	assign w2515 = ADi[0];
	assign w2535 = ADi[1];
	assign RDo[7] = w2658;
	assign w5298 = SD[7];
	assign w5299 = SD[6];
	assign w6728 = SD[5];
	assign w6730 = SD[4];
	assign w5300 = SD[3];
	assign w5297 = SD[2];
	assign w6729 = SD[1];
	assign w5296 = SD[0];
	assign CLK1 = 68K CPU CLOCK;
	assign CLK0 = w1413;
	assign w4498 = EDCLKi;
	assign EDCLKo = EDCLK_O;
	assign w4474 = MCLK;
	assign SUB_CLK = w4463;
	assign w4516 = nRES_PAD;
	assign w1441 = 68kCLKi;
	assign EDCLKd = w1497;
	assign CA_PAD_DIR = w2463;
	assign DB_PAD_DIR = w2464;
	assign w407 = SEL0_M3;
	assign w6734 = nPAL;
	assign w441 = nHL;
	assign SPA/Bo = w2838;
	assign w2781 = SPA/Bi;

	// Instances

	vdp_slatch g1 (.nQ(w355), .D(VPOS[7]), .C(w1568), .nC(w1569) );
	vdp_slatch g2 (.nQ(w1531), .D(HPOS[8]), .C(w376), .nC(w377) );
	vdp_slatch g3 (.nQ(w360), .D(w301), .C(w1470), .nC(w378) );
	vdp_slatch g4 (.D(w302), .C(w1566), .nC(w1567), .nQ(w6836) );
	vdp_slatch g5 (.nQ(w361), .D(w362), .C(w1564), .nC(w1565) );
	vdp_slatch g6 (.nQ(w304), .D(w305), .C(w1562), .nC(w1563) );
	vdp_slatch g7 (.nQ(w363), .D(w362), .C(w379), .nC(w380) );
	vdp_slatch g8 (.nQ(w366), .D(w305), .C(w381), .nC(w382) );
	vdp_slatch g9 (.nQ(w364), .D(w362), .C(w430), .nC(w1467) );
	vdp_slatch g10 (.nQ(w367), .D(w305), .C(w1466), .nC(w387) );
	vdp_slatch g11 (.nQ(w365), .D(w362), .C(w385), .nC(w384) );
	vdp_slatch g12 (.nQ(w307), .D(w305), .C(w383), .nC(w1465) );
	vdp_slatch g13 (.Q(w305), .D(w160), .C(w369), .nC(w368) );
	vdp_slatch g14 (.Q(w362), .D(w934), .C(w372), .nC(w371) );
	vdp_sr_bit g15 (.D(w308), .C2(HCLK2), .C1(HCLK1), .Q(FIFOo[7]), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g16 (.A(1'b1), .nZ(w160), .nE(w1464) );
	vdp_notif0 g17 (.A(w307), .nZ(w308), .nE(w2030) );
	vdp_notif0 g18 (.A(w365), .nZ(w359), .nE(w386) );
	vdp_notif0 g19 (.A(w306), .nZ(AD_DATA[7]), .nE(w1609) );
	vdp_notif0 g20 (.A(w367), .nZ(w308), .nE(w1561) );
	vdp_notif0 g21 (.A(w364), .nZ(w359), .nE(w1608) );
	vdp_notif0 g22 (.A(w1537), .nZ(AD_DATA[7]), .nE(w404) );
	vdp_notif0 g23 (.A(w366), .nZ(w308), .nE(w403) );
	vdp_notif0 g24 (.A(w363), .nZ(w359), .nE(w1468) );
	vdp_notif0 g25 (.A(w1536), .nZ(AD_DATA[7]), .nE(w418) );
	vdp_notif0 g26 (.A(w304), .nZ(w308), .nE(w396) );
	vdp_notif0 g27 (.A(w303), .nZ(AD_DATA[7]), .nE(w416) );
	vdp_notif0 g28 (.A(w360), .nZ(w160), .nE(w1606) );
	vdp_notif0 g29 (.nZ(w358), .nE(w397), .A(w6836) );
	vdp_notif0 g30 (.A(w361), .nZ(w359), .nE(w1607) );
	vdp_notif0 g31 (.A(w355), .nZ(w358), .nE(w1605) );
	vdp_notif0 g32 (.A(w433), .nZ(w160), .nE(w398) );
	vdp_aon22 g33 (.Z(w433), .A1(w1531), .A2(w1570), .B1(w402), .B2(w355) );
	vdp_aon22 g34 (.A2(w400), .B1(w401), .B2(AD_DATA[7]), .A1(w359), .Z(w301) );
	vdp_aon22 g35 (.A2(w6742), .B1(w6743), .B2(w359), .A1(AD_DATA[7]), .Z(w302) );
	vdp_aon22 g36 (.Z(w303), .A2(w399), .B1(w1571), .B2(w304), .A1(w361) );
	vdp_aon22 g37 (.Z(w1536), .A2(w423), .B1(w422), .B2(w363), .A1(w366) );
	vdp_aon22 g38 (.Z(w1537), .A2(w431), .B1(w432), .B2(w364), .A1(w367) );
	vdp_aon22 g39 (.Z(w306), .A2(w6738), .B1(w6739), .B2(w307), .A1(w365) );
	vdp_aon22 g40 (.Z(w934), .A1(w358), .A2(w370), .B1(w374), .B2(w160) );
	vdp_slatch g41 (.nQ(w223), .D(VPOS[6]), .C(w1568), .nC(w1569) );
	vdp_slatch g42 (.nQ(w225), .D(HPOS[7]), .C(w376), .nC(w377) );
	vdp_slatch g43 (.nQ(w227), .D(w263), .C(w1470), .nC(w378) );
	vdp_slatch g44 (.nQ(w265), .D(w1437), .C(w1566), .nC(w1567) );
	vdp_slatch g45 (.nQ(w228), .D(w229), .C(w1564), .nC(w1565) );
	vdp_slatch g46 (.nQ(w267), .D(w268), .C(w1562), .nC(w1563) );
	vdp_slatch g47 (.nQ(w230), .D(w229), .C(w379), .nC(w380) );
	vdp_slatch g48 (.nQ(w232), .D(w268), .C(w381), .nC(w382) );
	vdp_slatch g49 (.nQ(w233), .D(w229), .C(w430), .nC(w1467) );
	vdp_slatch g50 (.nQ(w235), .D(w268), .C(w1466), .nC(w387) );
	vdp_slatch g51 (.nQ(w236), .D(w229), .C(w385), .nC(w384) );
	vdp_slatch g52 (.nQ(w270), .D(w268), .C(w383), .nC(w1465) );
	vdp_slatch g53 (.Q(w268), .D(DB[6]), .C(w369), .nC(w368) );
	vdp_slatch g54 (.Q(w229), .D(w271), .C(w372), .nC(w371) );
	vdp_sr_bit g55 (.D(w264), .Q(FIFOo[6]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g56 (.A(1'b1), .nZ(DB[6]), .nE(w1464) );
	vdp_notif0 g57 (.A(w270), .nZ(w264), .nE(w2030) );
	vdp_notif0 g58 (.A(w236), .nZ(RD_DATA[6]), .nE(w386) );
	vdp_notif0 g59 (.A(w269), .nZ(AD_DATA[6]), .nE(w1609) );
	vdp_notif0 g60 (.A(w235), .nZ(w264), .nE(w1561) );
	vdp_notif0 g61 (.A(w233), .nZ(RD_DATA[6]), .nE(w1608) );
	vdp_notif0 g62 (.A(w234), .nZ(AD_DATA[6]), .nE(w404) );
	vdp_notif0 g63 (.A(w232), .nZ(w264), .nE(w403) );
	vdp_notif0 g64 (.A(w230), .nZ(RD_DATA[6]), .nE(w1468) );
	vdp_notif0 g65 (.A(w231), .nZ(AD_DATA[6]), .nE(w418) );
	vdp_notif0 g66 (.A(w267), .nZ(w264), .nE(w396) );
	vdp_notif0 g67 (.A(w266), .nZ(AD_DATA[6]), .nE(w416) );
	vdp_notif0 g68 (.A(w227), .nZ(DB[6]), .nE(w1606) );
	vdp_notif0 g69 (.A(w265), .nZ(DB[14]), .nE(w397) );
	vdp_notif0 g70 (.A(w228), .nZ(RD_DATA[6]), .nE(w1607) );
	vdp_notif0 g71 (.A(w223), .nZ(DB[14]), .nE(w1605) );
	vdp_notif0 g72 (.A(w226), .nZ(DB[6]), .nE(w398) );
	vdp_aon22 g73 (.A2(w1570), .B1(w402), .B2(w223), .A1(w225), .Z(w226) );
	vdp_aon22 g74 (.Z(w263), .A2(w400), .B1(w401), .B2(AD_DATA[6]), .A1(RD_DATA[6]) );
	vdp_aon22 g75 (.Z(w1437), .A2(w6742), .B1(w6743), .B2(RD_DATA[6]), .A1(AD_DATA[6]) );
	vdp_aon22 g76 (.Z(w266), .A2(w399), .B1(w1571), .B2(w267), .A1(w228) );
	vdp_aon22 g77 (.Z(w231), .A2(w423), .B1(w422), .B2(w232), .A1(w230) );
	vdp_aon22 g78 (.Z(w234), .A2(w431), .B1(w432), .B2(w235), .A1(w233) );
	vdp_aon22 g79 (.Z(w269), .A2(w6738), .B1(w6739), .B2(w270), .A1(w236) );
	vdp_aon22 g80 (.Z(w271), .A1(DB[14]), .A2(w370), .B1(w374), .B2(DB[6]) );
	vdp_slatch g81 (.nQ(w339), .D(VPOS[5]), .C(w1568), .nC(w1569) );
	vdp_slatch g82 (.nQ(w1532), .D(HPOS[6]), .C(w376), .nC(w377) );
	vdp_slatch g83 (.nQ(w344), .D(w292), .C(w1470), .nC(w378) );
	vdp_slatch g84 (.D(w293), .C(w1566), .nC(w1567), .nQ(w6837) );
	vdp_slatch g85 (.nQ(w345), .D(w351), .C(w1564), .nC(w1565) );
	vdp_slatch g86 (.nQ(w295), .D(w296), .C(w1562), .nC(w1563) );
	vdp_slatch g87 (.nQ(w347), .D(w351), .C(w379), .nC(w380) );
	vdp_slatch g88 (.nQ(w346), .D(w296), .C(w381), .nC(w382) );
	vdp_slatch g89 (.nQ(w349), .D(w351), .C(w430), .nC(w1467) );
	vdp_slatch g90 (.nQ(w352), .D(w296), .C(w1466), .nC(w387) );
	vdp_slatch g91 (.nQ(w353), .D(w351), .C(w385), .nC(w384) );
	vdp_slatch g92 (.nQ(w298), .D(w296), .C(w383), .nC(w1465) );
	vdp_slatch g93 (.Q(w296), .D(DB[5]), .C(w369), .nC(w368) );
	vdp_slatch g94 (.Q(w351), .D(w299), .C(w372), .nC(w371) );
	vdp_sr_bit g95 (.D(w300), .Q(FIFOo[5]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g96 (.A(1'b1), .nZ(DB[5]), .nE(w1464) );
	vdp_notif0 g97 (.A(w298), .nZ(w300), .nE(w2030) );
	vdp_notif0 g98 (.A(w353), .nZ(RD_DATA[5]), .nE(w386) );
	vdp_notif0 g99 (.A(w297), .nZ(w291), .nE(w1609) );
	vdp_notif0 g100 (.A(w352), .nZ(w300), .nE(w1561) );
	vdp_notif0 g101 (.A(w349), .nZ(RD_DATA[5]), .nE(w1608) );
	vdp_notif0 g102 (.A(w350), .nZ(w291), .nE(w404) );
	vdp_notif0 g103 (.A(w346), .nZ(w300), .nE(w403) );
	vdp_notif0 g104 (.A(w347), .nZ(RD_DATA[5]), .nE(w1468) );
	vdp_notif0 g105 (.A(w348), .nZ(w291), .nE(w418) );
	vdp_notif0 g106 (.A(w295), .nZ(w300), .nE(w396) );
	vdp_notif0 g107 (.A(w294), .nZ(w291), .nE(w416) );
	vdp_notif0 g108 (.A(w344), .nZ(DB[5]), .nE(w1606) );
	vdp_notif0 g109 (.nZ(DB[13]), .nE(w397), .A(w6837) );
	vdp_notif0 g110 (.A(w345), .nZ(RD_DATA[5]), .nE(w1607) );
	vdp_notif0 g111 (.A(w339), .nZ(DB[13]), .nE(w1605) );
	vdp_notif0 g112 (.A(w343), .nZ(DB[5]), .nE(w398) );
	vdp_aon22 g113 (.Z(w343), .A1(w1532), .A2(w1570), .B1(w402), .B2(w339) );
	vdp_aon22 g114 (.A2(w400), .B1(w401), .B2(w291), .A1(RD_DATA[5]), .Z(w292) );
	vdp_aon22 g115 (.A2(w6742), .B1(w6743), .B2(RD_DATA[5]), .A1(w291), .Z(w293) );
	vdp_aon22 g116 (.Z(w294), .A2(w399), .B1(w1571), .B2(w295), .A1(w345) );
	vdp_aon22 g117 (.Z(w348), .A2(w423), .B1(w422), .B2(w347), .A1(w346) );
	vdp_aon22 g118 (.Z(w350), .A2(w431), .B1(w432), .B2(w349), .A1(w352) );
	vdp_aon22 g119 (.Z(w297), .A2(w6738), .B1(w6739), .B2(w298), .A1(w353) );
	vdp_aon22 g120 (.Z(w299), .A1(DB[13]), .A2(w370), .B1(w374), .B2(DB[5]) );
	vdp_slatch g121 (.nQ(w208), .D(VPOS[4]), .C(w1568), .nC(w1569) );
	vdp_slatch g122 (.nQ(w210), .D(HPOS[5]), .C(w376), .nC(w377) );
	vdp_slatch g123 (.nQ(w1572), .D(w255), .C(w1470), .nC(w378) );
	vdp_slatch g124 (.D(w1535), .C(w1566), .nC(w1567), .nQ(w6838) );
	vdp_slatch g125 (.nQ(w212), .D(w213), .C(w1564), .nC(w1565) );
	vdp_slatch g126 (.nQ(w258), .D(w259), .C(w1562), .nC(w1563) );
	vdp_slatch g127 (.nQ(w214), .D(w213), .C(w379), .nC(w380) );
	vdp_slatch g128 (.nQ(w216), .D(w259), .C(w381), .nC(w382) );
	vdp_slatch g129 (.nQ(w217), .D(w213), .C(w430), .nC(w1467) );
	vdp_slatch g130 (.nQ(w219), .D(w259), .C(w1466), .nC(w387) );
	vdp_slatch g131 (.nQ(w220), .D(w213), .C(w385), .nC(w384) );
	vdp_slatch g132 (.nQ(w261), .D(w259), .C(w383), .nC(w1465) );
	vdp_slatch g133 (.Q(w259), .D(DB[4]), .C(w369), .nC(w368) );
	vdp_slatch g134 (.Q(w213), .D(w262), .C(w372), .nC(w371) );
	vdp_sr_bit g135 (.D(w256), .Q(FIFOo[4]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g136 (.A(1'b1), .nZ(DB[4]), .nE(w1464) );
	vdp_notif0 g137 (.A(w261), .nZ(w256), .nE(w2030) );
	vdp_notif0 g138 (.A(w220), .nZ(RD_DATA[4]), .nE(w386) );
	vdp_notif0 g139 (.A(w260), .nZ(AD_DATA[4]), .nE(w1609) );
	vdp_notif0 g140 (.A(w219), .nZ(w256), .nE(w1561) );
	vdp_notif0 g141 (.A(w217), .nZ(RD_DATA[4]), .nE(w1608) );
	vdp_notif0 g142 (.A(w218), .nZ(AD_DATA[4]), .nE(w404) );
	vdp_notif0 g143 (.A(w216), .nZ(w256), .nE(w403) );
	vdp_notif0 g144 (.A(w214), .nZ(RD_DATA[4]), .nE(w1468) );
	vdp_notif0 g145 (.A(w215), .nZ(AD_DATA[4]), .nE(w418) );
	vdp_notif0 g146 (.A(w258), .nZ(w256), .nE(w396) );
	vdp_notif0 g147 (.A(w257), .nZ(AD_DATA[4]), .nE(w416) );
	vdp_notif0 g148 (.A(w1572), .nZ(DB[4]), .nE(w1606) );
	vdp_notif0 g149 (.nZ(DB[12]), .nE(w397), .A(w6838) );
	vdp_notif0 g150 (.A(w212), .nZ(RD_DATA[4]), .nE(w1607) );
	vdp_notif0 g151 (.A(w208), .nZ(DB[12]), .nE(w1605) );
	vdp_notif0 g152 (.A(w211), .nZ(DB[4]), .nE(w398) );
	vdp_aon22 g153 (.A2(w1570), .B1(w402), .B2(w208), .A1(w210), .Z(w211) );
	vdp_aon22 g154 (.Z(w255), .A2(w400), .B1(w401), .B2(AD_DATA[4]), .A1(RD_DATA[4]) );
	vdp_aon22 g155 (.Z(w1535), .A2(w6742), .B1(w6743), .B2(RD_DATA[4]), .A1(AD_DATA[4]) );
	vdp_aon22 g156 (.Z(w257), .A2(w399), .B1(w1571), .B2(w258), .A1(w212) );
	vdp_aon22 g157 (.Z(w215), .A2(w423), .B1(w422), .B2(w216), .A1(w214) );
	vdp_aon22 g158 (.Z(w218), .A2(w431), .B1(w432), .B2(w219), .A1(w217) );
	vdp_aon22 g159 (.Z(w260), .A2(w6738), .B1(w6739), .B2(w261), .A1(w220) );
	vdp_aon22 g160 (.Z(w262), .A1(DB[12]), .A2(w370), .B1(w374), .B2(DB[4]) );
	vdp_slatch g161 (.nQ(w322), .D(VPOS[3]), .C(w1568), .nC(w1569) );
	vdp_slatch g162 (.nQ(w1533), .D(HPOS[4]), .C(w376), .nC(w377) );
	vdp_slatch g163 (.nQ(w328), .D(w282), .C(w1470), .nC(w378) );
	vdp_slatch g164 (.D(w283), .C(w1566), .nC(w1567), .nQ(w6839) );
	vdp_slatch g165 (.nQ(w329), .D(w332), .C(w1564), .nC(w1565) );
	vdp_slatch g166 (.nQ(w285), .D(w286), .C(w1562), .nC(w1563) );
	vdp_slatch g167 (.nQ(w330), .D(w332), .C(w379), .nC(w380) );
	vdp_slatch g168 (.nQ(w331), .D(w286), .C(w381), .nC(w382) );
	vdp_slatch g169 (.nQ(w334), .D(w332), .C(w430), .nC(w1467) );
	vdp_slatch g170 (.nQ(w336), .D(w286), .C(w1466), .nC(w387) );
	vdp_slatch g171 (.nQ(w337), .D(w332), .C(w385), .nC(w384) );
	vdp_slatch g172 (.nQ(w288), .D(w286), .C(w383), .nC(w1465) );
	vdp_slatch g173 (.Q(w286), .D(w156), .C(w369), .nC(w368) );
	vdp_slatch g174 (.Q(w332), .D(w289), .C(w372), .nC(w371) );
	vdp_sr_bit g175 (.D(w290), .Q(FIFOo[3]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g176 (.A(1'b1), .nZ(w156), .nE(w1464) );
	vdp_notif0 g177 (.A(w288), .nZ(w290), .nE(w2030) );
	vdp_notif0 g178 (.A(w337), .nZ(w324), .nE(w386) );
	vdp_notif0 g179 (.A(w287), .nZ(AD_DATA[3]), .nE(w1609) );
	vdp_notif0 g180 (.A(w336), .nZ(w290), .nE(w1561) );
	vdp_notif0 g181 (.A(w334), .nZ(w324), .nE(w1608) );
	vdp_notif0 g182 (.A(w335), .nZ(AD_DATA[3]), .nE(w404) );
	vdp_notif0 g183 (.A(w331), .nZ(w290), .nE(w403) );
	vdp_notif0 g184 (.A(w330), .nZ(w324), .nE(w1468) );
	vdp_notif0 g185 (.A(w333), .nZ(AD_DATA[3]), .nE(w418) );
	vdp_notif0 g186 (.A(w285), .nZ(w290), .nE(w396) );
	vdp_notif0 g187 (.A(w284), .nZ(AD_DATA[3]), .nE(w416) );
	vdp_notif0 g188 (.A(w328), .nZ(w156), .nE(w1606) );
	vdp_notif0 g189 (.nZ(w325), .nE(w397), .A(w6839) );
	vdp_notif0 g190 (.A(w329), .nZ(w324), .nE(w1607) );
	vdp_notif0 g191 (.A(w322), .nZ(w325), .nE(w1605) );
	vdp_notif0 g192 (.A(w327), .nZ(w156), .nE(w398) );
	vdp_aon22 g193 (.Z(w327), .A1(w1533), .A2(w1570), .B1(w402), .B2(w322) );
	vdp_aon22 g194 (.A2(w400), .B1(w401), .B2(AD_DATA[3]), .A1(w324), .Z(w282) );
	vdp_aon22 g195 (.A2(w6742), .B1(w6743), .B2(w324), .A1(AD_DATA[3]), .Z(w283) );
	vdp_aon22 g196 (.Z(w284), .A2(w399), .B1(w1571), .B2(w285), .A1(w329) );
	vdp_aon22 g197 (.Z(w333), .A2(w423), .B1(w422), .B2(w330), .A1(w331) );
	vdp_aon22 g198 (.Z(w335), .A2(w431), .B1(w432), .B2(w334), .A1(w336) );
	vdp_aon22 g199 (.Z(w287), .A2(w6738), .B1(w6739), .B2(w288), .A1(w337) );
	vdp_aon22 g200 (.Z(w289), .A1(w325), .A2(w370), .B1(w374), .B2(w156) );
	vdp_slatch g201 (.nQ(w193), .D(VPOS[2]), .C(w1568), .nC(w1569) );
	vdp_slatch g202 (.nQ(w1573), .D(HPOS[3]), .C(w376), .nC(w377) );
	vdp_slatch g203 (.nQ(w195), .D(w246), .C(w1470), .nC(w378) );
	vdp_slatch g204 (.D(w1471), .C(w1566), .nC(w1567), .nQ(w6840) );
	vdp_slatch g205 (.nQ(w196), .D(w199), .C(w1564), .nC(w1565) );
	vdp_slatch g206 (.nQ(w249), .D(w250), .C(w1562), .nC(w1563) );
	vdp_slatch g207 (.nQ(w197), .D(w199), .C(w379), .nC(w380) );
	vdp_slatch g208 (.nQ(w200), .D(w250), .C(w381), .nC(w382) );
	vdp_slatch g209 (.nQ(w201), .D(w199), .C(w430), .nC(w1467) );
	vdp_slatch g210 (.nQ(w203), .D(w250), .C(w1466), .nC(w387) );
	vdp_slatch g211 (.nQ(w204), .D(w199), .C(w385), .nC(w384) );
	vdp_slatch g212 (.nQ(w252), .D(w250), .C(w383), .nC(w1465) );
	vdp_slatch g213 (.Q(w250), .D(DB[2]), .C(w369), .nC(w368) );
	vdp_slatch g214 (.Q(w199), .D(w253), .C(w372), .nC(w371) );
	vdp_sr_bit g215 (.D(w247), .Q(FIFOo[2]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g216 (.A(w205), .nZ(DB[2]), .nE(w1464) );
	vdp_notif0 g217 (.A(w252), .nZ(w247), .nE(w2030) );
	vdp_notif0 g218 (.A(w204), .nZ(RD_DATA[2]), .nE(w386) );
	vdp_notif0 g219 (.A(w251), .nZ(AD_DATA[2]), .nE(w1609) );
	vdp_notif0 g220 (.A(w203), .nZ(w247), .nE(w1561) );
	vdp_notif0 g221 (.A(w201), .nZ(RD_DATA[2]), .nE(w1608) );
	vdp_notif0 g222 (.A(w202), .nZ(AD_DATA[2]), .nE(w404) );
	vdp_notif0 g223 (.A(w200), .nZ(w247), .nE(w403) );
	vdp_notif0 g224 (.A(w197), .nZ(RD_DATA[2]), .nE(w1468) );
	vdp_notif0 g225 (.A(w198), .nZ(AD_DATA[2]), .nE(w418) );
	vdp_notif0 g226 (.A(w249), .nZ(w247), .nE(w396) );
	vdp_notif0 g227 (.A(w248), .nZ(AD_DATA[2]), .nE(w416) );
	vdp_notif0 g228 (.A(w195), .nZ(DB[2]), .nE(w1606) );
	vdp_notif0 g229 (.nZ(DB[10]), .nE(w397), .A(w6840) );
	vdp_notif0 g230 (.A(w196), .nZ(RD_DATA[2]), .nE(w1607) );
	vdp_notif0 g231 (.A(w193), .nZ(DB[10]), .nE(w1605) );
	vdp_notif0 g232 (.A(w194), .nZ(DB[2]), .nE(w398) );
	vdp_aon22 g233 (.A2(w1570), .B1(w402), .B2(w193), .A1(w1573), .Z(w194) );
	vdp_aon22 g234 (.Z(w246), .A2(w400), .B1(w401), .B2(AD_DATA[2]), .A1(RD_DATA[2]) );
	vdp_aon22 g235 (.Z(w1471), .A2(w6742), .B1(w6743), .B2(RD_DATA[2]), .A1(AD_DATA[2]) );
	vdp_aon22 g236 (.Z(w248), .A2(w399), .B1(w1571), .B2(w249), .A1(w196) );
	vdp_aon22 g237 (.Z(w198), .A2(w423), .B1(w422), .B2(w200), .A1(w197) );
	vdp_aon22 g238 (.Z(w202), .A2(w431), .B1(w432), .B2(w203), .A1(w201) );
	vdp_aon22 g239 (.Z(w251), .A2(w6738), .B1(w6739), .B2(w252), .A1(w204) );
	vdp_aon22 g240 (.Z(w253), .A1(DB[10]), .A2(w370), .B1(w374), .B2(DB[2]) );
	vdp_slatch g241 (.nQ(w309), .D(VPOS[1]), .C(w1568), .nC(w1569) );
	vdp_slatch g242 (.nQ(w1534), .D(HPOS[2]), .C(w376), .nC(w377) );
	vdp_slatch g243 (.nQ(w312), .D(w272), .C(w1470), .nC(w378) );
	vdp_slatch g244 (.D(w273), .C(w1566), .nC(w1567), .nQ(w6841) );
	vdp_slatch g245 (.nQ(w313), .D(w316), .C(w1564), .nC(w1565) );
	vdp_slatch g246 (.nQ(w275), .D(w276), .C(w1562), .nC(w1563) );
	vdp_slatch g247 (.nQ(w315), .D(w316), .C(w379), .nC(w380) );
	vdp_slatch g248 (.nQ(w314), .D(w276), .C(w381), .nC(w382) );
	vdp_slatch g249 (.nQ(w318), .D(w316), .C(w430), .nC(w1467) );
	vdp_slatch g250 (.nQ(w320), .D(w276), .C(w1466), .nC(w387) );
	vdp_slatch g251 (.nQ(w321), .D(w316), .C(w385), .nC(w384) );
	vdp_slatch g252 (.nQ(w278), .D(w276), .C(w383), .nC(w1465) );
	vdp_slatch g253 (.Q(w276), .D(DB[1]), .C(w369), .nC(w368) );
	vdp_slatch g254 (.Q(w316), .D(w280), .C(w372), .nC(w371) );
	vdp_sr_bit g255 (.D(w281), .Q(FIFOo[1]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g256 (.A(w1610), .nZ(DB[1]), .nE(w1464) );
	vdp_notif0 g257 (.A(w278), .nZ(w281), .nE(w2030) );
	vdp_notif0 g258 (.A(w321), .nZ(RD_DATA[1]), .nE(w386) );
	vdp_notif0 g259 (.A(w277), .nZ(AD_DATA[1]), .nE(w1609) );
	vdp_notif0 g260 (.A(w320), .nZ(w281), .nE(w1561) );
	vdp_notif0 g261 (.A(w318), .nZ(RD_DATA[1]), .nE(w1608) );
	vdp_notif0 g262 (.A(w319), .nZ(AD_DATA[1]), .nE(w404) );
	vdp_notif0 g263 (.A(w314), .nZ(w281), .nE(w403) );
	vdp_notif0 g264 (.A(w315), .nZ(RD_DATA[1]), .nE(w1468) );
	vdp_notif0 g265 (.A(w317), .nZ(AD_DATA[1]), .nE(w418) );
	vdp_notif0 g266 (.A(w275), .nZ(w281), .nE(w396) );
	vdp_notif0 g267 (.A(w274), .nZ(AD_DATA[1]), .nE(w416) );
	vdp_notif0 g268 (.A(w312), .nZ(DB[1]), .nE(w1606) );
	vdp_notif0 g269 (.nZ(DB[9]), .nE(w397), .A(w6841) );
	vdp_notif0 g270 (.A(w313), .nZ(RD_DATA[1]), .nE(w1607) );
	vdp_notif0 g271 (.A(w309), .nZ(DB[9]), .nE(w1605) );
	vdp_notif0 g272 (.A(w1469), .nZ(DB[1]), .nE(w398) );
	vdp_aon22 g273 (.Z(w1469), .A1(w1534), .A2(w1570), .B1(w402), .B2(w309) );
	vdp_aon22 g274 (.A2(w400), .B1(w401), .B2(AD_DATA[1]), .A1(RD_DATA[1]), .Z(w272) );
	vdp_aon22 g275 (.A2(w6742), .B1(w6743), .B2(RD_DATA[1]), .A1(AD_DATA[1]), .Z(w273) );
	vdp_aon22 g276 (.Z(w274), .A2(w399), .B1(w1571), .B2(w275), .A1(w313) );
	vdp_aon22 g277 (.Z(w317), .A2(w423), .B1(w422), .B2(w315), .A1(w314) );
	vdp_aon22 g278 (.Z(w319), .A2(w431), .B1(w432), .B2(w318), .A1(w320) );
	vdp_aon22 g279 (.Z(w277), .A2(w6738), .B1(w6739), .B2(w278), .A1(w321) );
	vdp_aon22 g280 (.Z(w280), .A1(DB[9]), .A2(w370), .B1(w374), .B2(DB[1]) );
	vdp_slatch g281 (.nQ(w178), .D(w176), .C(w1568), .nC(w1569) );
	vdp_slatch g282 (.D(HPOS[1]), .nQ(w1463), .C(w376), .nC(w377) );
	vdp_slatch g283 (.nQ(w180), .D(w238), .C(w1470), .nC(w378) );
	vdp_slatch g284 (.D(w1438), .C(w1566), .nC(w1567), .nQ(w6842) );
	vdp_slatch g285 (.nQ(w181), .D(w185), .C(w1564), .nC(w1565) );
	vdp_slatch g286 (.nQ(w241), .D(w242), .C(w1562), .nC(w1563) );
	vdp_slatch g287 (.nQ(w182), .D(w185), .C(w379), .nC(w380) );
	vdp_slatch g288 (.nQ(w184), .D(w242), .C(w381), .nC(w382) );
	vdp_slatch g289 (.nQ(w186), .D(w185), .C(w430), .nC(w1467) );
	vdp_slatch g290 (.nQ(w188), .D(w242), .C(w1466), .nC(w387) );
	vdp_slatch g291 (.nQ(w189), .D(w185), .C(w385), .nC(w384) );
	vdp_slatch g292 (.nQ(w244), .D(w242), .C(w383), .nC(w1465) );
	vdp_slatch g293 (.Q(w242), .D(DB[0]), .C(w369), .nC(w368) );
	vdp_slatch g294 (.D(w245), .Q(w185), .C(w372), .nC(w371) );
	vdp_sr_bit g295 (.D(w239), .C2(HCLK2), .C1(HCLK1), .Q(FIFOo[0]), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g296 (.A(1'b1), .nZ(DB[0]), .nE(w1464) );
	vdp_notif0 g297 (.A(w244), .nZ(w239), .nE(w2030) );
	vdp_notif0 g298 (.A(w189), .nZ(RD_DATA[0]), .nE(w386) );
	vdp_notif0 g299 (.A(w243), .nZ(AD_DATA[0]), .nE(w1609) );
	vdp_notif0 g300 (.A(w188), .nZ(w239), .nE(w1561) );
	vdp_notif0 g301 (.A(w186), .nZ(RD_DATA[0]), .nE(w1608) );
	vdp_notif0 g302 (.A(w187), .nZ(AD_DATA[0]), .nE(w404) );
	vdp_notif0 g303 (.A(w184), .nZ(w239), .nE(w403) );
	vdp_notif0 g304 (.A(w182), .nZ(RD_DATA[0]), .nE(w1468) );
	vdp_notif0 g305 (.A(w183), .nZ(AD_DATA[0]), .nE(w418) );
	vdp_notif0 g306 (.A(w241), .nZ(w239), .nE(w396) );
	vdp_notif0 g307 (.A(w240), .nZ(AD_DATA[0]), .nE(w416) );
	vdp_notif0 g308 (.A(w180), .nZ(DB[0]), .nE(w1606) );
	vdp_notif0 g309 (.nZ(DB[8]), .nE(w397), .A(w6842) );
	vdp_notif0 g310 (.A(w181), .nZ(RD_DATA[0]), .nE(w1607) );
	vdp_notif0 g311 (.A(w178), .nZ(DB[8]), .nE(w1605) );
	vdp_notif0 g312 (.A(w179), .nZ(DB[0]), .nE(w398) );
	vdp_aon22 g313 (.A2(w1570), .B1(w402), .B2(w178), .A1(w1463), .Z(w179) );
	vdp_aon22 g314 (.Z(w238), .A2(w400), .B1(w401), .B2(AD_DATA[0]), .A1(RD_DATA[0]) );
	vdp_aon22 g315 (.Z(w1438), .A2(w6742), .B1(w6743), .B2(RD_DATA[0]), .A1(AD_DATA[0]) );
	vdp_aon22 g316 (.Z(w240), .A2(w399), .B1(w1571), .B2(w241), .A1(w181) );
	vdp_aon22 g317 (.Z(w183), .A2(w423), .B1(w422), .B2(w184), .A1(w182) );
	vdp_aon22 g318 (.Z(w187), .A2(w431), .B1(w432), .B2(w188), .A1(w186) );
	vdp_aon22 g319 (.Z(w243), .A2(w6738), .B1(w6739), .B2(w244), .A1(w189) );
	vdp_aon22 g320 (.Z(w245), .A1(DB[8]), .A2(w370), .B1(w374), .B2(DB[0]) );
	vdp_not g321 (.A(w279), .nZ(w1610) );
	vdp_not g322 (.A(w254), .nZ(w205) );
	vdp_not g323 (.A(w406), .nZ(w1605) );
	vdp_not g324 (.A(w410), .nZ(w398) );
	vdp_not g325 (.A(w415), .nZ(w1606) );
	vdp_not g326 (.A(w415), .nZ(w397) );
	vdp_sr_bit g327 (.D(w414), .C2(HCLK2), .C1(HCLK1), .Q(w950), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g328 (.D(w460), .Q(w429), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g329 (.D(w429), .Q(w426), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g330 (.D(w426), .Q(w420), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g331 (.D(w424), .Q(w466), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g332 (.D(w466), .Q(w421), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g333 (.D(w467), .Q(w414), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g334 (.D(w417), .Q(w411), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g335 (.A(w449), .nZ(w1607) );
	vdp_not g336 (.A(w449), .nZ(w416) );
	vdp_not g337 (.A(w449), .nZ(w396) );
	vdp_not g338 (.A(w451), .nZ(w1468) );
	vdp_not g339 (.A(w451), .nZ(w418) );
	vdp_not g340 (.A(w451), .nZ(w403) );
	vdp_not g341 (.A(w463), .nZ(w1608) );
	vdp_not g342 (.A(w463), .nZ(w404) );
	vdp_not g343 (.A(w463), .nZ(w1561) );
	vdp_not g344 (.A(w452), .nZ(w386) );
	vdp_not g345 (.A(w452), .nZ(w1609) );
	vdp_not g346 (.A(w452), .nZ(w2030) );
	vdp_not g347 (.A(w428), .nZ(w1464) );
	vdp_not g348 (.A(w426), .nZ(w405) );
	vdp_not g349 (.A(w407), .nZ(w408) );
	vdp_comp_str g350 (.A(w442), .Z(w1568), .nZ(w1569) );
	vdp_comp_str g351 (.A(w443), .Z(w376), .nZ(w377) );
	vdp_comp_str g352 (.A(w412), .Z(w1470), .nZ(w378) );
	vdp_comp_str g353 (.A(w413), .Z(w1566), .nZ(w1567) );
	vdp_comp_str g354 (.A(w468), .Z(w1564), .nZ(w1565) );
	vdp_comp_str g355 (.A(w468), .Z(w1562), .nZ(w1563) );
	vdp_comp_str g356 (.A(w465), .Z(w379), .nZ(w380) );
	vdp_comp_str g357 (.A(w465), .Z(w381), .nZ(w382) );
	vdp_comp_str g358 (.A(w509), .Z(w430), .nZ(w1467) );
	vdp_comp_str g359 (.A(w509), .Z(w1466), .nZ(w387) );
	vdp_comp_str g360 (.A(w459), .Z(w385), .nZ(w384) );
	vdp_comp_str g361 (.A(w459), .Z(w383), .nZ(w1465) );
	vdp_comp_str g362 (.A(w470), .Z(w369), .nZ(w368) );
	vdp_comp_str g363 (.A(w470), .Z(w372), .nZ(w371) );
	vdp_comp_we g364 (.A(w407), .Z(w370), .nZ(w374) );
	vdp_comp_we g365 (.A(w448), .Z(w6738), .nZ(w6739) );
	vdp_comp_we g366 (.A(w448), .Z(w431), .nZ(w432) );
	vdp_comp_we g367 (.A(w448), .Z(w423), .nZ(w422) );
	vdp_comp_we g368 (.A(w448), .Z(w399), .nZ(w1571) );
	vdp_comp_we g369 (.A(w453), .Z(w6742), .nZ(w6743) );
	vdp_comp_we g370 (.A(w409), .Z(w400), .nZ(w401) );
	vdp_comp_we g371 (.A(w446), .Z(w1570), .nZ(w402) );
	vdp_and g372 (.Z(w412), .B(HCLK1), .A(w411) );
	vdp_and g373 (.Z(w413), .B(HCLK1), .A(w414) );
	vdp_and g374 (.Z(w417), .B(w421), .A(w419) );
	vdp_and g375 (.Z(w467), .B(w421), .A(w425) );
	vdp_nand g376 (.Z(w425), .B(w453), .A(w405) );
	vdp_nand g377 (.Z(w419), .B(w453), .A(w426) );
	vdp_and3 g378 (.Z(w453), .B(w439), .A(w407), .C(w440) );
	vdp_and3 g379 (.Z(w409), .B(w408), .A(w420), .C(128k) );
	vdp_not g380 (.A(128k), .nZ(w440) );
	vdp_sr_bit g381 (.D(w437), .C2(HCLK2), .C1(HCLK1), .Q(w436), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g382 (.D(w1447), .Q(w474), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g383 (.D(w1526), .C2(HCLK2), .C1(HCLK1), .Q(w500), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g384 (.A(w501), .nZ(w427) );
	vdp_fa g385 (.SUM(w461), .A(w500), .B(1'b0), .CI(w502) );
	vdp_not g386 (.A(w437), .nZ(w435) );
	vdp_not g387 (.A(M5), .nZ(w473) );
	vdp_not g388 (.A(w445), .nZ(w443) );
	vdp_not g389 (.A(w455), .nZ(w456) );
	vdp_not g390 (.A(w507), .nZ(w458) );
	vdp_not g391 (.A(w500), .nZ(w457) );
	vdp_slatch g392 (.Q(w494), .D(w498), .C(w480), .nC(w434) );
	vdp_slatch g393 (.Q(w1514), .D(w498), .C(w492), .nC(w464) );
	vdp_slatch g394 (.Q(w495), .D(w498), .C(w478), .nC(w450) );
	vdp_slatch g395 (.Q(w496), .D(w498), .C(w476), .nC(w447) );
	vdp_slatch g396 (.Q(w497), .D(w471), .C(w480), .nC(w434) );
	vdp_slatch g397 (.Q(w499), .D(w471), .C(w492), .nC(w464) );
	vdp_slatch g398 (.Q(w1513), .D(w471), .E(w478), .nE(w450) );
	vdp_slatch g399 (.Q(w493), .D(w471), .C(w476), .nC(w447) );
	vdp_slatch g400 (.Q(w485), .D(w472), .C(w480), .nC(w434) );
	vdp_slatch g401 (.Q(w479), .D(w472), .C(w492), .nC(w464) );
	vdp_slatch g402 (.Q(w483), .D(w472), .C(w478), .nC(w450) );
	vdp_slatch g403 (.Q(w486), .D(w472), .C(w476), .nC(w447) );
	vdp_comp_dff g404 (.D(w441), .C2(HCLK2), .C1(HCLK1), .Q(w437), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and g405 (.Z(w1447), .B(w435), .A(w436) );
	vdp_or g406 (.Z(w442), .B(w473), .A(w443) );
	vdp_or g407 (.Z(w446), .B(CA[0]), .A(w407) );
	vdp_and3 g408 (.Z(w449), .B(w501), .A(w457), .C(w507) );
	vdp_and3 g409 (.Z(w451), .B(w501), .A(w458), .C(w500) );
	vdp_and3 g410 (.Z(w452), .B(w457), .A(w458), .C(w501) );
	vdp_xor g411 (.Z(w454), .B(w505), .A(w504) );
	vdp_aon22 g412 (.Z(w448), .A1(w456), .A2(w505), .B1(w524), .B2(w455) );
	vdp_and3 g413 (.Z(w463), .B(w500), .A(w507), .C(w501) );
	vdp_comp_str g414 (.A(w509), .Z(w480), .nZ(w434) );
	vdp_comp_str g415 (.A(w459), .Z(w476), .nZ(w447) );
	vdp_comp_str g416 (.A(w468), .Z(w478), .nZ(w450) );
	vdp_comp_str g417 (.A(w465), .Z(w492), .nZ(w464) );
	vdp_nand g418 (.Z(w455), .B(w506), .A(w454) );
	vdp_and g419 (.Z(w1526), .B(w503), .A(w461) );
	vdp_aoi21 g420 (.Z(w445), .B(w444), .A1(HCLK1), .A2(w474) );
	vdp_nor g421 (.Z(w444), .B(w477), .A(w473) );
	vdp_nor g422 (.Z(w439), .B(w471), .A(w472) );
	vdp_not g423 (.A(w488), .nZ(w551) );
	vdp_not g424 (.A(w487), .nZ(w555) );
	vdp_nor g425 (.Z(w615), .A(w535), .B(w488) );
	vdp_or g426 (.A(w1446), .Z(w489), .B(w490) );
	vdp_comp_we g427 (.A(w1516), .nZ(w481), .Z(w529) );
	vdp_aon22 g428 (.Z(w487), .A1(w529), .A2(w472), .B1(w481), .B2(w491) );
	vdp_aon22 g429 (.Z(w554), .A1(w529), .A2(w514), .B1(w481), .B2(w489) );
	vdp_aon22 g430 (.Z(w544), .A1(w529), .A2(w540), .B1(w481), .B2(w504) );
	vdp_aon22 g431 (.Z(w488), .A1(w529), .A2(w471), .B1(w481), .B2(w536) );
	vdp_aon22 g432 (.Z(w550), .A1(w529), .A2(w534), .B1(w481), .B2(w505) );
	vdp_aon22 g433 (.Z(w535), .A1(w529), .A2(w498), .B1(w481), .B2(w528) );
	vdp_and g434 (.Z(w549), .A(w527), .B(w526) );
	vdp_and g435 (.Z(w484), .A(w527), .B(w507) );
	vdp_and g436 (.Z(w548), .A(w500), .B(w526) );
	vdp_and g437 (.Z(w482), .A(w500), .B(w507) );
	vdp_and g438 (.Z(w1448), .A(w503), .B(w522) );
	vdp_fa g439 (.SUM(w522), .A(w507), .B(w508), .CO(w502), .CI(w523) );
	vdp_sr_bit g440 (.D(w1448), .C2(HCLK2), .C1(HCLK1), .Q(w507), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g441 (.A(w525), .nZ(w1450) );
	vdp_not g442 (.A(w515), .nZ(w518) );
	vdp_and g443 (.Z(w508), .A(w584), .B(w1450) );
	vdp_and3 g444 (.Z(w465), .B(w516), .A(w515), .C(w519) );
	vdp_and3 g445 (.Z(w509), .B(w516), .A(w515), .C(w517) );
	vdp_xor g446 (.Z(w521), .A(w500), .B(w515) );
	vdp_not g447 (.A(w507), .nZ(w526) );
	vdp_not g448 (.A(w500), .nZ(w527) );
	vdp_not g449 (.A(w506), .nZ(w1449) );
	vdp_and5 g450 (.Z(w38), .A(w552), .B(w544), .C(w556), .D(w555), .E(w488) );
	vdp_and5 g451 (.Z(w37), .A(w552), .B(w550), .C(w556), .D(w555), .E(w488) );
	vdp_aon2222 g452 (.C2(w545), .B2(w543), .A2(w542), .C1(w548), .B1(w484), .A1(w549), .Z(w490), .D2(w546), .D1(w482) );
	vdp_aon2222 g453 (.C2(w479), .B2(w483), .A2(w486), .C1(w548), .B1(w484), .A1(w549), .Z(w491), .D2(w485), .D1(w482) );
	vdp_aon2222 g454 (.C2(w1461), .B2(w539), .A2(w1462), .C1(w548), .B1(w484), .A1(w549), .Z(w504), .D2(w537), .D1(w482) );
	vdp_aon2222 g455 (.C2(w499), .B2(w1513), .A2(w493), .C1(w548), .B1(w484), .A1(w549), .Z(w536), .D2(w497), .D1(w482) );
	vdp_aon2222 g456 (.C2(w1515), .B2(w533), .A2(w530), .C1(w548), .B1(w484), .A1(w549), .Z(w505), .D2(w547), .D1(w482) );
	vdp_aon2222 g457 (.C2(w1514), .B2(w495), .A2(w496), .C1(w548), .B1(w484), .A1(w549), .Z(w528), .D2(w494), .D1(w482) );
	vdp_nor g458 (.Z(w525), .A(w1449), .B(w454) );
	vdp_or g459 (.Z(w470), .B(w512), .A(w978) );
	vdp_cnt_bit g460 (.R(SYSRES), .Q(w515), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2), .CI(w513) );
	vdp_cnt_bit g461 (.R(SYSRES), .Q(w517), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2), .CI(w577), .CO(w513) );
	vdp_not g462 (.A(w517), .nZ(w519) );
	vdp_not g463 (.A(w1451), .nZ(w516) );
	vdp_and3 g464 (.Z(w459), .B(w516), .A(w518), .C(w519) );
	vdp_and3 g465 (.Z(w468), .B(w516), .A(w518), .C(w517) );
	vdp_xor g466 (.Z(w520), .A(w507), .B(w517) );
	vdp_fa g467 (.SUM(w1575), .A(w585), .B(w524), .CO(w523), .CI(1'b0) );
	vdp_and g468 (.Z(w585), .A(w525), .B(w584) );
	vdp_and g469 (.Z(w1460), .A(w503), .B(w1575) );
	vdp_sr_bit g470 (.D(w1460), .C2(HCLK2), .C1(HCLK1), .Q(w524), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g471 (.A(w1458), .nZ(w570) );
	vdp_comp_str g472 (.A(w459), .Z(w564), .nZ(w541) );
	vdp_comp_str g473 (.A(w468), .Z(w572), .nZ(w531) );
	vdp_comp_str g474 (.A(w465), .Z(w571), .nZ(w538) );
	vdp_comp_str g475 (.A(w509), .Z(w573), .nZ(w532) );
	vdp_slatch g476 (.Q(w547), .D(w534), .C(w573), .nC(w532) );
	vdp_slatch g477 (.Q(w1515), .D(w534), .C(w571), .nC(w538) );
	vdp_slatch g478 (.Q(w533), .D(w534), .C(w572), .nC(w531) );
	vdp_slatch g479 (.Q(w530), .D(w534), .C(w564), .nC(w541) );
	vdp_slatch g480 (.Q(w537), .D(w540), .C(w573), .nC(w532) );
	vdp_slatch g481 (.Q(w1461), .D(w540), .C(w571), .nC(w538) );
	vdp_slatch g482 (.Q(w539), .D(w540), .C(w572), .nC(w531) );
	vdp_slatch g483 (.Q(w1462), .D(w540), .C(w564), .nC(w541) );
	vdp_slatch g484 (.Q(w546), .D(w514), .C(w573), .nC(w532) );
	vdp_slatch g485 (.Q(w545), .D(w514), .C(w571), .nC(w538) );
	vdp_slatch g486 (.Q(w543), .D(w514), .C(w572), .nC(w531) );
	vdp_slatch g487 (.Q(w542), .D(w514), .C(w564), .nC(w541) );
	vdp_and5 g488 (.Z(w175), .A(w552), .B(w544), .C(w555), .D(w535), .E(w551) );
	vdp_and5 g489 (.Z(w174), .A(w552), .B(w550), .C(w555), .D(w535), .E(w551) );
	vdp_not g490 (.A(M5), .nZ(w1446) );
	vdp_not g491 (.A(w535), .nZ(w556) );
	vdp_not g492 (.A(w553), .nZ(w552) );
	vdp_oai21 g493 (.A1(w589), .Z(w553), .A2(w584), .B(w554) );
	vdp_and3 g494 (.Z(w575), .B(w584), .A(w506), .C(w524) );
	vdp_nor g495 (.Z(w1459), .A(w574), .B(w524) );
	vdp_nor g496 (.Z(w582), .A(w521), .B(w520) );
	vdp_aoi21 g497 (.A1(DCLK1), .Z(w1451), .A2(w512), .B(w576) );
	vdp_comb1 g498 (.Z(w1458), .A1(w584), .B(w586), .A2(w1459), .C(HCLK1) );
	vdp_not g499 (.A(w562), .nZ(w35) );
	vdp_not g500 (.A(w1518), .nZ(w557) );
	vdp_not g501 (.A(128k), .nZ(w560) );
	vdp_not g502 (.A(w559), .nZ(w133) );
	vdp_not g503 (.A(w1519), .nZ(w134) );
	vdp_not g504 (.A(w1520), .nZ(w558) );
	vdp_not g505 (.A(VRAMA[0]), .nZ(w1521) );
	vdp_not g506 (.A(w566), .nZ(w565) );
	vdp_not g507 (.A(w500), .nZ(w611) );
	vdp_not g508 (.A(w507), .nZ(w613) );
	vdp_not g509 (.A(w587), .nZ(w610) );
	vdp_not g510 (.A(w407), .nZ(w609) );
	vdp_not g511 (.A(128k), .nZ(w1525) );
	vdp_not g512 (.A(w524), .nZ(w605) );
	vdp_not g513 (.A(SYSRES), .nZ(w503) );
	vdp_not g514 (.A(w593), .nZ(w1453) );
	vdp_not g515 (.A(w34), .nZ(w1452) );
	vdp_not g516 (.A(w583), .nZ(w601) );
	vdp_not g517 (.A(w576), .nZ(w580) );
	vdp_not g518 (.A(w580), .nZ(w581) );
	vdp_sr_bit g519 (.D(w1454), .C2(HCLK2), .C1(HCLK1), .Q(w584), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g520 (.D(w1457), .Q(w589), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_slatch g521 (.Q(w460), .D(VRAMA[0]), .C(w601), .nC(w583) );
	vdp_and g522 (.A(w32), .Z(w1454), .B(w1453) );
	vdp_and g523 (.A(w1452), .Z(w501), .B(w3) );
	vdp_and g524 (.A(w3), .Z(w583), .B(HCLK1) );
	vdp_and g525 (.A(w593), .Z(w34), .B(w591) );
	vdp_and g526 (.A(w592), .Z(w36), .B(w593) );
	vdp_and g527 (.A(w592), .B(w575) );
	vdp_or g528 (.A(w579), .Z(w577), .B(w512) );
	vdp_or g529 (.A(w581), .Z(w949), .B(1'b0) );
	vdp_or g530 (.A(SYSRES), .Z(w603), .B(w596) );
	vdp_and g531 (.A(w584), .Z(w1455), .B(DMA_BUSY) );
	vdp_and g532 (.A(w615), .Z(w506), .B(w1524) );
	vdp_and g533 (.A(w1525), .Z(w1524), .B(w407) );
	vdp_or g534 (.A(w575), .Z(w608), .B(w574) );
	vdp_or g535 (.A(DMA_BUSY), .Z(w1522), .B(w569) );
	vdp_or g536 (.A(DMA_BUSY), .Z(w1523), .B(w568) );
	vdp_and g537 (.A(M5), .Z(w587), .B(w612) );
	vdp_or g538 (.A(w544), .Z(w561), .B(w560) );
	vdp_and g539 (.A(w550), .Z(w1517), .B(128k) );
	vdp_aon22 g540 (.Z(w534), .A2(w1522), .B1(w609), .B2(w587), .A1(w407) );
	vdp_aon22 g541 (.Z(w540), .A2(w1523), .B1(w610), .B2(w609), .A1(w407) );
	vdp_and3 g542 (.A(w32), .Z(w1457), .B(w36), .C(w1456) );
	vdp_rs_ff g543 (.Q(w1456), .R(w603), .S(w1455) );
	vdp_oai21 g544 (.A1(VRAMA[0]), .Z(w566), .A2(128k), .B(w595) );
	vdp_oai21 g545 (.A1(128k), .Z(w1520), .A2(w1521), .B(w595) );
	vdp_aoi21 g546 (.A1(w550), .Z(w1519), .A2(w563), .B(w565) );
	vdp_aoi21 g547 (.A1(w544), .Z(w559), .A2(w563), .B(w558) );
	vdp_aoi21 g548 (.A1(w563), .Z(w1518), .A2(w561), .B(w595) );
	vdp_aoi21 g549 (.A1(w563), .Z(w562), .A2(w1517), .B(w595) );
	vdp_and4 g550 (.A(w552), .Z(w563), .B(w556), .C(w551), .D(w555) );
	vdp_not g551 (.A(w639), .nZ(w1445) );
	vdp_not g552 (.A(w651), .nZ(w650) );
	vdp_and3 g553 (.A(w605), .Z(w606), .B(w641), .C(w650) );
	vdp_and3 g554 (.A(w613), .Z(w628), .B(w616), .C(w611) );
	vdp_and3 g555 (.A(w507), .Z(w632), .B(w616), .C(w611) );
	vdp_and3 g556 (.A(w613), .Z(w621), .B(w616), .C(w500) );
	vdp_and3 g557 (.A(w507), .Z(w625), .B(w616), .C(w500) );
	vdp_or g558 (.A(w607), .Z(w638), .B(w640) );
	vdp_or g559 (.A(w607), .Z(w644), .B(w648) );
	vdp_or g560 (.A(w674), .Z(w594), .B(w647) );
	vdp_and3 g561 (.Z(w592), .B(DMA_BUSY), .A(w673), .C(w646) );
	vdp_or3 g562 (.Z(w598), .B(w589), .A(w595), .C(w645) );
	vdp_and g563 (.A(w599), .Z(w512), .B(w600) );
	vdp_and g564 (.A(w584), .Z(w616), .B(w605) );
	vdp_bufif0 g565 (.A(w597), .Z(VRAMA[8]), .nE(w652) );
	vdp_aoi221 g566 (.Z(w639), .A2(w606), .B1(w593), .B2(w582), .A1(w582), .C(SYSRES) );
	vdp_aon33 g567 (.Z(w675), .A2(w582), .B1(w1555), .B2(w582), .A1(w649), .A3(w1555), .B3(w602) );
	vdp_not g568 (.A(w608), .nZ(w1473) );
	vdp_comp_str g569 (.A(w570), .Z(w1474), .nZ(w635) );
	vdp_not g570 (.A(w632), .nZ(w634) );
	vdp_comp_str g571 (.A(w468), .Z(w1476), .nZ(w1475) );
	vdp_not g572 (.A(w608), .nZ(w854) );
	vdp_comp_str g573 (.A(w570), .Z(w636), .nZ(w637) );
	vdp_not g574 (.A(w586), .nZ(w652) );
	vdp_not g575 (.A(w632), .nZ(w1556) );
	vdp_comp_str g576 (.A(w468), .Z(w1477), .nZ(w633) );
	vdp_not g577 (.A(w628), .nZ(w627) );
	vdp_comp_str g578 (.A(w459), .Z(w1478), .nZ(w1560) );
	vdp_not g579 (.A(w628), .nZ(w629) );
	vdp_comp_str g580 (.A(w509), .Z(w1479), .nZ(w626) );
	vdp_comp_str g581 (.A(w459), .Z(w630), .nZ(w631) );
	vdp_not g582 (.A(w621), .nZ(w618) );
	vdp_comp_str g583 (.A(w465), .Z(w619), .nZ(w620) );
	vdp_not g584 (.A(w621), .nZ(w853) );
	vdp_comp_str g585 (.A(w465), .Z(w1558), .nZ(w1559) );
	vdp_not g586 (.A(w625), .nZ(w622) );
	vdp_comp_str g587 (.A(w509), .Z(w623), .nZ(w624) );
	vdp_not g588 (.A(w625), .nZ(w1557) );
	vdp_sr_bit g589 (.D(w1445), .Q(w593), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g590 (.D(w641), .Q(w651), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g591 (.D(w584), .Q(w641), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g592 (.D(w675), .Q(w649), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g593 (.D(w577), .Q(w602), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_not g594 (.A(SYSRES), .nZ(w1555) );
	vdp_not g595 (.A(w1527), .nZ(w645) );
	vdp_sr_bit g596 (.D(w599), .Q(w600), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g597 (.D(w590), .C2(HCLK2), .C1(HCLK1), .Q(w596), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_dlatch_inv g598 (.D(w599), .C(HCLK2), .Q(w1527), .nC(nHCLK2) );
	vdp_slatch g599 (.D(w663), .C(w619), .nC(w620), .nQ(w6758) );
	vdp_slatch g600 (.D(w617), .C(w1558), .nC(w1559), .nQ(w6759) );
	vdp_slatch g601 (.D(w663), .C(w623), .nC(w624), .nQ(w6778) );
	vdp_slatch g602 (.D(w617), .C(w1479), .nC(w626), .nQ(w6776) );
	vdp_slatch g603 (.D(w663), .C(w1478), .nC(w1560), .nQ(w6792) );
	vdp_slatch g604 (.D(w617), .C(w630), .nC(w631), .nQ(w6794) );
	vdp_slatch g605 (.D(w663), .C(w1477), .nC(w633), .nQ(w6812) );
	vdp_slatch g606 (.D(w617), .C(w1476), .nC(w1475), .nQ(w6810) );
	vdp_slatch g607 (.D(VRAMA[9]), .C(w1474), .nC(w635), .nQ(w6826) );
	vdp_slatch g608 (.D(VRAMA[7]), .C(w636), .nC(w637), .nQ(w6827) );
	vdp_notif0 g609 (.nZ(VRAMA[7]), .nE(w854), .A(w6827) );
	vdp_notif0 g610 (.nZ(VRAMA[9]), .nE(w1473), .A(w6826) );
	vdp_notif0 g611 (.nZ(VRAMA[7]), .nE(w634), .A(w6810) );
	vdp_notif0 g612 (.nZ(VRAMA[9]), .nE(w1556), .A(w6812) );
	vdp_notif0 g613 (.nZ(VRAMA[7]), .nE(w629), .A(w6794) );
	vdp_notif0 g614 (.nZ(VRAMA[9]), .nE(w622), .A(w6778) );
	vdp_notif0 g615 (.nZ(VRAMA[7]), .nE(w1557), .A(w6776) );
	vdp_notif0 g616 (.nZ(VRAMA[9]), .nE(w627), .A(w6792) );
	vdp_notif0 g617 (.nZ(VRAMA[9]), .nE(w618), .A(w6758) );
	vdp_notif0 g618 (.nZ(VRAMA[7]), .nE(w853), .A(w6759) );
	vdp_bufif0 g619 (.A(w663), .Z(VRAMA[9]), .nE(w652) );
	vdp_bufif0 g620 (.A(w617), .Z(VRAMA[7]), .nE(w652) );
	vdp_bufif0 g621 (.A(w656), .Z(VRAMA[8]), .nE(w1509) );
	vdp_bufif0 g622 (.A(w656), .Z(CA[8]), .nE(w856) );
	vdp_bufif0 g623 (.A(w655), .Z(VRAMA[7]), .nE(w1507) );
	vdp_bufif0 g624 (.A(w655), .Z(CA[7]), .nE(w855) );
	vdp_slatch g625 (.Q(w673), .D(w617), .nQ(w670), .C(w1600), .nC(w1601) );
	vdp_not g626 (.A(w612), .nZ(w668) );
	vdp_not g627 (.A(w617), .nZ(w676) );
	vdp_and3 g628 (.Z(w674), .B(w646), .A(w670), .C(DMA_BUSY) );
	vdp_nand g629 (.A(w666), .Z(w696), .B(w667) );
	vdp_cnt_bit_load g630 (.D(w612), .nL(w1603), .L(w1612), .R(1'b0), .Q(w656), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w638), .CO(w660) );
	vdp_cnt_bit_load g631 (.D(w617), .nL(w1444), .L(w810), .R(1'b0), .Q(w655), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w658), .CO(w640) );
	vdp_cnt_bit_load g632 (.D(w668), .nL(w1602), .L(w818), .R(1'b0), .Q(w666), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w644), .CO(w665) );
	vdp_cnt_bit_load g633 (.D(w676), .nL(w799), .L(w800), .R(1'b0), .Q(w669), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w671), .CO(w648) );
	vdp_slatch g634 (.D(w684), .C(w619), .nC(w620), .nQ(w6757) );
	vdp_slatch g635 (.D(w661), .C(w1558), .nC(w1559), .nQ(w6760) );
	vdp_slatch g636 (.D(w684), .C(w623), .nC(w624), .nQ(w6777) );
	vdp_slatch g637 (.D(w661), .C(w1479), .nC(w626), .nQ(w6775) );
	vdp_slatch g638 (.D(w684), .C(w1478), .nC(w1560), .nQ(w6791) );
	vdp_slatch g639 (.D(w661), .C(w630), .nC(w631), .nQ(w6793) );
	vdp_slatch g640 (.D(w684), .C(w1477), .nC(w633), .nQ(w6811) );
	vdp_slatch g641 (.D(w661), .C(w1476), .nC(w1475), .nQ(w6809) );
	vdp_slatch g642 (.D(VRAMA[10]), .C(w1474), .nC(w635), .nQ(w6825) );
	vdp_slatch g643 (.D(VRAMA[6]), .C(w636), .nC(w637), .nQ(w6828) );
	vdp_notif0 g644 (.nZ(VRAMA[6]), .nE(w854), .A(w6828) );
	vdp_notif0 g645 (.nZ(VRAMA[10]), .nE(w1473), .A(w6825) );
	vdp_notif0 g646 (.nZ(VRAMA[6]), .nE(w634), .A(w6809) );
	vdp_notif0 g647 (.nZ(VRAMA[10]), .nE(w1556), .A(w6811) );
	vdp_notif0 g648 (.nZ(VRAMA[6]), .nE(w629), .A(w6793) );
	vdp_notif0 g649 (.nZ(VRAMA[10]), .nE(w622), .A(w6777) );
	vdp_notif0 g650 (.nZ(VRAMA[6]), .nE(w1557), .A(w6775) );
	vdp_notif0 g651 (.nZ(VRAMA[10]), .nE(w627), .A(w6791) );
	vdp_notif0 g652 (.nZ(VRAMA[10]), .nE(w618), .A(w6757) );
	vdp_notif0 g653 (.nZ(VRAMA[6]), .nE(w853), .A(w6760) );
	vdp_bufif0 g654 (.A(w684), .Z(VRAMA[10]), .nE(w652) );
	vdp_bufif0 g655 (.A(w661), .Z(VRAMA[6]), .nE(w1510) );
	vdp_bufif0 g656 (.A(w654), .Z(VRAMA[9]), .nE(w1509) );
	vdp_bufif0 g657 (.A(w654), .Z(CA[9]), .nE(w856) );
	vdp_bufif0 g658 (.A(w678), .Z(VRAMA[6]), .nE(w1507) );
	vdp_bufif0 g659 (.A(w678), .Z(CA[6]), .nE(w855) );
	vdp_slatch g660 (.Q(w691), .D(w661), .nQ(w646), .C(w1600), .nC(w1601) );
	vdp_not g661 (.A(w685), .nZ(w687) );
	vdp_not g662 (.A(w661), .nZ(w689) );
	vdp_and3 g663 (.Z(w647), .B(DMA_BUSY), .A(w691), .C(w670) );
	vdp_cnt_bit_load g664 (.D(w685), .nL(w1603), .L(w1612), .R(1'b0), .Q(w654), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w660), .CO(w680) );
	vdp_cnt_bit_load g665 (.D(w661), .nL(w1444), .L(w810), .R(1'b0), .Q(w678), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w679), .CO(w658) );
	vdp_cnt_bit_load g666 (.D(w687), .nL(w1602), .L(w818), .R(1'b0), .Q(w667), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w665), .CO(w686) );
	vdp_cnt_bit_load g667 (.D(w689), .nL(w799), .L(w800), .R(1'b0), .Q(w688), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w692), .CO(w671) );
	vdp_nand3 g668 (.Z(w695), .B(w688), .A(w694), .C(w669) );
	vdp_slatch g669 (.D(w708), .C(w619), .nC(w620), .nQ(w6756) );
	vdp_slatch g670 (.D(w681), .C(w1558), .nC(w1559), .nQ(w6761) );
	vdp_slatch g671 (.D(w708), .C(w623), .nC(w624), .nQ(w6779) );
	vdp_slatch g672 (.D(w681), .C(w1479), .nC(w626), .nQ(w6774) );
	vdp_slatch g673 (.D(w708), .C(w1478), .nC(w1560), .nQ(w6790) );
	vdp_slatch g674 (.D(w708), .C(w1477), .nC(w633), .nQ(w6813) );
	vdp_slatch g675 (.D(w681), .C(w1476), .nC(w1475), .nQ(w6808) );
	vdp_slatch g676 (.D(VRAMA[11]), .C(w1474), .nC(w635), .nQ(w6824) );
	vdp_slatch g677 (.D(VRAMA[5]), .C(w636), .nC(w637), .nQ(w6829) );
	vdp_notif0 g678 (.nZ(VRAMA[5]), .nE(w854), .A(w6829) );
	vdp_notif0 g679 (.nZ(VRAMA[11]), .nE(w1473), .A(w6824) );
	vdp_notif0 g680 (.nZ(VRAMA[5]), .nE(w634), .A(w6808) );
	vdp_notif0 g681 (.nZ(VRAMA[11]), .nE(w1556), .A(w6813) );
	vdp_notif0 g682 (.nZ(VRAMA[5]), .nE(w629), .A(w6795) );
	vdp_notif0 g683 (.nZ(VRAMA[11]), .nE(w622), .A(w6779) );
	vdp_notif0 g684 (.nZ(VRAMA[5]), .nE(w1557), .A(w6774) );
	vdp_notif0 g685 (.nZ(VRAMA[11]), .nE(w627), .A(w6790) );
	vdp_notif0 g686 (.nZ(VRAMA[11]), .nE(w618), .A(w6756) );
	vdp_notif0 g687 (.nZ(VRAMA[5]), .nE(w853), .A(w6761) );
	vdp_bufif0 g688 (.A(w708), .Z(VRAMA[11]), .nE(w652) );
	vdp_bufif0 g689 (.A(w681), .Z(VRAMA[5]), .nE(w1510) );
	vdp_bufif0 g690 (.A(w677), .Z(VRAMA[10]), .nE(w1509) );
	vdp_bufif0 g691 (.A(w677), .Z(CA[10]), .nE(w856) );
	vdp_bufif0 g692 (.A(w710), .Z(VRAMA[5]), .nE(w1507) );
	vdp_bufif0 g693 (.A(w710), .Z(CA[5]), .nE(w855) );
	vdp_slatch g694 (.Q(CA[18]), .D(w698), .C(w1600), .nC(w1601) );
	vdp_not g695 (.A(w698), .nZ(w703) );
	vdp_not g696 (.A(w681), .nZ(w702) );
	vdp_and3 g697 (.Z(w591), .B(DMA_BUSY), .A(w691), .C(w673) );
	vdp_cnt_bit_load g698 (.D(w698), .nL(w1603), .L(w1612), .R(1'b0), .Q(w677), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w680), .CO(w713) );
	vdp_cnt_bit_load g699 (.D(w681), .nL(w1444), .L(w810), .R(1'b0), .Q(w710), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w709), .CO(w679) );
	vdp_cnt_bit_load g700 (.D(w703), .nL(w1602), .L(w818), .R(1'b0), .Q(w693), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w686), .CO(w704) );
	vdp_cnt_bit_load g701 (.D(w702), .nL(w799), .L(w800), .R(1'b0), .Q(w694), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w699), .CO(w692) );
	vdp_nand3 g702 (.Z(w707), .B(w705), .A(w706), .C(w693) );
	vdp_slatch g703 (.D(w722), .C(w619), .nC(w620), .nQ(w6755) );
	vdp_slatch g704 (.D(w725), .C(w1558), .nC(w1559), .nQ(w6762) );
	vdp_slatch g705 (.D(w722), .C(w623), .nC(w624), .nQ(w6780) );
	vdp_slatch g706 (.D(w725), .C(w1479), .nC(w626), .nQ(w6773) );
	vdp_slatch g707 (.D(w722), .C(w1478), .nC(w1560), .nQ(w6789) );
	vdp_slatch g708 (.D(w722), .C(w1477), .nC(w633), .nQ(w6814) );
	vdp_slatch g709 (.D(w725), .C(w1476), .nC(w1475), .nQ(w6807) );
	vdp_slatch g710 (.D(VRAMA[12]), .C(w1474), .nC(w635), .nQ(w6823) );
	vdp_slatch g711 (.D(VRAMA[4]), .C(w636), .nC(w637), .nQ(w6830) );
	vdp_notif0 g712 (.nZ(VRAMA[4]), .nE(w854), .A(w6830) );
	vdp_notif0 g713 (.nZ(VRAMA[12]), .nE(w1473), .A(w6823) );
	vdp_notif0 g714 (.nZ(VRAMA[4]), .nE(w634), .A(w6807) );
	vdp_notif0 g715 (.nZ(VRAMA[12]), .nE(w1556), .A(w6814) );
	vdp_notif0 g716 (.nZ(VRAMA[4]), .nE(w629), .A(w6796) );
	vdp_notif0 g717 (.nZ(VRAMA[12]), .nE(w622), .A(w6780) );
	vdp_notif0 g718 (.nZ(VRAMA[4]), .nE(w1557), .A(w6773) );
	vdp_notif0 g719 (.nZ(VRAMA[12]), .nE(w627), .A(w6789) );
	vdp_notif0 g720 (.nZ(VRAMA[12]), .nE(w618), .A(w6755) );
	vdp_notif0 g721 (.nZ(VRAMA[4]), .nE(w853), .A(w6762) );
	vdp_bufif0 g722 (.A(w722), .Z(VRAMA[12]), .nE(w652) );
	vdp_bufif0 g723 (.A(w725), .Z(VRAMA[4]), .nE(w1510) );
	vdp_bufif0 g724 (.A(w712), .Z(VRAMA[11]), .nE(w1509) );
	vdp_bufif0 g725 (.A(w712), .Z(CA[11]), .nE(w856) );
	vdp_bufif0 g726 (.A(w723), .Z(VRAMA[4]), .nE(w1507) );
	vdp_bufif0 g727 (.A(w723), .Z(CA[4]), .nE(w855) );
	vdp_slatch g728 (.Q(CA[19]), .D(w719), .C(w1600), .nC(w1601) );
	vdp_not g729 (.A(w719), .nZ(w724) );
	vdp_not g730 (.A(w725), .nZ(w726) );
	vdp_and g731 (.Z(w590), .B(w701), .A(w734) );
	vdp_cnt_bit_load g732 (.D(w719), .nL(w1603), .L(w1612), .R(1'b0), .Q(w712), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w713), .CO(w718) );
	vdp_cnt_bit_load g733 (.D(w725), .nL(w1444), .L(w810), .R(1'b0), .Q(w723), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w728), .CO(w709) );
	vdp_cnt_bit_load g734 (.D(w724), .nL(w1602), .L(w818), .R(1'b0), .Q(w705), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w704), .CO(w729) );
	vdp_cnt_bit_load g735 (.D(w726), .nL(w799), .L(w800), .R(1'b0), .Q(w732), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w733), .CO(w699) );
	vdp_nor3 g736 (.Z(w701), .B(w707), .A(w731), .C(w696) );
	vdp_slatch g737 (.D(w740), .C(w619), .nC(w620), .nQ(w6754) );
	vdp_slatch g738 (.D(w719), .C(w1558), .nC(w1559), .nQ(w6763) );
	vdp_slatch g739 (.D(w740), .C(w623), .nC(w624), .nQ(w6781) );
	vdp_slatch g740 (.D(w719), .C(w1479), .nC(w626), .nQ(w6772) );
	vdp_slatch g741 (.D(w740), .C(w1478), .nC(w1560), .nQ(w6788) );
	vdp_slatch g742 (.D(w719), .C(w630), .nC(w631), .nQ(w6798) );
	vdp_slatch g743 (.D(w740), .C(w1477), .nC(w633), .nQ(w6816) );
	vdp_slatch g744 (.D(w719), .C(w1476), .nC(w1475), .nQ(w6806) );
	vdp_slatch g745 (.D(VRAMA[13]), .C(w1474), .nC(w635), .nQ(w6822) );
	vdp_slatch g746 (.D(VRAMA[3]), .C(w636), .nC(w637), .nQ(w6831) );
	vdp_notif0 g747 (.nZ(VRAMA[3]), .nE(w854), .A(w6831) );
	vdp_notif0 g748 (.nZ(VRAMA[13]), .nE(w1473), .A(w6822) );
	vdp_notif0 g749 (.nZ(VRAMA[3]), .nE(w634), .A(w6806) );
	vdp_notif0 g750 (.nZ(VRAMA[13]), .nE(w1556), .A(w6816) );
	vdp_notif0 g751 (.nZ(VRAMA[3]), .nE(w629), .A(w6798) );
	vdp_notif0 g752 (.nZ(VRAMA[13]), .nE(w622), .A(w6781) );
	vdp_notif0 g753 (.nZ(VRAMA[3]), .nE(w1557), .A(w6772) );
	vdp_notif0 g754 (.nZ(VRAMA[13]), .nE(w627), .A(w6788) );
	vdp_notif0 g755 (.nZ(VRAMA[13]), .nE(w618), .A(w6754) );
	vdp_notif0 g756 (.nZ(VRAMA[3]), .nE(w853), .A(w6763) );
	vdp_bufif0 g757 (.A(w740), .Z(VRAMA[13]), .nE(w652) );
	vdp_bufif0 g758 (.A(w719), .Z(VRAMA[3]), .nE(w1510) );
	vdp_bufif0 g759 (.A(w717), .Z(VRAMA[12]), .nE(w1509) );
	vdp_bufif0 g760 (.A(w717), .Z(CA[12]), .nE(w856) );
	vdp_bufif0 g761 (.A(w748), .Z(VRAMA[3]), .nE(w1507) );
	vdp_bufif0 g762 (.A(w748), .Z(CA[3]), .nE(w855) );
	vdp_slatch g763 (.Q(w755), .D(w725), .C(w1600), .nC(w1601) );
	vdp_not g764 (.A(w725), .nZ(w742) );
	vdp_not g765 (.A(w719), .nZ(w743) );
	vdp_cnt_bit_load g766 (.D(w725), .nL(w1603), .L(w1612), .R(1'b0), .Q(w717), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w718), .CO(w739) );
	vdp_cnt_bit_load g767 (.D(w719), .nL(w1444), .L(w810), .R(1'b0), .Q(w748), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w737), .CO(w728) );
	vdp_cnt_bit_load g768 (.D(w742), .nL(w1602), .L(w818), .R(1'b0), .Q(w706), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w729), .CO(w747) );
	vdp_cnt_bit_load g769 (.D(w743), .nL(w799), .L(w800), .R(1'b0), .Q(w752), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w744), .CO(w733) );
	vdp_nor3 g770 (.Z(w734), .B(w753), .A(w751), .C(w695) );
	vdp_bufif0 g771 (.A(w755), .Z(CA[20]), .nE(w797) );
	vdp_slatch g772 (.D(w759), .C(w619), .nC(w620), .nQ(w6753) );
	vdp_slatch g773 (.D(w698), .C(w1558), .nC(w1559), .nQ(w6764) );
	vdp_slatch g774 (.D(w759), .C(w623), .nC(w624), .nQ(w6782) );
	vdp_slatch g775 (.D(w698), .C(w1479), .nC(w626), .nQ(w6771) );
	vdp_slatch g776 (.D(w759), .C(w1478), .nC(w1560), .nQ(w6787) );
	vdp_slatch g777 (.D(w698), .C(w630), .nC(w631), .nQ(w6797) );
	vdp_slatch g778 (.D(w759), .C(w1477), .nC(w633), .nQ(w6815) );
	vdp_slatch g779 (.D(w698), .C(w1476), .nC(w1475), .nQ(w6805) );
	vdp_slatch g780 (.D(VRAMA[14]), .C(w1474), .nC(w635), .nQ(w6821) );
	vdp_slatch g781 (.D(VRAMA[2]), .nC(w637), .C(w636), .nQ(w6832) );
	vdp_notif0 g782 (.nZ(VRAMA[2]), .nE(w854), .A(w6832) );
	vdp_notif0 g783 (.nZ(VRAMA[14]), .nE(w1473), .A(w6821) );
	vdp_notif0 g784 (.nZ(VRAMA[2]), .nE(w634), .A(w6805) );
	vdp_notif0 g785 (.nZ(VRAMA[14]), .nE(w1556), .A(w6815) );
	vdp_notif0 g786 (.nZ(VRAMA[2]), .nE(w629), .A(w6797) );
	vdp_notif0 g787 (.nZ(VRAMA[14]), .nE(w622), .A(w6782) );
	vdp_notif0 g788 (.nZ(VRAMA[2]), .nE(w1557), .A(w6771) );
	vdp_notif0 g789 (.nZ(VRAMA[14]), .nE(w627), .A(w6787) );
	vdp_notif0 g790 (.nZ(VRAMA[14]), .nE(w618), .A(w6753) );
	vdp_notif0 g791 (.nZ(VRAMA[2]), .nE(w853), .A(w6764) );
	vdp_bufif0 g792 (.A(w759), .Z(VRAMA[14]), .nE(w1508) );
	vdp_bufif0 g793 (.A(w698), .Z(VRAMA[2]), .nE(w1510) );
	vdp_bufif0 g794 (.A(w738), .Z(VRAMA[13]), .nE(w1509) );
	vdp_bufif0 g795 (.A(w738), .Z(CA[13]), .nE(w856) );
	vdp_bufif0 g796 (.A(w760), .Z(VRAMA[2]), .nE(w1507) );
	vdp_bufif0 g797 (.A(w760), .Z(CA[2]), .nE(w855) );
	vdp_slatch g798 (.Q(w767), .D(w681), .C(w1600), .nC(w1601) );
	vdp_not g799 (.A(w681), .nZ(w761) );
	vdp_not g800 (.A(w698), .nZ(w762) );
	vdp_cnt_bit_load g801 (.D(w681), .nL(w1603), .L(w1612), .R(1'b0), .Q(w738), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w739), .CO(w773) );
	vdp_cnt_bit_load g802 (.D(w698), .nL(w1444), .L(w810), .R(1'b0), .Q(w760), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w772), .CO(w737) );
	vdp_cnt_bit_load g803 (.D(w761), .nL(w1602), .L(w818), .R(1'b0), .Q(w771), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w747), .CO(w763) );
	vdp_cnt_bit_load g804 (.D(w762), .nL(w799), .L(w800), .R(1'b0), .Q(w769), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w775), .CO(w744) );
	vdp_nand3 g805 (.Z(w753), .B(w752), .A(w769), .C(w732) );
	vdp_bufif0 g806 (.A(w767), .Z(CA[21]), .nE(w797) );
	vdp_slatch g807 (.D(w780), .C(w619), .nC(w620), .nQ(w6752) );
	vdp_slatch g808 (.D(w685), .C(w1558), .nC(w1559), .nQ(w6765) );
	vdp_slatch g809 (.D(w780), .C(w623), .nC(w624), .nQ(w6784) );
	vdp_slatch g810 (.D(w685), .C(w1479), .nC(w626), .nQ(w6770) );
	vdp_slatch g811 (.D(w780), .C(w1478), .nC(w1560), .nQ(w6786) );
	vdp_slatch g812 (.D(w685), .C(w630), .nC(w631), .nQ(w6800) );
	vdp_slatch g813 (.D(w780), .C(w1477), .nC(w633), .nQ(w6817) );
	vdp_slatch g814 (.D(w685), .C(w1476), .nC(w1475), .nQ(w6804) );
	vdp_slatch g815 (.D(VRAMA[15]), .C(w1474), .nC(w635), .nQ(w6820) );
	vdp_slatch g816 (.D(VRAMA[1]), .C(w636), .nC(w637), .nQ(w6833) );
	vdp_notif0 g817 (.nZ(VRAMA[1]), .nE(w854), .A(w6833) );
	vdp_notif0 g818 (.nZ(VRAMA[15]), .nE(w1473), .A(w6820) );
	vdp_notif0 g819 (.nZ(VRAMA[1]), .nE(w634), .A(w6804) );
	vdp_notif0 g820 (.nZ(VRAMA[15]), .nE(w1556), .A(w6817) );
	vdp_notif0 g821 (.nZ(VRAMA[1]), .nE(w629), .A(w6800) );
	vdp_notif0 g822 (.nZ(VRAMA[15]), .nE(w622), .A(w6784) );
	vdp_notif0 g823 (.nZ(VRAMA[1]), .nE(w1557), .A(w6770) );
	vdp_notif0 g824 (.nZ(VRAMA[15]), .nE(w627), .A(w6786) );
	vdp_notif0 g825 (.nZ(VRAMA[15]), .nE(w618), .A(w6752) );
	vdp_notif0 g826 (.nZ(VRAMA[1]), .nE(w853), .A(w6765) );
	vdp_bufif0 g827 (.A(w780), .Z(VRAMA[15]), .nE(w1508) );
	vdp_bufif0 g828 (.A(w685), .Z(VRAMA[1]), .nE(w1510) );
	vdp_bufif0 g829 (.A(w756), .Z(VRAMA[14]), .nE(w1509) );
	vdp_bufif0 g830 (.A(w756), .Z(CA[14]), .nE(w856) );
	vdp_bufif0 g831 (.A(w782), .Z(VRAMA[1]), .nE(w1507) );
	vdp_bufif0 g832 (.A(w782), .Z(CA[1]), .nE(w855) );
	vdp_slatch g833 (.Q(w1511), .D(w685), .C(w1600), .nC(w1601) );
	vdp_not g834 (.A(w661), .nZ(w785) );
	vdp_not g835 (.A(w685), .nZ(w788) );
	vdp_cnt_bit_load g836 (.D(w661), .nL(w1603), .L(w1612), .R(1'b0), .Q(w756), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w773), .CO(w789) );
	vdp_cnt_bit_load g837 (.D(w685), .nL(w1444), .L(w810), .R(1'b0), .Q(w782), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w790), .CO(w772) );
	vdp_cnt_bit_load g838 (.D(w785), .nL(w1602), .L(w818), .R(1'b0), .Q(w770), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w763), .CO(w783) );
	vdp_cnt_bit_load g839 (.D(w788), .nL(w799), .L(w800), .R(1'b0), .Q(w787), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w786), .CO(w775) );
	vdp_nand3 g840 (.Z(w731), .B(w770), .A(w771), .C(w784) );
	vdp_bufif0 g841 (.A(w1511), .Z(CA[17]), .nE(w797) );
	vdp_slatch g842 (.nQ(w781), .D(w794), .C(w619), .nC(w620) );
	vdp_slatch g843 (.D(w612), .C(w1558), .nC(w1559), .nQ(w6766) );
	vdp_slatch g844 (.D(w794), .C(w623), .nC(w624), .nQ(w6783) );
	vdp_slatch g845 (.D(w612), .C(w1479), .nC(w626), .nQ(w6769) );
	vdp_slatch g846 (.D(w794), .C(w1478), .nC(w1560), .nQ(w6785) );
	vdp_slatch g847 (.D(w612), .C(w630), .nC(w631), .nQ(w6799) );
	vdp_slatch g848 (.D(w794), .C(w1477), .nC(w633), .nQ(w6818) );
	vdp_slatch g849 (.D(w612), .C(w1476), .nC(w1475), .nQ(w6803) );
	vdp_slatch g850 (.D(VRAMA[16]), .C(w1474), .nC(w635), .nQ(w6819) );
	vdp_slatch g851 (.Q(w6834), .D(VRAMA[0]), .C(w636), .nC(w637) );
	vdp_notif0 g852 (.nZ(VRAMA[0]), .nE(w854), .A(w6834) );
	vdp_notif0 g853 (.nZ(VRAMA[16]), .nE(w1473), .A(w6819) );
	vdp_notif0 g854 (.nZ(VRAMA[0]), .nE(w634), .A(w6803) );
	vdp_notif0 g855 (.nZ(VRAMA[16]), .nE(w1556), .A(w6818) );
	vdp_notif0 g856 (.nZ(VRAMA[0]), .nE(w629), .A(w6799) );
	vdp_notif0 g857 (.nZ(VRAMA[16]), .nE(w622), .A(w6783) );
	vdp_notif0 g858 (.nZ(VRAMA[0]), .nE(w1557), .A(w6769) );
	vdp_notif0 g859 (.nZ(VRAMA[16]), .nE(w627), .A(w6785) );
	vdp_notif0 g860 (.A(w781), .nZ(VRAMA[16]), .nE(w618) );
	vdp_notif0 g861 (.nZ(VRAMA[0]), .nE(w853), .A(w6766) );
	vdp_bufif0 g862 (.A(w794), .Z(VRAMA[16]), .nE(w1508) );
	vdp_bufif0 g863 (.A(w612), .Z(VRAMA[0]), .nE(w1510) );
	vdp_bufif0 g864 (.A(w776), .Z(VRAMA[15]), .nE(w1509) );
	vdp_bufif0 g865 (.A(w776), .Z(CA[15]), .nE(w856) );
	vdp_bufif0 g866 (.A(w804), .Z(VRAMA[0]), .nE(w1507) );
	vdp_bufif0 g867 (.A(w804), .Z(CA[0]), .nE(w855) );
	vdp_slatch g868 (.Q(w795), .D(w612), .C(w1600), .nC(w1601) );
	vdp_not g869 (.A(w617), .nZ(w1604) );
	vdp_not g870 (.A(w612), .nZ(w1481) );
	vdp_cnt_bit_load g871 (.D(w617), .nL(w1603), .L(w1612), .R(1'b0), .Q(w776), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w789) );
	vdp_cnt_bit_load g872 (.D(w612), .nL(w1444), .L(w810), .R(1'b0), .Q(w804), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w802), .CO(w790) );
	vdp_cnt_bit_load g873 (.D(w1604), .nL(w1602), .L(w818), .R(1'b0), .Q(w784), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w783) );
	vdp_cnt_bit_load g874 (.D(w1481), .nL(w799), .L(w800), .R(1'b0), .Q(w1480), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w802), .CO(w786) );
	vdp_nand3 g875 (.Z(w751), .B(w787), .A(w598), .C(w1439) );
	vdp_bufif0 g876 (.A(w795), .Z(CA[16]), .nE(w797) );
	vdp_slatch g877 (.D(VRAMA[8]), .C(w636), .nC(w637), .nQ(w6835) );
	vdp_slatch g878 (.D(w597), .C(w1476), .nC(w1475), .nQ(w6802) );
	vdp_slatch g879 (.D(w597), .C(w630), .nC(w631), .nQ(w6801) );
	vdp_slatch g880 (.D(w597), .C(w1479), .nC(w626), .nQ(w6768) );
	vdp_slatch g881 (.D(w597), .C(w1558), .nC(w1559), .nQ(w6767) );
	vdp_notif0 g882 (.nZ(VRAMA[8]), .nE(w853), .A(w6767) );
	vdp_notif0 g883 (.nZ(VRAMA[8]), .nE(w1557), .A(w6768) );
	vdp_notif0 g884 (.nZ(VRAMA[8]), .nE(w629), .A(w6801) );
	vdp_notif0 g885 (.nZ(VRAMA[8]), .nE(w634), .A(w6802) );
	vdp_notif0 g886 (.nZ(VRAMA[8]), .nE(w854), .A(w6835) );
	vdp_bufif0 g887 (.A(w795), .Z(VRAMA[16]), .nE(w1509) );
	vdp_not g888 (.A(w1472), .nZ(w1508) );
	vdp_not g889 (.A(w586), .nZ(w1510) );
	vdp_not g890 (.A(w33), .nZ(w1509) );
	vdp_not g891 (.A(w594), .nZ(w856) );
	vdp_not g892 (.A(w33), .nZ(w1507) );
	vdp_not g893 (.A(w594), .nZ(w855) );
	vdp_not g894 (.A(w594), .nZ(w797) );
	vdp_not g895 (.A(w1480), .nZ(w1439) );
	vdp_not g896 (.A(w798), .nZ(w1443) );
	vdp_not g897 (.A(M5), .nZ(w815) );
	vdp_and4 g898 (.Z(w811), .B(w684), .A(w820), .D(w597), .C(w821) );
	vdp_and4 g899 (.Z(w812), .B(w684), .A(w820), .D(w823), .C(w663) );
	vdp_and4 g900 (.B(w824), .A(w805), .D(w823), .C(w821), .Z(w814) );
	vdp_and4 g901 (.B(w824), .A(w805), .D(w597), .C(w821), .Z(w813) );
	vdp_and4 g902 (.Z(w808), .B(w821), .A(w597), .D(w825), .C(w684) );
	vdp_and4 g903 (.Z(w806), .B(w663), .A(w823), .D(w805), .C(w824) );
	vdp_and4 g904 (.Z(w807), .B(w663), .A(w597), .D(w825), .C(w684) );
	vdp_and4 g905 (.B(w828), .A(M5), .D(w708), .C(w829), .Z(w820) );
	vdp_comp_str g906 (.A(w831), .Z(w1600), .nZ(w1601) );
	vdp_comp_we g907 (.A(w1485), .Z(w1612), .nZ(w1603) );
	vdp_comp_we g908 (.A(w809), .Z(w810), .nZ(w1444) );
	vdp_comp_we g909 (.A(w832), .Z(w818), .nZ(w1602) );
	vdp_comp_we g910 (.A(w833), .Z(w800), .nZ(w799) );
	vdp_and g911 (.Z(w607), .B(w598), .A(w798) );
	vdp_and g912 (.Z(w802), .B(w598), .A(w1443) );
	vdp_or g913 (.Z(w831), .B(w807), .A(SYSRES) );
	vdp_or g914 (.Z(w809), .B(w808), .A(SYSRES) );
	vdp_or g915 (.Z(w1472), .B(w815), .A(w586) );
	vdp_or g916 (.B(w813), .A(SYSRES), .Z(w87) );
	vdp_or g917 (.B(w814), .A(SYSRES), .Z(w86) );
	vdp_or g918 (.Z(w85), .B(w812), .A(SYSRES) );
	vdp_or g919 (.Z(w68), .B(w811), .A(SYSRES) );
	vdp_or g920 (.B(w1482), .A(SYSRES), .Z(w72) );
	vdp_and4 g921 (.B(w684), .A(w822), .D(w597), .C(w663), .Z(w840) );
	vdp_or g922 (.B(w840), .A(SYSRES), .Z(w73) );
	vdp_and4 g923 (.B(w824), .A(w825), .D(w823), .C(w663), .Z(w839) );
	vdp_or g924 (.B(w839), .A(SYSRES), .Z(w75) );
	vdp_and4 g925 (.B(w824), .A(w825), .D(w597), .C(w821), .Z(w838) );
	vdp_or g926 (.B(w838), .A(SYSRES), .Z(w74) );
	vdp_and4 g927 (.B(w824), .A(w825), .D(w823), .C(w821), .Z(w1483) );
	vdp_or g928 (.B(w1483), .A(SYSRES), .Z(w69) );
	vdp_and4 g929 (.B(w684), .A(w822), .D(w823), .C(w663), .Z(w837) );
	vdp_or g930 (.B(w837), .A(SYSRES), .Z(w143) );
	vdp_and4 g931 (.B(w684), .A(w822), .D(w597), .C(w821), .Z(w836) );
	vdp_or g932 (.B(w836), .A(SYSRES), .Z(w142) );
	vdp_or g933 (.B(w841), .A(SYSRES), .Z(w71) );
	vdp_and4 g934 (.B(w684), .A(w822), .D(w823), .C(w821), .Z(w1482) );
	vdp_or g935 (.B(w842), .A(SYSRES), .Z(w70) );
	vdp_and4 g936 (.B(w824), .A(w822), .D(w597), .C(w663), .Z(w841) );
	vdp_and4 g937 (.B(w824), .A(w822), .D(w823), .C(w663), .Z(w842) );
	vdp_and4 g938 (.B(w821), .A(w597), .D(w822), .C(w824), .Z(w844) );
	vdp_or g939 (.B(w844), .A(SYSRES), .Z(w1140) );
	vdp_and4 g940 (.B(w821), .A(w823), .D(w822), .C(w824), .Z(w1484) );
	vdp_or g941 (.B(w1484), .A(SYSRES), .Z(w1179) );
	vdp_and4 g942 (.B(w821), .A(w823), .D(w820), .C(w684), .Z(w843) );
	vdp_or g943 (.B(w843), .A(SYSRES), .Z(w1141) );
	vdp_and4 g944 (.B(w663), .A(w823), .D(w825), .C(w684), .Z(w845) );
	vdp_or g945 (.B(w845), .A(SYSRES), .Z(w1485) );
	vdp_and4 g946 (.B(w663), .A(w597), .D(w820), .C(w824), .Z(w1486) );
	vdp_or g947 (.B(w1486), .A(SYSRES), .Z(CA[14]) );
	vdp_and4 g948 (.B(w821), .A(w823), .D(w825), .C(w684), .Z(w846) );
	vdp_or g949 (.B(w846), .A(SYSRES), .Z(w832) );
	vdp_and4 g950 (.B(w663), .A(w597), .D(w825), .C(w824), .Z(w847) );
	vdp_or g951 (.B(w847), .A(SYSRES), .Z(w833) );
	vdp_and4 g952 (.B(w663), .A(w834), .D(w820), .C(w684), .Z(w848) );
	vdp_or g953 (.B(w848), .A(SYSRES), .Z(w849) );
	vdp_and4 g954 (.B(w830), .A(w828), .D(M5), .C(w722), .Z(w825) );
	vdp_and3 g955 (.B(w829), .A(w828), .C(w708), .Z(w805) );
	vdp_and3 g956 (.B(w830), .A(w828), .C(w829), .Z(w822) );
	vdp_or g957 (.Z(w850), .B(w851), .A(w6737) );
	vdp_and g958 (.B(w827), .A(HCLK1), .Z(w828) );
	vdp_dlatch_inv g959 (.D(w826), .C(DCLK2), .nQ(w851), .nC(nDCLK2) );
	vdp_dlatch_inv g960 (.D(w6736), .C(HCLK2), .nQ(w827), .nC(nHCLK2) );
	vdp_not g961 (.A(w722), .nZ(w829) );
	vdp_not g962 (.A(w708), .nZ(w830) );
	vdp_not g963 (.A(w663), .nZ(w821) );
	vdp_not g964 (.A(w684), .nZ(w824) );
	vdp_not g965 (.A(w597), .nZ(w823) );
	vdp_slatch g966 (.D(w681), .C(w630), .nC(w631), .nQ(w6795) );
	vdp_slatch g967 (.D(w725), .C(w630), .nC(w631), .nQ(w6796) );
	vdp_sr_bit g968 (.D(w851), .C2(DCLK2), .C1(DCLK1), .Q(w6737), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_dlatch_inv g969 (.D(w850), .C(DCLK1), .nQ(w6736), .nC(nDCLK1) );
	vdp_comp_str g970 (.A(w888), .Z(w858), .nZ(w866) );
	vdp_fa g971 (.SUM(w885), .A(w661), .B(w1577), .CO(w887), .CI(w883) );
	vdp_fa g972 (.SUM(w881), .A(w681), .B(w882), .CO(w883), .CI(w880) );
	vdp_fa g973 (.SUM(w878), .A(w725), .B(w879), .CO(w880), .CI(w875) );
	vdp_fa g974 (.SUM(w874), .A(w719), .B(w877), .CO(w875), .CI(w872) );
	vdp_fa g975 (.SUM(w870), .A(w698), .B(w871), .CO(w872), .CI(w869) );
	vdp_fa g976 (.SUM(w6740), .A(w685), .B(w868), .CO(w869), .CI(w865) );
	vdp_fa g977 (.SUM(w6741), .A(w612), .B(w862), .CO(w865), .CI(w860) );
	vdp_fa g978 (.SUM(w1487), .A(w617), .B(w1576), .CO(w889), .CI(w887) );
	vdp_slatch g979 (.Q(w886), .D(w160), .C(w858), .nC(w866) );
	vdp_aon22 g980 (.Z(w1587), .A1(w886), .A2(w857), .B1(w863), .B2(w1487) );
	vdp_slatch g981 (.Q(w884), .D(DB[6]), .C(w858), .nC(w866) );
	vdp_aon22 g982 (.Z(w1588), .A1(w884), .A2(w857), .B1(w863), .B2(w885) );
	vdp_slatch g983 (.Q(w1530), .D(DB[5]), .C(w858), .nC(w866) );
	vdp_aon22 g984 (.Z(w1589), .A1(w1530), .A2(w857), .B1(w863), .B2(w881) );
	vdp_slatch g985 (.Q(w876), .D(DB[4]), .C(w858), .nC(w866) );
	vdp_aon22 g986 (.Z(w1590), .A1(w876), .A2(w857), .B1(w863), .B2(w878) );
	vdp_slatch g987 (.Q(w873), .D(w156), .C(w858), .nC(w866) );
	vdp_aon22 g988 (.Z(w1591), .A1(w873), .A2(w857), .B1(w863), .B2(w874) );
	vdp_slatch g989 (.Q(w867), .D(DB[2]), .C(w858), .nC(w866) );
	vdp_aon22 g990 (.Z(w1592), .A1(w867), .A2(w857), .B1(w863), .B2(w870) );
	vdp_slatch g991 (.Q(w864), .D(DB[1]), .C(w858), .nC(w866) );
	vdp_aon22 g992 (.Z(w1593), .A1(w864), .A2(w857), .B1(w863), .B2(w6740) );
	vdp_slatch g993 (.Q(w859), .D(DB[0]), .C(w858), .nC(w866) );
	vdp_aon22 g994 (.Z(w1594), .A1(w859), .A2(w857), .B1(w863), .B2(w6741) );
	vdp_dff g995 (.Q(w612), .R(SYSRES), .C(w891), .D(w1594) );
	vdp_slatch g996 (.Q(w862), .D(w612), .C(w890), .nC(w861) );
	vdp_dff g997 (.Q(w685), .R(SYSRES), .D(w1593), .C(w891) );
	vdp_slatch g998 (.Q(w868), .D(w685), .C(w890), .nC(w861) );
	vdp_dff g999 (.Q(w698), .R(SYSRES), .C(w891), .D(w1592) );
	vdp_slatch g1000 (.Q(w871), .D(w698), .C(w890), .nC(w861) );
	vdp_dff g1001 (.Q(w719), .R(SYSRES), .D(w1591), .C(w891) );
	vdp_slatch g1002 (.Q(w877), .D(w719), .C(w890), .nC(w861) );
	vdp_dff g1003 (.Q(w725), .R(SYSRES), .C(w891), .D(w1590) );
	vdp_slatch g1004 (.Q(w879), .D(w725), .C(w890), .nC(w861) );
	vdp_dff g1005 (.Q(w681), .R(SYSRES), .C(w891), .D(w1589) );
	vdp_slatch g1006 (.Q(w882), .D(w681), .C(w890), .nC(w861) );
	vdp_dff g1007 (.Q(w661), .R(SYSRES), .C(w891), .D(w1588) );
	vdp_slatch g1008 (.Q(w1577), .D(w661), .C(w890), .nC(w861) );
	vdp_dff g1009 (.Q(w617), .R(SYSRES), .D(w1587), .C(w891) );
	vdp_slatch g1010 (.Q(w1576), .D(w617), .C(w890), .nC(w861) );
	vdp_comp_str g1011 (.A(w849), .Z(w890), .nZ(w861) );
	vdp_comp_we g1012 (.A(w894), .Z(w857), .nZ(w863) );
	vdp_dff g1013 (.Q(w794), .R(w898), .C(w891), .D(w1578) );
	vdp_dff g1014 (.Q(w780), .R(w898), .C(w891), .D(w1579) );
	vdp_dff g1015 (.Q(w759), .R(w898), .C(w891), .D(w1580) );
	vdp_dff g1016 (.Q(w740), .R(SYSRES), .C(w891), .D(w1581) );
	vdp_dff g1017 (.Q(w722), .R(SYSRES), .C(w891), .D(w1582) );
	vdp_dff g1018 (.Q(w708), .R(SYSRES), .C(w891), .D(w1583) );
	vdp_dff g1019 (.Q(w684), .R(SYSRES), .C(w891), .D(w1584) );
	vdp_dff g1020 (.Q(w663), .R(SYSRES), .C(w891), .D(w1585) );
	vdp_dff g1021 (.Q(w597), .R(SYSRES), .C(w891), .D(w1586) );
	vdp_not g1022 (.A(w920), .nZ(w891) );
	vdp_or g1023 (.Z(w898), .B(SYSRES), .A(w860) );
	vdp_not g1024 (.A(M5), .nZ(w860) );
	vdp_slatch g1025 (.Q(w917), .D(w932), .C(w931), .nC(w908) );
	vdp_aon22 g1026 (.Z(w1586), .A1(w921), .A2(w929), .B1(w895), .B2(w919) );
	vdp_slatch g1027 (.Q(w921), .D(w245), .C(w931), .nC(w908) );
	vdp_comp_str g1028 (.A(w936), .Z(w931), .nZ(w908) );
	vdp_comp_we g1029 (.A(w894), .Z(w929), .nZ(w895) );
	vdp_ha g1030 (.SUM(w919), .A(w597), .B(w889), .CO(w916) );
	vdp_slatch g1031 (.Q(w915), .D(w253), .C(w931), .nC(w908) );
	vdp_aon22 g1032 (.Z(w1585), .A1(w917), .A2(w929), .B1(w895), .B2(w918) );
	vdp_ha g1033 (.SUM(w918), .A(w663), .B(w916), .CO(w1597) );
	vdp_slatch g1034 (.Q(w913), .D(w289), .C(w931), .nC(w908) );
	vdp_aon22 g1035 (.Z(w1584), .A1(w915), .A2(w929), .B1(w895), .B2(w914) );
	vdp_ha g1036 (.SUM(w914), .A(w684), .B(w1597), .CO(w912) );
	vdp_slatch g1037 (.Q(w910), .D(w262), .C(w931), .nC(w908) );
	vdp_aon22 g1038 (.Z(w1583), .A1(w913), .A2(w929), .B1(w895), .B2(w911) );
	vdp_ha g1039 (.SUM(w911), .A(w708), .B(w912), .CO(w1596) );
	vdp_slatch g1040 (.Q(w907), .D(w299), .C(w931), .nC(w908) );
	vdp_aon22 g1041 (.Z(w1582), .A1(w910), .A2(w929), .B1(w895), .B2(w909) );
	vdp_ha g1042 (.SUM(w909), .A(w722), .B(w1596), .CO(w906) );
	vdp_aon22 g1043 (.Z(w1581), .A1(w907), .A2(w929), .B1(w895), .B2(w904) );
	vdp_ha g1044 (.SUM(w904), .A(w740), .B(w906), .CO(w905) );
	vdp_comp_str g1045 (.A(w930), .Z(w928), .nZ(w897) );
	vdp_aon22 g1046 (.Z(w1580), .A1(w903), .A2(w929), .B1(w895), .B2(w1595) );
	vdp_ha g1047 (.SUM(w1595), .A(w759), .B(w905), .CO(w900) );
	vdp_slatch_r g1048 (.Q(w903), .D(DB[0]), .R(w898), .C(w928), .nC(w897) );
	vdp_slatch_r g1049 (.Q(w902), .D(DB[1]), .R(w898), .C(w928), .nC(w897) );
	vdp_aon22 g1050 (.Z(w1579), .A1(w902), .A2(w929), .B1(w895), .B2(w901) );
	vdp_ha g1051 (.SUM(w901), .A(w780), .B(w900), .CO(w899) );
	vdp_slatch_r g1052 (.Q(w896), .D(DB[2]), .R(w898), .C(w928), .nC(w897) );
	vdp_aon22 g1053 (.Z(w1578), .A1(w896), .A2(w929), .B1(w895), .B2(w1529) );
	vdp_ha g1054 (.SUM(w1529), .A(w794), .B(w899) );
	vdp_and3 g1055 (.C(w925), .A(w923), .B(w924), .Z(w927) );
	vdp_sr_bit g1056 (.D(w1493), .C2(HCLK2), .C1(HCLK1), .nQ(w110), .nC1(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1057 (.D(w945), .Q(w1493), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK2), .nC1(nHCLK1) );
	vdp_not g1058 (.A(w972), .nZ(w947) );
	vdp_not g1059 (.A(w471), .nZ(w1494) );
	vdp_not g1060 (.A(w472), .nZ(w958) );
	vdp_not g1061 (.A(w923), .nZ(w959) );
	vdp_not g1062 (.A(w956), .nZ(w964) );
	vdp_not g1063 (.A(w514), .nZ(w941) );
	vdp_not g1064 (.A(w591), .nZ(w953) );
	vdp_not g1065 (.A(w979), .nZ(w967) );
	vdp_not g1066 (.A(w1495), .nZ(w970) );
	vdp_not g1067 (.A(w968), .nZ(w937) );
	vdp_slatch g1068 (.Q(w498), .D(w934), .C(w935), .nC(w948) );
	vdp_slatch g1069 (.Q(w514), .D(w271), .C(w935), .nC(w948) );
	vdp_comp_str g1070 (.A(w936), .Z(w935), .nZ(w948) );
	vdp_dlatch_inv g1071 (.D(w599), .C(DCLK1), .nQ(w968), .nC(nDCLK1) );
	vdp_dlatch_inv g1072 (.D(w967), .C(DCLK1), .nQ(w966), .nC(nDCLK1) );
	vdp_dlatch_inv g1073 (.D(w981), .C(DCLK2), .nQ(w979), .nC(nDCLK2) );
	vdp_dlatch_inv g1074 (.D(w986), .C(DCLK1), .nQ(w981), .nC(nDCLK1) );
	vdp_slatch g1075 (.Q(w986), .D(w943), .C(DCLK2), .nC(nDCLK2) );
	vdp_slatch g1076 (.Q(w943), .D(w980), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g1077 (.D(w586), .C(HCLK1), .nQ(w942), .nC(nHCLK1) );
	vdp_rs_FF g1078 (.nQ(w939), .R(w988), .S(w987), .Q(w951) );
	vdp_rs_FF g1079 (.Q(w963), .R(w961), .S(w940) );
	vdp_and3 g1080 (.C(w424), .A(w472), .B(w1494), .Z(w946) );
	vdp_and3 g1081 (.C(w958), .A(w471), .B(w424), .Z(w109) );
	vdp_comp_dff g1082 (.D(w962), .C2(HCLK2), .C1(HCLK1), .Q(w955), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_comp_dff g1083 (.D(w952), .C2(HCLK2), .C1(HCLK1), .Q(w954), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g1084 (.C(w32), .A(w951), .B(w593), .Z(w952) );
	vdp_and g1085 (.A(w160), .B(w971), .Z(w933) );
	vdp_and g1086 (.A(w942), .B(w986), .Z(w894) );
	vdp_and g1087 (.A(w954), .B(w953), .Z(w574) );
	vdp_and g1088 (.A(w591), .B(w954), .Z(w595) );
	vdp_and g1089 (.A(w955), .B(w953), .Z(w965) );
	vdp_and g1090 (.A(w591), .B(w955), .Z(w33) );
	vdp_or g1091 (.A(w955), .B(w977), .Z(w961) );
	vdp_or g1092 (.A(w955), .B(w574), .Z(w424) );
	vdp_or g1093 (.A(w591), .B(w453), .Z(w985) );
	vdp_aoi21 g1094 (.A1(w966), .B(SYSRES), .Z(w1495), .A2(w967) );
	vdp_or3 g1095 (.C(w938), .A(w960), .B(w927), .Z(w940) );
	vdp_or3 g1096 (.C(w595), .A(w965), .B(w589), .Z(w586) );
	vdp_or5 g1097 (.C(w949), .A(w937), .B(w586), .Z(w920), .D(w936), .E(w930) );
	vdp_nand3 g1098 (.C(w926), .A(w964), .B(w975), .Z(w826) );
	vdp_2a3oi g1099 (.A1(w925), .B(w982), .Z(w976), .A2(w975), .C(w924) );
	vdp_nand g1100 (.A(w498), .B(w941), .Z(w956) );
	vdp_nor g1101 (.A(w943), .B(w981), .Z(w926) );
	vdp_and4 g1102 (.C(w939), .A(w593), .B(w32), .Z(w962), .D(w963) );
	vdp_nor5 g1103 (.C(w514), .A(w990), .B(w976), .Z(w938), .D(w498), .E(w959) );
	vdp_and g1104 (.A(w591), .B(w990), .Z(w960) );
	vdp_not g1105 (.A(w579), .nZ(w1547) );
	vdp_not g1106 (.A(w1547), .nZ(w1025) );
	vdp_not g1107 (.A(w1006), .nZ(w1041) );
	vdp_not g1108 (.A(w981), .nZ(w1500) );
	vdp_not g1109 (.A(w986), .nZ(w1026) );
	vdp_not g1110 (.A(w1029), .nZ(w936) );
	vdp_not g1111 (.A(w407), .nZ(w957) );
	vdp_not g1112 (.A(w1015), .nZ(w1023) );
	vdp_not g1113 (.A(M5), .nZ(w925) );
	vdp_rs_FF g1114 (.Q(w975), .R(w973), .S(w936) );
	vdp_rs_FF g1115 (.Q(w924), .R(w973), .S(w1048) );
	vdp_rs_FF g1116 (.Q(w982), .R(w973), .S(w971) );
	vdp_rs_FF g1117 (.nQ(w984), .R(w983), .S(w950) );
	vdp_rs_FF g1118 (.Q(w1045), .R(w970), .S(w978) );
	vdp_rs_FF g1119 (.Q(w569), .R(w970), .S(w1039) );
	vdp_rs_FF g1120 (.Q(w568), .R(w970), .S(w996) );
	vdp_or g1121 (.A(w996), .B(w1039), .Z(w1047) );
	vdp_and g1122 (.A(w1045), .B(w923), .Z(w576) );
	vdp_and g1123 (.A(w1044), .B(w1045), .Z(w579) );
	vdp_and g1124 (.A(w1026), .B(w1500), .Z(w923) );
	vdp_and g1125 (.A(w1026), .B(w979), .Z(w1044) );
	vdp_and g1126 (.A(w981), .B(w979), .Z(w1013) );
	vdp_and g1127 (.A(w955), .B(w985), .Z(w987) );
	vdp_and g1128 (.A(w1009), .B(w997), .Z(w415) );
	vdp_and g1129 (.A(w957), .B(w888), .Z(w1054) );
	vdp_and g1130 (.A(w1032), .B(w1031), .Z(w978) );
	vdp_or g1131 (.A(w954), .B(w977), .Z(w988) );
	vdp_or g1132 (.A(w428), .B(w1028), .Z(w969) );
	vdp_or g1133 (.A(SYSRES), .B(w923), .Z(w983) );
	vdp_or g1134 (.A(SYSRES), .B(w986), .Z(w1051) );
	vdp_or g1135 (.A(w981), .B(w980), .Z(w1046) );
	vdp_or g1136 (.A(w1009), .B(w1032), .Z(w1052) );
	vdp_or g1137 (.A(w974), .B(SYSRES), .Z(w1019) );
	vdp_or g1138 (.A(SYSRES), .B(w1014), .Z(w1056) );
	vdp_or g1139 (.A(SYSRES), .B(w1013), .Z(w973) );
	vdp_and g1140 (.A(w972), .B(w946), .Z(w131) );
	vdp_and g1141 (.A(w946), .B(w947), .Z(w108) );
	vdp_and g1142 (.A(w923), .B(w1021), .Z(w1055) );
	vdp_nand g1143 (.A(w415), .B(w984), .Z(w1037) );
	vdp_nor g1144 (.A(w675), .B(w1025), .Z(w1038) );
	vdp_or5 g1145 (.C(w936), .A(w1024), .B(w1036), .Z(w1035), .D(w888), .E(w1040) );
	vdp_or3 g1146 (.C(w1027), .A(w1009), .B(w410), .Z(w1028) );
	vdp_nor g1147 (.A(w109), .B(w946), .Z(w945) );
	vdp_and3 g1148 (.C(w1057), .A(w1053), .B(w1011), .Z(w1030) );
	vdp_or4 g1149 (.C(w978), .A(w971), .B(w1008), .Z(w974), .D(w415) );
	vdp_and4 g1150 (.C(w1053), .A(w1032), .B(w1016), .Z(w888), .D(w1033) );
	vdp_aoi21 g1151 (.A1(w923), .B(SYSRES), .Z(w1015), .A2(w1022) );
	vdp_aoi21 g1152 (.A1(w888), .B(w1030), .Z(w1029), .A2(w407) );
	vdp_or5 g1153 (.C(w415), .A(w1008), .B(w971), .Z(w1014), .D(w978), .E(w936) );
	vdp_and5 g1154 (.C(w1020), .A(M5), .B(w1053), .Z(w971), .D(w1033), .E(w1032) );
	vdp_not g1155 (.A(CA[7]), .nZ(w1002) );
	vdp_not g1156 (.A(w1032), .nZ(w1010) );
	vdp_not g1157 (.A(w1010), .nZ(w994) );
	vdp_not g1158 (.A(w1009), .nZ(w993) );
	vdp_not g1159 (.A(w993), .nZ(w992) );
	vdp_slatch g1160 (.Q(w1034), .D(w995), .nC(w992), .C(w993) );
	vdp_slatch g1161 (.Q(w1053), .D(w995), .nC(w994), .C(w1010), .nQ(w1031) );
	vdp_rs_FF g1162 (.Q(w1017), .R(w1013), .S(w1019) );
	vdp_rs_FF g1163 (.Q(w1021), .R(w1056), .S(w1054), .nQ(w1022) );
	vdp_rs_FF g1164 (.Q(w1057), .R(w1023), .S(w1055), .nQ(w1033) );
	vdp_rs_FF g1165 (.Q(w1020), .R(w1018), .S(w1491), .nQ(w1016) );
	vdp_slatch_r g1166 (.Q(w990), .D(DB[6]), .C(w1012), .nC(w991), .R(w898) );
	vdp_slatch_r g1167 (.Q(w472), .D(DB[5]), .R(w898), .C(w1012), .nC(w991) );
	vdp_slatch_r g1168 (.Q(w471), .D(DB[4]), .R(w898), .C(w1012), .nC(w991) );
	vdp_comp_str g1169 (.A(w971), .Z(w1012), .nZ(w991) );
	vdp_not g1170 (.A(w1492), .nZ(w1018) );
	vdp_aoi21 g1171 (.A1(w923), .B(SYSRES), .Z(w1492), .A2(w1017) );
	vdp_and4 g1172 (.C(w956), .A(M5), .B(w975), .Z(w1491), .D(w923) );
	vdp_and g1173 (.A(w1009), .B(w1034), .Z(w1048) );
	vdp_rs_FF g1174 (.nQ(w1050), .R(w1049), .S(w1048) );
	vdp_rs_FF g1175 (.Q(w980), .R(w1051), .S(w1052) );
	vdp_not g1176 (.A(w995), .nZ(w1598) );
	vdp_not g1177 (.A(CA[2]), .nZ(w1081) );
	vdp_not g1178 (.A(CA[3]), .nZ(w1082) );
	vdp_aon22 g1179 (.Z(w995), .A1(CA[0]), .A2(w1109), .B1(w407), .B2(w1084) );
	vdp_and4 g1180 (.C(w1000), .A(w1002), .B(w1001), .Z(w1043), .D(w999) );
	vdp_and4 g1181 (.C(w1005), .A(w1004), .B(CA[7]), .Z(w1011), .D(w999) );
	vdp_and4 g1182 (.C(CA[3]), .A(w1041), .B(w1042), .Z(w1027), .D(CA[9]) );
	vdp_and4 g1183 (.C(CA[2]), .A(w1041), .B(w1042), .Z(w406), .D(w1082) );
	vdp_and4 g1184 (.C(w1006), .A(w1081), .B(CA[3]), .Z(w1003), .D(w1042) );
	vdp_or g1185 (.A(w1043), .B(w406), .Z(w410) );
	vdp_and g1186 (.A(w978), .B(w1038), .Z(w1036) );
	vdp_and g1187 (.A(w1028), .B(w1037), .Z(w1040) );
	vdp_and g1188 (.A(w407), .B(w1035), .Z(w1072) );
	vdp_or g1189 (.A(SYSRES), .B(w950), .Z(w1049) );
	vdp_or g1190 (.A(w1011), .B(w998), .Z(w1032) );
	vdp_or g1191 (.A(SYSRES), .B(w596), .Z(w977) );
	vdp_and3 g1192 (.C(w1080), .A(w971), .B(w1050), .Z(w1024) );
	vdp_and3 g1193 (.C(w1083), .A(w1046), .B(w1215), .Z(w1042) );
	vdp_and5 g1194 (.C(CA[2]), .A(w1006), .B(CA[3]), .Z(w1077), .D(w1598), .E(w1042) );
	vdp_and5 g1195 (.C(CA[2]), .A(w1006), .B(w995), .Z(w1076), .D(CA[3]), .E(w1042) );
	vdp_and5 g1196 (.C(w1081), .A(w1047), .B(w1041), .Z(w1007), .D(w1082), .E(w1042) );
	vdp_and5 g1197 (.C(w1082), .A(w1081), .B(w1047), .Z(w998), .D(w1006), .E(w1042) );
	vdp_nor5 g1198 (.C(w1073), .A(w1076), .B(w1077), .Z(w1059), .D(w1003), .E(w1072) );
	vdp_aon22 g1199 (.Z(w1070), .A1(w4), .A2(w1079), .B1(w27), .B2(w407) );
	vdp_aon22 g1200 (.Z(w176), .A1(w1062), .A2(VPOS[8]), .B1(w1067), .B2(VPOS[0]) );
	vdp_not g1201 (.A(w1062), .nZ(w1067) );
	vdp_not g1202 (.A(w407), .nZ(w1063) );
	vdp_not g1203 (.A(w407), .nZ(w1079) );
	vdp_not g1204 (.A(w1544), .nZ(w114) );
	vdp_not g1205 (.A(w1001), .nZ(w1004) );
	vdp_not g1206 (.A(w1489), .nZ(w1068) );
	vdp_not g1207 (.A(w995), .nZ(w997) );
	vdp_aoi21 g1208 (.A1(w996), .B(w1490), .Z(w1489), .A2(w1003) );
	vdp_and4 g1209 (.C(w1000), .A(w1004), .B(CA[7]), .Z(w1488), .D(w999) );
	vdp_and4 g1210 (.C(w1005), .A(w1002), .B(w1001), .Z(w1490), .D(w999) );
	vdp_slatch g1211 (.Q(w116), .D(w1000), .C(w1599), .nC(w1545) );
	vdp_comp_we g1212 (.A(w1061), .Z(w1599), .nZ(w1545) );
	vdp_and g1213 (.A(w47), .B(w1074), .Z(w1546) );
	vdp_and g1214 (.A(w995), .B(w1009), .Z(w1008) );
	vdp_or g1215 (.A(w1007), .B(w1488), .Z(w1009) );
	vdp_or g1216 (.A(w1073), .B(w1546), .Z(w1075) );
	vdp_or g1217 (.Z(w1069), .A(w7), .B(SYSRES) );
	vdp_and g1218 (.Z(w112), .A(w58), .B(w1070) );
	vdp_rs_FF g1219 (.Q(w1065), .R(w1069), .S(w112) );
	vdp_aoi221 g1220 (.Z(w1544), .A1(w113), .A2(1'b0), .B1(w1071), .B2(w1075), .C(w115) );
	vdp_aoi22 g1221 (.Z(w1060), .A1(w1066), .A2(w1063), .B1(w407), .B2(w1065) );
	vdp_comp_str g1222 (.Z(w1097), .A(w58), .nZ(w1098) );
	vdp_comp_str g1223 (.Z(w1123), .A(CA[14]), .nZ(w1124) );
	vdp_comp_str g1224 (.Z(w1133), .A(w1141), .nZ(w1134) );
	vdp_comp_str g1225 (.Z(w1130), .A(w1140), .nZ(w1129) );
	vdp_not g1226 (.A(w1139), .nZ(w1142) );
	vdp_not g1227 (.A(w1131), .nZ(w1144) );
	vdp_not g1228 (.A(w1128), .nZ(w1143) );
	vdp_not g1229 (.A(w1143), .nZ(w1108) );
	vdp_not g1230 (.A(w407), .nZ(w1109) );
	vdp_not g1231 (.A(w1144), .nZ(w1127) );
	vdp_not g1232 (.A(w1146), .nZ(w1126) );
	vdp_not g1233 (.A(w1145), .nZ(w1125) );
	vdp_aon222 g1234 (.C2(w1125), .B2(w1126), .A2(w1127), .C1(w1106), .B1(CA[15]), .A1(CA[7]), .Z(w1118) );
	vdp_aon222 g1235 (.C2(w1125), .B2(w1126), .A2(w1127), .C1(w1105), .B1(CA[13]), .A1(w1001), .Z(w1117) );
	vdp_aon222 g1236 (.C2(w1125), .B2(w1126), .A2(w1127), .C1(w1104), .B1(CA[12]), .A1(CA[5]), .Z(w1116) );
	vdp_aon222 g1237 (.C2(w1125), .B2(w1126), .A2(w1127), .C1(w1103), .B1(CA[11]), .A1(CA[4]), .Z(w1115) );
	vdp_aon222 g1238 (.C2(w1125), .B2(w1126), .A2(w1127), .C1(w1107), .B1(CA[10]), .A1(CA[3]), .Z(w1114) );
	vdp_aon222 g1239 (.C2(w1125), .B2(w1126), .A2(w1127), .C1(w1528), .B1(CA[9]), .A1(CA[2]), .Z(w1113) );
	vdp_aon222 g1240 (.C2(w1125), .B2(w1126), .A2(w1127), .C1(w1110), .B1(CA[8]), .A1(w1084), .Z(w1112) );
	vdp_aon222 g1241 (.C2(w1125), .B2(w1126), .A2(w1127), .C1(w1100), .B1(CA[14]), .A1(CA[0]), .Z(w1111) );
	vdp_aon222 g1242 (.C2(w1125), .B2(w1126), .A2(w1127), .C1(nHCLK1), .B1(1'b1), .A1(1'b0), .Z(w1128) );
	vdp_slatch g1243 (.Q(w1062), .D(w1120), .C(w1097), .nC(w1098) );
	vdp_slatch g1244 (.Q(w1096), .D(w1132), .C(w1097), .nC(w1098) );
	vdp_aon22 g1245 (.Z(w1099), .A1(COL[6]), .A2(w1135), .B1(w129), .B2(w1498) );
	vdp_not g1246 (.A(w1122), .nZ(w1094) );
	vdp_not g1247 (.A(w1135), .nZ(w1498) );
	vdp_and g1248 (.Z(w1), .A(w1096), .B(w1062) );
	vdp_and g1249 (.Z(w1095), .A(M5), .B(w1094) );
	vdp_and g1250 (.Z(w1499), .A(M5), .B(w1122) );
	vdp_and g1251 (.Z(128k), .A(M5), .B(w1121) );
	vdp_or3 g1252 (.Z(w1139), .A(w1136), .B(w1137), .C(w1405) );
	vdp_and g1253 (.Z(w1138), .A(w1136), .B(w1108) );
	vdp_nand g1254 (.Z(w1146), .A(w1144), .B(w1139) );
	vdp_nand g1255 (.Z(w1145), .A(w1144), .B(w1142) );
	vdp_slatch g1256 (.Q(w91), .D(w612), .C(w1123), .nC(w1124) );
	vdp_slatch g1257 (.Q(w93), .D(w685), .C(w1123), .nC(w1124) );
	vdp_slatch g1258 (.Q(w44), .D(w698), .C(w1123), .nC(w1124) );
	vdp_slatch g1259 (.Q(w1147), .D(w719), .C(w1123), .nC(w1124) );
	vdp_slatch g1260 (.Q(w111), .D(w725), .C(w1123), .nC(w1124) );
	vdp_slatch g1261 (.Q(w94), .D(w681), .C(w1123), .nC(w1124) );
	vdp_slatch g1262 (.Q(w1074), .D(w661), .C(w1123), .nC(w1124) );
	vdp_slatch g1263 (.Q(w1131), .D(w617), .C(w1123), .nC(w1124) );
	vdp_slatch g1264 (.Q(w1122), .D(w719), .C(w1130), .nC(w1129) );
	vdp_slatch g1265 (.Q(w1121), .D(w617), .C(w1130), .nC(w1129) );
	vdp_slatch g1266 (.Q(w19), .D(w725), .C(w1133), .nC(w1134) );
	vdp_slatch g1267 (.Q(w89), .D(w719), .C(w1133), .nC(w1134) );
	vdp_slatch g1268 (.Q(w1132), .D(w698), .C(w1133), .nC(w1134) );
	vdp_slatch g1269 (.Q(w1120), .D(w685), .C(w1133), .nC(w1134) );
	vdp_slatch g1270 (.Q(H40), .D(w612), .C(w1133), .nC(w1134) );
	vdp_slatch g1271 (.Q(w45), .D(w612), .C(w1130), .nC(w1129) );
	vdp_slatch g1272 (.Q(w132), .D(w685), .C(w1130), .nC(w1129) );
	vdp_slatch g1273 (.Q(M5), .D(w698), .C(w1130), .nC(w1129) );
	vdp_slatch g1274 (.Q(w1149), .D(w725), .C(w1130), .nC(w1129) );
	vdp_slatch g1275 (.Q(w1148), .D(w681), .C(w1130), .nC(w1129) );
	vdp_slatch g1276 (.Q(w1119), .D(w661), .C(w1130), .nC(w1129) );
	vdp_and g1277 (.Z(w119), .A(w1076), .B(w1158) );
	vdp_and g1278 (.Z(w123), .A(w1027), .B(w1158) );
	vdp_and g1279 (.Z(w118), .A(w1076), .B(w1159) );
	vdp_and g1280 (.Z(w122), .A(w1027), .B(w1159) );
	vdp_and g1281 (.Z(w120), .A(w1076), .B(w1153) );
	vdp_and g1282 (.Z(w121), .A(w1027), .B(w1153) );
	vdp_and g1283 (.Z(w57), .A(w1076), .B(w1154) );
	vdp_and g1284 (.Z(w48), .A(w1027), .B(w1154) );
	vdp_and g1285 (.Z(w90), .A(w1076), .B(w1156) );
	vdp_and g1286 (.Z(w88), .A(w1027), .B(w1156) );
	vdp_and g1287 (.Z(w92), .A(w1076), .B(w1157) );
	vdp_and g1288 (.Z(w1152), .A(w1027), .B(w1157) );
	vdp_and g1289 (.Z(w1175), .A(w1076), .B(w1161) );
	vdp_and g1290 (.Z(w1150), .A(w1076), .B(w1162) );
	vdp_and g1291 (.Z(w56), .A(w1076), .B(w1155) );
	vdp_and g1292 (.Z(w54), .A(w1027), .B(w1155) );
	vdp_dslatch g1293 (.D(COL[0]), .C(HCLK1), .Q(w1100), .nC(nHCLK1) );
	vdp_dslatch g1294 (.D(COL[1]), .Q(w1110), .C(HCLK1), .nC(nHCLK1) );
	vdp_dslatch g1295 (.D(COL[2]), .Q(w1528), .C(HCLK1), .nC(nHCLK1) );
	vdp_dslatch g1296 (.D(COL[3]), .Q(w1107), .C(HCLK1), .nC(nHCLK1) );
	vdp_dslatch g1297 (.D(COL[4]), .Q(w1103), .C(HCLK1), .nC(nHCLK1) );
	vdp_dslatch g1298 (.D(COL[5]), .Q(w1104), .C(HCLK1), .nC(nHCLK1) );
	vdp_dslatch g1299 (.D(w1099), .Q(w1105), .C(HCLK1), .nC(nHCLK1) );
	vdp_dslatch g1300 (.D(w130), .Q(w1106), .C(HCLK1), .nC(nHCLK1) );
	vdp_slatch g1301 (.Q(w52), .D(w681), .C(w1134), .nC(w1133) );
	vdp_slatch g1302 (.Q(w39), .D(w661), .C(w1134), .nC(w1133) );
	vdp_slatch g1303 (.Q(w1151), .D(w617), .C(w1134), .nC(w1133) );
	vdp_slatch g1304 (.Q(w23), .D(w719), .nC(w1183), .C(w1181) );
	vdp_slatch g1305 (.Q(w97), .D(w698), .nC(w1183), .C(w1181) );
	vdp_slatch g1306 (.Q(w477), .D(w685), .nC(w1183), .C(w1181) );
	vdp_slatch g1307 (.Q(w53), .D(w612), .nC(w1183), .C(w1181) );
	vdp_slatch g1308 (.Q(w95), .D(w617), .nC(w1183), .C(w1181) );
	vdp_slatch g1309 (.Q(w96), .D(w661), .nC(w1183), .C(w1181) );
	vdp_slatch g1310 (.Q(w59), .D(w681), .nC(w1183), .C(w1181) );
	vdp_slatch g1311 (.Q(w1180), .D(w725), .nC(w1183), .C(w1181) );
	vdp_slatch_r g1312 (.Q(w124), .D(DB[14]), .nC(w1174), .R(w1170), .C(w1178) );
	vdp_slatch_r g1313 (.Q(w128), .D(DB[13]), .R(w1170), .nC(w1174), .C(w1178) );
	vdp_slatch_r g1314 (.Q(w125), .D(DB[12]), .R(w1170), .nC(w1174), .C(w1178) );
	vdp_comp_str g1315 (.Z(w1181), .A(w1179), .nZ(w1183) );
	vdp_comp_str g1316 (.Z(w1177), .A(w1150), .nZ(w1176) );
	vdp_not g1317 (.A(w661), .nZ(w1496) );
	vdp_not g1318 (.A(w617), .nZ(w1198) );
	vdp_not g1319 (.A(w725), .nZ(w1184) );
	vdp_not g1320 (.A(w681), .nZ(w1182) );
	vdp_not g1321 (.A(w698), .nZ(w1199) );
	vdp_not g1322 (.A(w719), .nZ(w1185) );
	vdp_not g1323 (.A(w612), .nZ(w1193) );
	vdp_not g1324 (.A(w685), .nZ(w1194) );
	vdp_not g1325 (.A(w1168), .nZ(w1187) );
	vdp_not g1326 (.A(w1169), .nZ(w1172) );
	vdp_not g1327 (.A(w1160), .nZ(w1186) );
	vdp_not g1328 (.A(w1173), .nZ(w1188) );
	vdp_comp_str g1329 (.Z(DB[9]), .nZ(w1171), .A(w1077) );
	vdp_slatch_r g1330 (.Q(w1173), .R(w1170), .D(w325), .nC(w1171), .C(DB[9]) );
	vdp_slatch_r g1331 (.Q(w1160), .D(DB[10]), .nC(w1171), .R(w1170), .C(DB[9]) );
	vdp_and4 g1332 (.Z(w1505), .A(w1168), .B(w1169), .C(w1173), .D(w1160) );
	vdp_and4 g1333 (.Z(w1153), .A(w1173), .B(w1186), .C(w1172), .D(w1187) );
	vdp_and4 g1334 (.Z(w1159), .A(w1188), .B(w1160), .C(w1169), .D(w1168) );
	vdp_and4 g1335 (.Z(w1158), .A(w1188), .B(w1160), .C(w1169), .D(w1187) );
	vdp_and4 g1336 (.Z(w1157), .A(w1188), .B(w1160), .C(w1172), .D(w1168) );
	vdp_and4 g1337 (.Z(w1156), .A(w1188), .B(w1160), .C(w1172), .D(w1187) );
	vdp_and4 g1338 (.Z(w1154), .A(w1188), .B(w1186), .C(w1169), .D(w1168) );
	vdp_and4 g1339 (.Z(w1155), .A(w1188), .B(w1186), .C(w1169), .D(w1187) );
	vdp_and4 g1340 (.Z(w1162), .A(w1188), .B(w1186), .C(w1172), .D(w1168) );
	vdp_and4 g1341 (.Z(w1161), .A(w1188), .B(w1186), .C(w1172), .D(w1187) );
	vdp_nand g1342 (.Z(w1442), .A(w1505), .B(w1076) );
	vdp_slatch_r g1343 (.Q(w1168), .D(DB[8]), .R(w1170), .C(DB[9]), .nC(w1171) );
	vdp_slatch_r g1344 (.Q(w1167), .D(w325), .R(w1170), .C(w1178), .nC(w1174) );
	vdp_slatch_r g1345 (.nC(w1190), .Q(w1169), .D(DB[9]), .R(w1170), .C(w1171) );
	vdp_slatch_r g1346 (.Q(w1166), .D(DB[10]), .R(w1170), .C(w1178), .nC(w1174) );
	vdp_slatch_r g1347 (.Q(w99), .D(DB[8]), .R(w1170), .C(w1178), .nC(w1174) );
	vdp_slatch_r g1348 (.Q(w1165), .D(DB[9]), .R(w1170), .C(w1178), .nC(w1174) );
	vdp_slatch_r g1349 (.Q(w98), .D(w160), .R(w1170), .C(w1178), .nC(w1174) );
	vdp_slatch_r g1350 (.Q(w100), .D(DB[5]), .R(w1170), .C(w1178), .nC(w1174) );
	vdp_slatch_r g1351 (.Q(w101), .D(DB[6]), .R(w1170), .C(w1178), .nC(w1174) );
	vdp_slatch_r g1352 (.Q(w972), .D(DB[4]), .R(w1170), .C(w1178), .nC(w1174) );
	vdp_slatch_r g1353 (.Q(w1196), .D(DB[2]), .R(w1170), .C(w1178), .nC(w1174) );
	vdp_slatch_r g1354 (.Q(w1197), .D(w156), .R(w1170), .C(w1178), .nC(w1174) );
	vdp_slatch_r g1355 (.Q(w1135), .D(DB[0]), .R(w1170), .C(w1178), .nC(w1174) );
	vdp_slatch_r g1356 (.Q(w798), .D(DB[1]), .R(w1170), .C(w1178), .nC(w1174) );
	vdp_slatch_r g1357 (.Q(w105), .D(DB[9]), .R(w1170), .C(w1177), .nC(w1176) );
	vdp_slatch_r g1358 (.Q(w106), .D(DB[10]), .R(w1170), .C(w1177), .nC(w1176) );
	vdp_slatch_r g1359 (.Q(w103), .D(w160), .R(w1170), .C(w1177), .nC(w1176) );
	vdp_slatch_r g1360 (.Q(w104), .D(DB[8]), .R(w1170), .C(w1177), .nC(w1176) );
	vdp_slatch_r g1361 (.Q(w51), .D(DB[5]), .R(w1170), .C(w1177), .nC(w1176) );
	vdp_slatch_r g1362 (.Q(w41), .D(DB[6]), .R(w1170), .C(w1177), .nC(w1176) );
	vdp_slatch_r g1363 (.Q(w40), .D(w156), .R(w1170), .C(w1177), .nC(w1176) );
	vdp_slatch_r g1364 (.Q(w42), .D(DB[4]), .R(w1170), .C(w1177), .nC(w1176) );
	vdp_slatch_r g1365 (.Q(w1497), .D(DB[1]), .R(w1170), .C(w1177), .nC(w1176) );
	vdp_slatch_r g1366 (.Q(w55), .D(DB[2]), .R(w1170), .C(w1177), .nC(w1176) );
	vdp_slatch_r g1367 (.Q(w43), .D(DB[0]), .R(w1170), .C(w1177), .nC(w1176) );
	vdp_comp_str g1368 (.Z(w1178), .nZ(w1174), .A(w1175) );
	vdp_notif0 g1369 (.A(VPOS[9]), .nZ(DB[10]), .nE(w1191) );
	vdp_notif0 g1370 (.A(VPOS[8]), .nZ(DB[9]), .nE(w1191) );
	vdp_bufif0 g1371 (.A(w593), .Z(DB[9]), .nE(w1224) );
	vdp_bufif0 g1372 (.A(w675), .Z(DB[8]), .nE(w1224) );
	vdp_bufif0 g1373 (.A(w1223), .Z(DB[1]), .nE(w1224) );
	vdp_bufif0 g1374 (.A(w1225), .Z(DB[0]), .nE(w1224) );
	vdp_bufif0 g1375 (.A(w1204), .Z(w160), .nE(w1224) );
	vdp_bufif0 g1376 (.A(w1203), .Z(DB[6]), .nE(w1224) );
	vdp_bufif0 g1377 (.A(w1202), .Z(DB[5]), .nE(w1224) );
	vdp_bufif0 g1378 (.A(ODD/EVEN), .Z(DB[4]), .nE(w1224) );
	vdp_bufif0 g1379 (.A(w46), .Z(w156), .nE(w1224) );
	vdp_bufif0 g1380 (.A(w21), .Z(DB[2]), .nE(w1224) );
	vdp_slatch_r g1381 (.Q(w80), .D(DB[4]), .R(w1170), .C(w1171), .nC(w1190) );
	vdp_slatch_r g1382 (.Q(w81), .D(DB[5]), .R(w1170), .C(w1171), .nC(w1190) );
	vdp_slatch_r g1383 (.Q(w83), .D(w160), .R(w1170), .C(w1171), .nC(w1190) );
	vdp_slatch_r g1384 (.Q(w82), .D(DB[6]), .R(w1170), .C(w1171), .nC(w1190) );
	vdp_slatch_r g1385 (.Q(w76), .D(DB[0]), .R(w1170), .C(w1171), .nC(w1190) );
	vdp_slatch_r g1386 (.Q(w77), .D(DB[1]), .R(w1170), .C(w1171), .nC(w1190) );
	vdp_slatch_r g1387 (.Q(w79), .D(w156), .R(w1170), .C(w1171), .nC(w1190) );
	vdp_slatch_r g1388 (.Q(w78), .D(DB[2]), .R(w1170), .C(w1171), .nC(w1190) );
	vdp_notif0 g1389 (.A(HPOS[0]), .nZ(DB[8]), .nE(w1191) );
	vdp_not g1390 (.A(w407), .nZ(w1506) );
	vdp_comp_str g1391 (.Z(w1192), .A(w806), .nZ(w1195) );
	vdp_slatch_r g1392 (.Q(w1208), .D(w1193), .R(w1211), .C(w1192), .nC(w1195) );
	vdp_slatch_r g1393 (.Q(w1219), .D(w1199), .R(w1211), .C(w1192), .nC(w1195) );
	vdp_slatch_r g1394 (.Q(w1226), .D(w1194), .R(w1211), .C(w1192), .nC(w1195) );
	vdp_slatch_r g1395 (.Q(w1213), .D(w1496), .R(w1211), .C(w1192), .nC(w1195) );
	vdp_slatch_r g1396 (.Q(w1220), .D(w1185), .R(w1211), .C(w1192), .nC(w1195) );
	vdp_slatch_r g1397 (.Q(w1212), .D(w1182), .R(w1211), .C(w1192), .nC(w1195) );
	vdp_slatch_r g1398 (.Q(w1221), .D(w1184), .R(w1211), .C(w1192), .nC(w1195) );
	vdp_slatch_r g1399 (.Q(w1214), .D(w1198), .R(w1211), .C(w1192), .nC(w1195) );
	vdp_aon22 g1400 (.Z(w1223), .A1(w593), .A2(w1206), .B1(w1207), .B2(DMA_BUSY) );
	vdp_aon22 g1401 (.Z(w1225), .A1(w675), .A2(w1206), .B1(w1207), .B2(w1205) );
	vdp_and3 g1402 (.C(w1196), .A(w410), .B(w1506), .Z(w1201) );
	vdp_not g1403 (.A(w1201), .nZ(w1191) );
	vdp_not g1404 (.A(w1008), .nZ(w1224) );
	vdp_cnt_bit_load g1405 (.V(w1214), .nL(w1231), .L(w1209), .R(1'b0), .Q(w1232), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1260) );
	vdp_cnt_bit_load g1406 (.V(w1213), .nL(w1231), .L(w1209), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1538), .CO(w1260) );
	vdp_cnt_bit_load g1407 (.V(w1212), .nL(w1231), .L(w1209), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1259), .CO(w1538) );
	vdp_cnt_bit_load g1408 (.V(w1221), .nL(w1231), .L(w1209), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1258), .CO(w1259) );
	vdp_cnt_bit_load g1409 (.V(w1220), .nL(w1231), .L(w1209), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1257), .CO(w1258) );
	vdp_cnt_bit_load g1410 (.V(w1219), .nL(w1231), .L(w1209), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1548), .CO(w1257) );
	vdp_cnt_bit_load g1411 (.V(w1226), .nL(w1231), .L(w1209), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1256), .CO(w1548) );
	vdp_cnt_bit_load g1412 (.V(w1208), .nL(w1231), .L(w1209), .R(1'b0), .CI(w1228), .CO(w1256), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g1413 (.D(w1502), .C2(HCLK2), .C1(HCLK1), .Q(w1233), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_rs_FF g1414 (.Q(w1203), .R(w1249), .S(w1250) );
	vdp_rs_FF g1415 (.Q(w1204), .R(w1248), .S(w112) );
	vdp_rs_FF g1416 (.Q(w1202), .R(w1249), .S(w126) );
	vdp_not g1417 (.A(M5), .nZ(w1247) );
	vdp_not g1418 (.A(w1204), .nZ(w1227) );
	vdp_not g1419 (.A(w1210), .nZ(w1216) );
	vdp_not g1420 (.A(CA[21]), .nZ(w1503) );
	vdp_not g1421 (.A(w407), .nZ(w1217) );
	vdp_not g1422 (.A(w1252), .nZ(w1218) );
	vdp_comp_we g1423 (.Z(w1231), .A(w1501), .nZ(w1209) );
	vdp_or g1424 (.A(w1252), .B(w1233), .Z(w1501) );
	vdp_and g1425 (.A(w1218), .B(w1232), .Z(w1502) );
	vdp_and g1426 (.A(w1227), .B(w127), .Z(w1250) );
	vdp_or g1427 (.A(w1197), .B(w4), .Z(w1228) );
	vdp_not g1428 (.A(w1206), .nZ(w1207) );
	vdp_nor3 g1429 (.A(w407), .B(w1247), .Z(w1206), .C(CA[1]) );
	vdp_nor3 g1430 (.A(w1197), .B(w5), .Z(w1252), .C(w31) );
	vdp_nor g1431 (.A(w1255), .B(w1234), .Z(w1215) );
	vdp_or5 g1432 (.A(w1217), .B(CA[4]), .C(CA[5]), .D(CA[15]), .Z(w1255), .E(CA[6]) );
	vdp_or5 g1433 (.A(CA[16]), .B(CA[17]), .C(CA[20]), .D(w1216), .Z(w1234), .E(w1503) );
	vdp_rs_FF g1434 (.Q(w1240), .R(w1293), .S(w1502) );
	vdp_rs_FF g1435 (.Q(w1294), .R(w1277), .S(w1504) );
	vdp_dff g1436 (.Q(w1297), .R(w1253), .C(w1243), .D(w1236) );
	vdp_dff g1437 (.Q(w1296), .R(w1253), .C(w1243), .D(w1235) );
	vdp_dff g1438 (.Q(w1298), .R(w1253), .C(w1243), .D(w1237) );
	vdp_rs_FF g1439 (.Q(w1554), .R(w1292), .S(w1553) );
	vdp_rs_FF g1440 (.Q(w1264), .R(w1265), .S(w1551) );
	vdp_dlatch_inv g1441 (.D(w1271), .Q(w1272), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g1442 (.D(w1265), .C(DCLK1), .Q(w1271), .nC(nDCLK1) );
	vdp_dlatch_inv g1443 (.D(w1275), .Q(w1249), .C(HCLK1), .nC(nHCLK1) );
	vdp_not g1444 (.A(w1288), .nZ(w1261) );
	vdp_not g1445 (.A(w673), .nZ(w1239) );
	vdp_not g1446 (.A(w1242), .nZ(w1237) );
	vdp_not g1447 (.A(w1241), .nZ(w1236) );
	vdp_not g1448 (.A(w1251), .nZ(w1253) );
	vdp_not g1449 (.A(w1268), .nZ(w1243) );
	vdp_not g1450 (.A(w1244), .nZ(w50) );
	vdp_not g1451 (.A(w1246), .nZ(w1245) );
	vdp_sr_bit g1452 (.D(w1273), .C2(HCLK2), .C1(HCLK1), .Q(w1292), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and g1453 (.A(M5), .B(w1264), .Z(w1268) );
	vdp_and g1454 (.A(w407), .B(w1263), .Z(w1083) );
	vdp_and g1455 (.A(w1244), .B(w1083), .Z(w1552) );
	vdp_or g1456 (.A(w428), .B(w1552), .Z(w1551) );
	vdp_or g1457 (.A(w1008), .B(SYSRES), .Z(w1553) );
	vdp_and g1458 (.A(w1247), .B(w1249), .Z(w1276) );
	vdp_or g1459 (.A(w1296), .B(w1276), .Z(w1277) );
	vdp_and g1460 (.A(M5), .B(w474), .Z(w1504) );
	vdp_and g1461 (.A(w1149), .B(M5), .Z(w1238) );
	vdp_or g1462 (.A(w1298), .B(w1276), .Z(w1248) );
	vdp_or g1463 (.A(w1297), .B(w1276), .Z(w1293) );
	vdp_comp_DFF g1464 (.D(w1554), .C2(HCLK2), .C1(HCLK1), .Q(w1273), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_comp_DFF g1465 (.D(w1268), .C2(DCLK2), .C1(DCLK1), .Q(w1265), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_nor g1466 (.A(w1273), .B(SYSRES), .Z(w1274) );
	vdp_nand g1467 (.A(w1292), .B(w1274), .Z(w1275) );
	vdp_nand g1468 (.A(w1204), .B(w1148), .Z(w1242) );
	vdp_and3 g1469 (.A(w1238), .B(w933), .Z(w1287), .C(w1239) );
	vdp_and3 g1470 (.A(w1238), .B(w933), .Z(w1286), .C(w673) );
	vdp_and4 g1471 (.A(w1241), .B(w1147), .C(w1242), .D(w1294), .Z(w1235) );
	vdp_nand3 g1472 (.C(w1240), .A(w1242), .B(w1180), .Z(w1241) );
	vdp_aoi21 g1473 (.A1(w1272), .B(SYSRES), .Z(w1251), .A2(w1271) );
	vdp_dff g1474 (.Q(w1317), .R(w1303), .C(w1300), .D(w1285) );
	vdp_dff g1475 (.Q(w1313), .R(w1303), .C(w1300), .D(w1312) );
	vdp_dff g1476 (.Q(w1282), .R(w1303), .C(w1300), .D(w1280) );
	vdp_dff g1477 (.Q(w1290), .R(w1303), .C(w1300), .D(w1289) );
	vdp_dff g1478 (.Q(w1291), .R(w1303), .C(w1300), .D(w1279) );
	vdp_dff g1479 (.Q(w1269), .R(w1303), .C(w1300), .D(w1308) );
	vdp_dff g1480 (.Q(w1266), .R(w1303), .C(w1300), .D(w1306) );
	vdp_dff g1481 (.Q(w1299), .R(1'b0), .C(w1300), .D(w1262) );
	vdp_ha g1482 (.SUM(w1306), .A(w1266), .B(w1261), .CO(w1267) );
	vdp_ha g1483 (.SUM(w1308), .A(w1269), .B(w1267), .CO(w1270) );
	vdp_ha g1484 (.SUM(w1279), .A(w1291), .B(w1270), .CO(w1278) );
	vdp_ha g1485 (.SUM(w1289), .A(w1290), .B(w1278), .CO(w1283) );
	vdp_ha g1486 (.SUM(w1280), .A(w1282), .B(w1283), .CO(w1281) );
	vdp_ha g1487 (.SUM(w1285), .A(w1317), .B(w1281), .CO(w1284) );
	vdp_ha g1488 (.SUM(w1312), .A(w1313), .B(w1284) );
	vdp_and3 g1489 (.A(w1313), .B(w1282), .Z(w1310), .C(w1317) );
	vdp_and4 g1490 (.C(w1269), .A(w1290), .B(w1310), .Z(w1316), .D(w1291) );
	vdp_nand g1491 (.A(w1299), .B(w407), .Z(w1440) );
	vdp_dff g1492 (.Q(w1325), .R(1'b0), .C(w1300), .D(w1305) );
	vdp_dff g1493 (.Q(w1305), .R(w1307), .C(w1300), .D(w1330) );
	vdp_dff g1494 (.Q(w1330), .R(w1307), .C(w1328), .D(w1309) );
	vdp_dff g1495 (.Q(w1309), .R(w1307), .C(w1300), .D(w1334) );
	vdp_dff g1496 (.Q(w1334), .R(w1307), .C(w1300), .D(w1335) );
	vdp_dff g1497 (.Q(w1335), .R(w1307), .C(w1300), .D(1'b1) );
	vdp_dff g1498 (.Q(w1541), .R(w1344), .C(w1318), .D(w1310) );
	vdp_dff g1499 (.Q(w1318), .R(1'b0), .C(w1300), .D(w1316) );
	vdp_dff g1500 (.Q(w1337), .R(w1315), .C(w1338), .D(w1310) );
	vdp_dff g1501 (.Q(w1314), .R(w1329), .C(w1342), .D(1'b1) );
	vdp_or g1502 (.A(SYSRES), .B(w1314), .Z(w1315) );
	vdp_or g1503 (.A(w1307), .B(w1325), .Z(w1340) );
	vdp_not g1504 (.A(w1325), .nZ(w1302) );
	vdp_not g1505 (.A(w1541), .nZ(w1307) );
	vdp_nand3 g1506 (.A(w407), .B(w1323), .Z(w1303), .C(w1302) );
	vdp_not g1507 (.nZ(w1328), .A(w1324) );
	vdp_not g1508 (.nZ(w1300), .A(w1301) );
	vdp_dff g1509 (.Q(w1327), .R(1'b0), .C(w1328), .D(w1350) );
	vdp_dff g1510 (.Q(w1353), .R(w1329), .C(w1328), .D(w1333) );
	vdp_dff g1511 (.Q(w1333), .R(w1329), .C(w1300), .D(w1355) );
	vdp_dff g1512 (.Q(w1355), .R(w1329), .C(w1328), .D(w1332) );
	vdp_dff g1513 (.Q(w1332), .R(w1329), .C(w1328), .D(w1343) );
	vdp_dff g1514 (.Q(w1343), .R(w1329), .C(w1300), .D(w47) );
	vdp_dff g1515 (.Q(w1360), .R(w1359), .C(w1328), .D(w1137) );
	vdp_dff g1516 (.Q(w1137), .R(w1359), .C(w1300), .D(w1339) );
	vdp_not g1517 (.A(w1347), .nZ(w113) );
	vdp_not g1518 (.A(w1006), .nZ(w1322) );
	vdp_not g1519 (.A(w1333), .nZ(w1331) );
	vdp_not g1520 (.A(w1330), .nZ(w1549) );
	vdp_not g1521 (.A(w1339), .nZ(w1359) );
	vdp_not g1522 (.A(w1083), .nZ(w1342) );
	vdp_not g1523 (.A(w1244), .nZ(w1542) );
	vdp_and g1524 (.A(w1340), .B(w1083), .Z(w1339) );
	vdp_and g1525 (.A(w1341), .B(w1339), .Z(w1338) );
	vdp_and g1526 (.A(w1360), .B(w1338), .Z(w47) );
	vdp_and g1527 (.A(w1334), .B(w1549), .Z(w1351) );
	vdp_and g1528 (.A(w1335), .B(w1549), .Z(w1352) );
	vdp_and g1529 (.A(w1326), .B(w996), .Z(w1349) );
	vdp_and g1530 (.A(w1326), .B(w1039), .Z(w1321) );
	vdp_and g1531 (.A(w1006), .B(w1327), .Z(w1326) );
	vdp_and g1532 (.A(w113), .B(w1137), .Z(w1071) );
	vdp_nand g1533 (.A(w1332), .B(w1331), .Z(w1323) );
	vdp_nor g1534 (.A(w1329), .B(w1343), .Z(w1354) );
	vdp_or3 g1535 (.C(w1337), .A(SYSRES), .B(w1325), .Z(w1344) );
	vdp_oai21 g1536 (.A1(w1039), .B(w1322), .Z(w1347), .A2(w996) );
	vdp_dff g1537 (.Q(w1368), .R(1'b0), .C(w1300), .D(w1246) );
	vdp_rs_FF g1538 (.nQ(w1080), .R(w1369), .S(w1366) );
	vdp_not g1539 (.A(w1374), .nZ(w1061) );
	vdp_not g1540 (.A(w617), .nZ(w1365) );
	vdp_and3 g1541 (.C(w1365), .A(w831), .B(M5), .Z(w1366) );
	vdp_or g1542 (.A(w1246), .B(SYSRES), .Z(w1369) );
	vdp_and g1543 (.A(w1386), .B(w594), .Z(w1387) );
	vdp_not g1544 (.A(w1341), .nZ(w1389) );
	vdp_and4 g1545 (.C(CA[21]), .A(w1210), .B(CA[20]), .Z(w1341), .D(w1542) );
	vdp_dff g1546 (.Q(w1429), .R(1'b0), .C(w1374), .D(w1414) );
	vdp_dff g1547 (.Q(w1409), .R(1'b0), .C(w1374), .D(w1408) );
	vdp_dff g1548 (.Q(w1348), .R(1'b0), .C(w1395), .D(w1396) );
	vdp_dff g1549 (.Q(w1408), .R(1'b0), .C(w1395), .D(w1348) );
	vdp_dff g1550 (.Q(w1421), .R(w1422), .C(HCLK2), .D(w1424) );
	vdp_dff g1551 (.Q(DMA_BUSY), .R(w1422), .C(HCLK2), .D(w1421) );
	vdp_rs_FF g1552 (.Q(w1288), .R(w1422), .S(w1357) );
	vdp_rs_FF g1553 (.Q(w1543), .R(w1422), .S(w1286) );
	vdp_rs_FF g1554 (.Q(w1262), .R(w1358), .S(w1287) );
	vdp_sr_bit g1555 (.D(w594), .Q(w1386), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1556 (.D(w1550), .Q(w1420), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_dlatch_inv g1557 (.D(w1385), .nQ(w1363), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g1558 (.D(w1384), .nQ(w1385), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g1559 (.D(w1371), .C(HCLK1), .nQ(w1384), .nC(nHCLK1) );
	vdp_aon22 g1560 (.Z(w1416), .A2(w1362), .B1(w1384), .B2(w1425), .A1(w1363) );
	vdp_sr_bit g1561 (.D(w1426), .Q(w1431), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1562 (.D(w1388), .Q(w1426), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1563 (.D(VRAM_REFRESH), .C2(HCLK2), .C1(HCLK1), .Q(w1388), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_aon22 g1564 (.Z(w1404), .A2(w1354), .B1(w1432), .B2(w1435), .A1(w1402) );
	vdp_not g1565 (.A(w1540), .nZ(w1073) );
	vdp_not g1566 (.A(w1354), .nZ(w1435) );
	vdp_not g1567 (.A(w1420), .nZ(w1425) );
	vdp_not g1568 (.A(w1361), .nZ(w1403) );
	vdp_not g1569 (.A(w1337), .nZ(w1329) );
	vdp_or g1570 (.A(w1288), .B(w1543), .Z(w1424) );
	vdp_or g1571 (.A(SYSRES), .B(w596), .Z(w1422) );
	vdp_or g1572 (.A(w1357), .B(w1422), .Z(w1358) );
	vdp_or g1573 (.A(w1237), .B(w1235), .Z(w279) );
	vdp_or g1574 (.A(w1237), .B(w1236), .Z(w254) );
	vdp_and g1575 (.A(w1420), .B(w647), .Z(w1362) );
	vdp_or g1576 (.A(w1363), .B(w1426) );
	vdp_and g1577 (.A(w1323), .B(w1338), .Z(w1402) );
	vdp_and g1578 (.A(w1355), .B(w1338), .Z(w1432) );
	vdp_and g1579 (.A(w1338), .B(w1329), .Z(w115) );
	vdp_and g1580 (.A(w1000), .B(w116), .Z(w1415) );
	vdp_or g1581 (.A(w1349), .B(w1005), .Z(w1411) );
	vdp_aon22 g1582 (.Z(w1419), .A2(w1074), .B1(w1356), .B2(w1407), .A1(w1406) );
	vdp_and g1583 (.A(w1414), .B(w1429), .Z(w1136) );
	vdp_and g1584 (.A(w1427), .B(w1436), .Z(w1417) );
	vdp_and g1585 (.A(w1436), .B(w1430), .Z(w1414) );
	vdp_not g1586 (.A(w1430), .nZ(w1427) );
	vdp_not g1587 (.A(w1428), .nZ(w1436) );
	vdp_not g1588 (.A(w1385), .nZ(w1423) );
	vdp_not g1589 (.A(w1400), .nZ(w1418) );
	vdp_and g1590 (.A(w1412), .B(w1376), .Z(w1375) );
	vdp_and g1591 (.A(w1412), .B(w1378), .Z(w999) );
	vdp_and g1592 (.A(w1412), .B(w1380), .Z(w1005) );
	vdp_and g1593 (.A(w1412), .B(w1377), .Z(w1000) );
	vdp_and g1594 (.A(w1412), .B(w1379), .Z(w1396) );
	vdp_and g1595 (.A(w999), .B(w1396), .Z(w428) );
	vdp_and g1596 (.A(w407), .B(w1390), .Z(w996) );
	vdp_and g1597 (.A(w407), .B(w1381), .Z(w1039) );
	vdp_not g1598 (.A(w407), .nZ(w1412) );
	vdp_nand g1599 (.A(w1408), .B(w1409), .Z(w1430) );
	vdp_nand g1600 (.A(w675), .B(w1373), .Z(w1372) );
	vdp_nand g1601 (.A(w407), .B(w254), .Z(w1383) );
	vdp_nand g1602 (.A(w279), .B(w407), .Z(w1382) );
	vdp_or3 g1603 (.C(w1237), .A(w1236), .B(w1235), .Z(w1066) );
	vdp_and3 g1604 (.C(w1363), .A(w594), .B(w1420), .Z(w599) );
	vdp_aoi21 g1605 (.A2(w1362), .B(w1423), .Z(w1361), .A1(w1384) );
	vdp_nor g1606 (.A(w1388), .B(w1431), .Z(w1373) );
	vdp_nand g1607 (.A(w113), .B(w1389), .Z(w1400) );
	vdp_nand3 g1608 (.C(w1372), .A(w3), .B(w1387), .Z(w1371) );
	vdp_2a3oi g1609 (.A1(w1423), .B(w674), .Z(w1370), .A2(w1384), .C(w1420) );
	vdp_nor4 g1610 (.C(VRAM_REFRESH), .A(w1426), .B(w1388), .Z(w1550), .D(w1431) );
	vdp_comb1 g1611 (.A1(CA[15]), .B(w1427), .Z(w1428), .A2(CA[14]), .C(w1375) );
	vdp_aon22 g1612 (.Z(w1346), .A2(w1074), .B1(w1356), .B2(w1401), .A1(w1539) );
	vdp_not g1613 (.A(w1074), .nZ(w1356) );
	vdp_or4 g1614 (.C(w1403), .A(w1436), .B(w1402), .Z(w1539), .D(w1351) );
	vdp_or4 g1615 (.C(w1363), .A(w1418), .B(w1415), .Z(w1407), .D(w1363) );
	vdp_or3 g1616 (.C(w1404), .A(w1414), .B(w1405), .Z(w1401) );
	vdp_comb1 g1617 (.A1(w1137), .B(w1333), .Z(w1540), .A2(w1354), .C(w1338) );
	vdp_and6 g1618 (.C(w1398), .A(w1299), .B(w1397), .Z(w1357), .D(w1368), .E(w407), .F(w1342) );
	vdp_or5 g1619 (.C(w1416), .A(w1408), .B(w47), .Z(w1406), .D(w1352), .E(w1138) );
	vdp_or5 g1620 (.C(w1363), .A(w1417), .B(w114), .Z(w1410), .D(w1351), .E(w1415) );
	vdp_aoi22 g1621 (.Z(w1350), .A2(w47), .B1(w1353), .B2(w1338), .A1(w1354) );
	vdp_g1622 g1622 (.Z(w308), .A(w427) );
	vdp_g1623 g1623 (.Z(w264), .A(w427) );
	vdp_g1624 g1624 (.A(w427), .Z(w300) );
	vdp_g1625 g1625 (.A(w427), .Z(w256) );
	vdp_g1626 g1626 (.Z(w290), .A(w427) );
	vdp_g1627 g1627 (.Z(w247), .A(w427) );
	vdp_g1628 g1628 (.Z(w281), .A(w427) );
	vdp_g1629 g1629 (.Z(w239), .A(w427) );
	vdp_aon22 g1630 (.Z(w1405), .A2(w1362), .B1(w1362), .B2(w1423), .A1(w1363) );
	vdp_comp_we g1631 (.nZ(w1374), .Z(w1395), .A(w1413) );
	vdp_comp_we g1632 (.nZ(w1301), .Z(w1324), .A(w1441) );
	vdp_not g1633 (.nZ(w1630), .A(w1994) );
	vdp_not g1634 (.nZ(w1632), .A(w1633) );
	vdp_sr_bit g1635 (.Q(w5), .D(w1989), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1636 (.Q(w1638), .D(w1836), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1637 (.Q(w1614), .D(w1837), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1638 (.Q(w1670), .D(w1635), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1639 (.Q(w1615), .D(w1838), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1640 (.Q(w1619), .D(w1839), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1641 (.Q(w1815), .D(w1826), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1642 (.Q(w1646), .D(w1644), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1643 (.Q(w1643), .D(w1827), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1644 (.Q(w1620), .D(w1828), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1645 (.Q(w1653), .D(w1853), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1646 (.Q(w1651), .D(w1648), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1647 (.Q(w1648), .D(w2005), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1648 (.Q(w1652), .D(w1655), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1649 (.Q(w1625), .D(w1955), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_not g1650 (.nZ(w1644), .A(w1654) );
	vdp_not g1651 (.nZ(w58), .A(w1643) );
	vdp_not g1652 (.nZ(w1629), .A(w1643) );
	vdp_not g1653 (.nZ(w1622), .A(ODD/EVEN) );
	vdp_not g1654 (.nZ(w1631), .A(w1062) );
	vdp_not g1655 (.nZ(w2005), .A(w1990) );
	vdp_not g1656 (.nZ(w1657), .A(w1658) );
	vdp_not g1657 (.nZ(w1645), .A(w1991) );
	vdp_not g1658 (.nZ(w1650), .A(w1651) );
	vdp_not g1659 (.nZ(w1627), .A(w53) );
	vdp_and g1660 (.Z(w1649), .A(w1849), .B(w1653) );
	vdp_nor g1661 (.Z(w1647), .A(SYSRES), .B(w1619) );
	vdp_oai21 g1662 (.Z(w1990), .B(w1647), .A2(w1657), .A1(w1648) );
	vdp_oai21 g1663 (.Z(w1658), .B(w1656), .A2(w1655), .A1(w1853) );
	vdp_aoi21 g1664 (.Z(w1991), .B(SYSRES), .A2(w1652), .A1(w1849) );
	vdp_and g1665 (.Z(w1626), .A(w1629), .B(w27) );
	vdp_and3 g1666 (.Z(w1849), .A(w1650), .B(w53), .C(w1648) );
	vdp_or g1667 (.Z(w1628), .A(SYSRES), .B(w1629) );
	vdp_and g1668 (.Z(w1955), .A(w1623), .B(w1633) );
	vdp_and g1669 (.Z(w1634), .A(w1626), .B(w1627) );
	vdp_and g1670 (.Z(w1623), .A(w1626), .B(w53) );
	vdp_and g1671 (.Z(w1618), .A(w1613), .B(w1620) );
	vdp_or g1672 (.Z(w1617), .A(SYSRES), .B(w1618) );
	vdp_2?3?I g1673 (.Z(w1994), .A1(w1632), .A2(w1623), .C(SYSRES), .B(w1631) );
	vdp_or g1674 (.Z(w1613), .A(w1621), .B(w1622) );
	vdp_or g1675 (.Z(w1616), .A(SYSRES), .B(w1668) );
	vdp_and g1676 (.Z(w1668), .A(w1613), .B(w1615) );
	vdp_and g1677 (.Z(w1639), .A(w1613), .B(w1638) );
	vdp_and g1678 (.Z(w1637), .A(w1613), .B(w1614) );
	vdp_or g1679 (.Z(w1942), .A(w1668), .B(SYSRES) );
	vdp_and g1680 (.Z(w1855), .A(w1635), .B(M5) );
	vdp_not g1681 (.nZ(w46), .A(w1641) );
	vdp_not g1682 (.nZ(w1641), .A(w1640) );
	vdp_not g1683 (.nZ(w1674), .A(w1640) );
	vdp_not g1684 (.nZ(w1989), .A(w1825) );
	vdp_and g1685 (.Z(w1743), .A(M5), .B(w1636) );
	vdp_or g1686 (.Z(w1642), .A(SYSRES), .B(w1639) );
	vdp_oai21 g1687 (.Z(w1640), .B(w1119), .A2(w31), .A1(w5) );
	vdp_RS g1688 (.Q(w1636), .S(w1637), .R(w1642) );
	vdp_RS g1689 (.Q(w1624), .R(w1616), .S(w1618) );
	vdp_RS g1690 (.Q(w31), .S(w1646), .R(w1628) );
	vdp_RS g1691 (.Q(w20), .R(w1619), .S(w1617) );
	vdp_TFF g1692 (.C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .CI(w1634), .R(w1630), .A(w1625), .Q(ODD/EVEN) );
	vdp_cnt_bit_load g1693 (.D(w1845), .Q(w1707), .nL(w1972), .L(w1830), .CI(w1847), .nC1(nHCLK1), .CO(w1939), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g1694 (.Q(w1621), .D(w1933), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1695 (.Q(w2003), .D(w1950), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1696 (.Q(w32), .D(w2017), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1697 (.Q(w27), .D(w1929), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1698 (.Q(VRAM_REFRESH), .D(w1693), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1699 (.Q(w1710), .D(w1692), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1700 (.Q(w1703), .D(w1691), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1701 (.Q(w1678), .D(w1930), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1702 (.Q(w1704), .D(w1719), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1703 (.Q(w1655), .D(w1932), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1704 (.Q(w1852), .D(w1934), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1705 (.Q(w1735), .D(w1928), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1706 (.Q(w1853), .D(w1924), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1707 (.Q(w1719), .D(w1982), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1708 (.Q(w1871), .D(w1879), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1709 (.Q(w1714), .D(w1689), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1710 (.Q(w1734), .D(w1880), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1711 (.Q(w2015), .D(w2018), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1712 (.Q(w1768), .D(w1764), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1713 (.Q(w1716), .D(w1874), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1714 (.Q(w9), .D(w1873), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1715 (.Q(w1732), .D(w1778), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1716 (.Q(w1729), .D(w1931), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1717 (.Q(w1748), .D(w1878), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1718 (.Q(w1740), .D(w1755), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1719 (.Q(w1799), .D(w1744), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1720 (.Q(w29), .D(w1770), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1721 (.Q(w22), .D(w1675), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1722 (.Q(w1763), .D(w1953), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1723 (.Q(w1984), .D(w1805), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1724 (.Q(w1801), .D(w1875), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1725 (.Q(w1759), .D(w1922), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1726 (.Q(w1785), .D(w1808), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1727 (.Q(w30), .D(w1952), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1728 (.Q(w1787), .D(w1877), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1729 (.Q(w1788), .D(w1876), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1730 (.Q(w1813), .D(w1757), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1731 (.Q(w1760), .D(w1925), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1732 (.Q(w1669), .D(w2010), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1733 (.Q(w1746), .D(w2009), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1734 (.Q(w1800), .D(w1756), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1735 (.Q(w1761), .D(w1758), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1736 (.Q(w1804), .D(w1926), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1737 (.Q(w1782), .D(w1923), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1738 (.Q(w25), .D(w1676), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1739 (.Q(w1783), .D(w1669), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1740 (.Q(w1814), .D(w1769), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1741 (.Q(w1865), .D(w1921), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_not g1742 (.nZ(w1699), .A(M5) );
	vdp_not g1743 (.nZ(w6), .A(w1957) );
	vdp_not g1744 (.nZ(w7), .A(w1678) );
	vdp_not g1745 (.nZ(w1872), .A(w1673) );
	vdp_not g1746 (.nZ(w1682), .A(w53) );
	vdp_not g1747 (.nZ(w1684), .A(w1951) );
	vdp_not g1748 (.nZ(w1774), .A(w1) );
	vdp_not g1749 (.nZ(w1724), .A(w1690) );
	vdp_not g1750 (.nZ(w1705), .A(w1704) );
	vdp_not g1751 (.nZ(w1717), .A(w1678) );
	vdp_not g1752 (.nZ(w1718), .A(w44) );
	vdp_not g1753 (.nZ(w8), .A(w1712) );
	vdp_not g1754 (.nZ(w1701), .A(w39) );
	vdp_not g1755 (.nZ(w2014), .A(w53) );
	vdp_not g1756 (.nZ(w13), .A(w1978) );
	vdp_not g1757 (.nZ(w1979), .A(w1729) );
	vdp_not g1758 (.nZ(w1982), .A(w1739) );
	vdp_not g1759 (.nZ(w1773), .A(w1695) );
	vdp_not g1760 (.nZ(w2001), .A(w1694) );
	vdp_not g1761 (.nZ(w1722), .A(H40) );
	vdp_not g1762 (.nZ(w14), .A(w1771) );
	vdp_not g1763 (.nZ(w1971), .A(w1681) );
	vdp_not g1764 (.nZ(w1810), .A(w1742) );
	vdp_not g1765 (.nZ(w1789), .A(w1775) );
	vdp_not g1766 (.nZ(w1806), .A(w52) );
	vdp_not g1767 (.nZ(w1751), .A(w1927) );
	vdp_not g1768 (.nZ(w12), .A(w1958) );
	vdp_not g1769 (.nZ(w1816), .A(w1814) );
	vdp_not g1770 (.nZ(w1715), .A(w42) );
	vdp_not g1771 (.nZ(w1733), .A(w51) );
	vdp_not g1772 (.nZ(w1679), .A(w41) );
	vdp_not g1773 (.nZ(w1940), .A(w19) );
	vdp_not g1774 (.nZ(w2002), .A(w45) );
	vdp_not g1775 (.nZ(w2004), .A(M5) );
	vdp_not g1776 (.nZ(w1997), .A(w1752) );
	vdp_not g1777 (.nZ(w1829), .A(w1780) );
	vdp_not g1778 (.nZ(w1975), .A(w1949) );
	vdp_not g1779 (.nZ(w1831), .A(w1095) );
	vdp_not g1780 (.nZ(w1848), .A(w1846) );
	vdp_not g1781 (.nZ(w1842), .A(w1499) );
	vdp_not g1782 (.nZ(w1843), .A(w1205) );
	vdp_aon22 g1783 (.Z(w2023), .B1(w1833), .A1(w1832), .A2(DB[4]), .B2(w1831) );
	vdp_aon22 g1784 (.Z(w1964), .B1(w1833), .A1(w1832), .A2(DB[5]), .B2(w1820) );
	vdp_aon22 g1785 (.Z(w1965), .B1(w1833), .A1(w1832), .B2(w1975), .A2(DB[6]) );
	vdp_aon22 g1786 (.Z(w1961), .B2(1'b1), .A2(w160), .B1(w1833), .A1(w1832) );
	vdp_aon22 g1787 (.Z(w1960), .B2(1'b1), .A2(DB[8]), .B1(w1833), .A1(w1832) );
	vdp_aon22 g1788 (.Z(w1822), .B2(1'b1), .B1(w1680), .A2(DB[8]), .A1(w1954) );
	vdp_aon22 g1789 (.Z(w1974), .B2(w1819), .A2(w156), .B1(w1833), .A1(w1832) );
	vdp_aon22 g1790 (.Z(w1840), .A2(DB[2]), .B2(w1843), .B1(w1833), .A1(w1832) );
	vdp_aon22 g1791 (.Z(w1841), .A2(DB[1]), .B2(w1818), .B1(w1833), .A1(w1832) );
	vdp_aon22 g1792 (.Z(w1966), .A1(w1954), .B1(w1680), .B2(1'b1), .A2(w160) );
	vdp_aon22 g1793 (.Z(w21), .A1(w2004), .B2(w1821), .B1(M5), .A2(w1799) );
	vdp_aon22 g1794 (.Z(w1792), .B1(w1680), .A1(w1954), .A2(DB[6]), .B2(1'b1) );
	vdp_aon22 g1795 (.Z(w1767), .B1(w1783), .B2(w1784), .A2(w1866), .A1(w1781) );
	vdp_not g1796 (.nZ(w1784), .A(w1781) );
	vdp_aon22 g1797 (.Z(w1967), .B1(w1680), .A1(w1954), .B2(1'b0), .A2(w1941) );
	vdp_not g1798 (.nZ(w1811), .A(w1809) );
	vdp_aon22 g1799 (.Z(w2011), .B1(w1954), .A1(w1680), .B2(w1971), .A2(DB[4]) );
	vdp_aon22 g1800 (.Z(w1968), .B2(w1970), .B1(w1680), .A2(w156), .A1(w1954) );
	vdp_aon22 g1801 (.Z(w1765), .A2(w1727), .B2(w1709), .A1(w1767), .B1(w1766) );
	vdp_aon22 g1802 (.Z(w1969), .A2(DB[2]), .B2(w1736), .A1(w1954), .B1(w1680) );
	vdp_aon22 g1803 (.Z(w1980), .B2(w1871), .B1(w44), .A2(w1718), .A1(w1717) );
	vdp_aon22 g1804 (.Z(w1708), .B1(w1956), .A1(HCLK2), .B2(w1701), .A2(w39) );
	vdp_aon22 g1805 (.Z(w1995), .A1(w1954), .B1(w1680), .B2(w1720), .A2(DB[1]) );
	vdp_aon22 g1806 (.Z(w1685), .A2(DB[0]), .B1(w1680), .B2(w1681), .A1(w1954) );
	vdp_not g1807 (.nZ(w4), .A(w1852) );
	vdp_not g1808 (.nZ(w3), .A(w1716) );
	vdp_RS g1809 (.Q(w1762), .S(w1812), .R(w1945) );
	vdp_RS g1810 (.Q(w1798), .R(w1801), .S(w1803) );
	vdp_RS g1811 (.Q(w1744), .S(w1985), .R(w1761) );
	vdp_RS g1812 (.Q(w1943), .R(w1944), .S(w1740) );
	vdp_RS g1813 (.Q(w1745), .R(w1735), .S(w2008) );
	vdp_aon22 g1814 (.Z(w1845), .A2(DB[0]), .B2(w1817), .B1(w1833), .A1(w1832) );
	vdp_notif0 g1815 (.nZ(DB[1]), .A(VRAM_REFRESH), .nE(w1696) );
	vdp_notif0 g1816 (.nZ(DB[0]), .A(w32), .nE(w1696) );
	vdp_notif0 g1817 (.nZ(w160), .A(w27), .nE(w1697) );
	vdp_notif0 g1818 (.A(w7), .nZ(DB[6]), .nE(w1697) );
	vdp_notif0 g1819 (.A(w6), .nZ(DB[2]), .nE(w1696) );
	vdp_notif0 g1820 (.A(w8), .nZ(w156), .nE(w1696) );
	vdp_notif0 g1821 (.nZ(DB[5]), .A(w14), .nE(w1696) );
	vdp_notif0 g1822 (.A(w13), .nZ(DB[4]), .nE(w1696) );
	vdp_notif0 g1823 (.A(w16), .nZ(DB[5]), .nE(w1697) );
	vdp_notif0 g1824 (.nZ(w160), .A(w9), .nE(w1696) );
	vdp_notif0 g1825 (.nZ(DB[6]), .A(w3), .nE(w1696) );
	vdp_notif0 g1826 (.nZ(DB[4]), .A(w17), .nE(w1697) );
	vdp_notif0 g1827 (.nZ(DB[9]), .A(w29), .nE(w1696) );
	vdp_notif0 g1828 (.nZ(DB[8]), .A(w22), .nE(w1696) );
	vdp_notif0 g1829 (.nZ(w156), .A(w11), .nE(w1697) );
	vdp_notif0 g1830 (.nZ(DB[2]), .A(w28), .nE(w1697) );
	vdp_notif0 g1831 (.nZ(DB[10]), .A(w30), .nE(w1696) );
	vdp_notif0 g1832 (.nZ(w325), .A(w12), .nE(w1696) );
	vdp_notif0 g1833 (.nZ(DB[12]), .A(w24), .nE(w1696) );
	vdp_notif0 g1834 (.nZ(DB[13]), .A(w25), .nE(w1696) );
	vdp_notif0 g1835 (.nZ(DB[1]), .A(w15), .nE(w1697) );
	vdp_notif0 g1836 (.nZ(DB[0]), .A(w10), .nE(w1697) );
	vdp_not g1837 (.nZ(VPOS[9]), .A(w1963) );
	vdp_not g1838 (.nZ(VPOS[8]), .A(w1962) );
	vdp_not g1839 (.nZ(VPOS[7]), .A(w1753) );
	vdp_not g1840 (.nZ(HPOS[7]), .A(w1997) );
	vdp_not g1841 (.nZ(HPOS[8]), .A(w1829) );
	vdp_not g1842 (.nZ(HPOS[6]), .A(w1751) );
	vdp_not g1843 (.nZ(VPOS[6]), .A(w1998) );
	vdp_not g1844 (.nZ(VPOS[5]), .A(w1999) );
	vdp_not g1845 (.nZ(HPOS[5]), .A(w1789) );
	vdp_not g1846 (.nZ(HPOS[4]), .A(w1810) );
	vdp_not g1847 (.nZ(VPOS[4]), .A(w2000) );
	vdp_not g1848 (.nZ(HPOS[3]), .A(w2001) );
	vdp_not g1849 (.nZ(VPOS[3]), .A(w1737) );
	vdp_not g1850 (.nZ(HPOS[2]), .A(w1773) );
	vdp_not g1851 (.nZ(VPOS[2]), .A(w1725) );
	vdp_not g1852 (.nZ(HPOS[1]), .A(w1724) );
	vdp_not g1853 (.nZ(VPOS[1]), .A(w1683) );
	vdp_not g1854 (.nZ(HPOS[0]), .A(w1684) );
	vdp_not g1855 (.nZ(VPOS[0]), .A(w1677) );
	vdp_aoi22 g1856 (.Z(w1956), .A1(w1698), .B1(w1700), .B2(w1709), .A2(w1699) );
	vdp_aon22 g1857 (.Z(w1726), .A2(w1699), .B1(w1728), .B2(w1709), .A1(w1769) );
	vdp_aoi22 g1858 (.Z(w1677), .B2(w1774), .B1(w1707), .A1(ODD/EVEN), .A2(w1) );
	vdp_aoi22 g1859 (.Z(w1683), .B2(w1774), .B1(w1850), .A1(w1707), .A2(w1) );
	vdp_aoi22 g1860 (.Z(w1725), .A2(w1), .A1(w1850), .B2(w1774), .B1(w1948) );
	vdp_aoi22 g1861 (.Z(w1737), .A1(w1948), .B2(w1774), .A2(w1), .B1(w1835) );
	vdp_aoi22 g1862 (.Z(w2000), .B1(w1947), .A1(w1835), .A2(w1), .B2(w1774) );
	vdp_aoi22 g1863 (.Z(w1999), .B1(w1791), .A1(w1947), .A2(w1), .B2(w1774) );
	vdp_aoi22 g1864 (.Z(w1998), .A2(w1), .B2(w1774), .B1(w1754), .A1(w1791) );
	vdp_aoi22 g1865 (.Z(w1753), .B2(w1774), .A1(w1754), .B1(w1824), .A2(w1) );
	vdp_aoi22 g1866 (.Z(w1962), .B2(w1774), .A2(w1), .A1(w1824), .B1(w1851) );
	vdp_aoi22 g1867 (.Z(w1963), .B1(1'b0), .A2(w1), .B2(w1774), .A1(w1851) );
	vdp_comp_ g1868 (.Q(w1656), .D(w1702), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_comp_ g1869 (.Q(w1807), .D(w1986), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_cnt_bit g1870 (.CI(w1988), .Q(w1866), .nEN(SYSRES), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g1871 (.nZ(w1959), .A(w55) );
	vdp_and g1872 (.Z(w1794), .A(w1809), .B(w1745) );
	vdp_and g1873 (.Z(w1795), .A(w1809), .B(w1745) );
	vdp_and g1874 (.Z(w1797), .A(w2013), .B(w1798) );
	vdp_and g1875 (.Z(w1798), .A(w1798), .B(w1811) );
	vdp_and g1876 (.Z(w1796), .A(w1855), .B(w1762) );
	vdp_and g1877 (.Z(w2013), .A(w1854), .B(w1743) );
	vdp_and g1878 (.Z(w1736), .A(w53), .B(w1722) );
	vdp_and g1879 (.Z(w16), .A(w1980), .B(w1713) );
	vdp_and g1880 (.Z(w1720), .A(w1682), .B(w1722) );
	vdp_and g1881 (.Z(w26), .A(w1641), .B(w1943) );
	vdp_and g1882 (.Z(w1721), .A(w52), .B(w1807) );
	vdp_and g1883 (.Z(w1747), .A(w1940), .B(w53) );
	vdp_and g1884 (.Z(w15), .A(w1713), .B(w1804) );
	vdp_and g1885 (.Z(w1779), .A(w2002), .B(w1747) );
	vdp_and g1886 (.Z(w10), .A(w1865), .B(w1713) );
	vdp_and g1887 (.Z(w1973), .A(w1815), .B(w4) );
	vdp_or g1888 (.Z(w1820), .A(w1946), .B(w1949) );
	vdp_or g1889 (.Z(w1819), .A(w1976), .B(w1949) );
	vdp_and g1890 (.Z(w1781), .A(M5), .B(w23) );
	vdp_and g1891 (.Z(w1988), .A(w1816), .B(w1769) );
	vdp_or g1892 (.Z(w1803), .A(SYSRES), .B(w1802) );
	vdp_or g1893 (.Z(w28), .A(w1788), .B(w1787) );
	vdp_or g1894 (.Z(w24), .A(w1782), .B(w1788) );
	vdp_or g1895 (.Z(w2010), .A(w1794), .B(w1798) );
	vdp_or g1896 (.Z(w1812), .A(w1800), .B(w1759) );
	vdp_or g1897 (.Z(w1945), .A(SYSRES), .B(w1802) );
	vdp_or g1898 (.Z(w1802), .A(w1748), .B(w1813) );
	vdp_or g1899 (.Z(w1985), .A(w1760), .B(SYSRES) );
	vdp_or g1900 (.Z(w1970), .A(w1681), .B(w2012) );
	vdp_or g1901 (.Z(w1944), .A(SYSRES), .B(w1759) );
	vdp_or g1902 (.Z(w1983), .A(w1721), .B(w1656) );
	vdp_or g1903 (.Z(w1931), .A(w1984), .B(w1805) );
	vdp_and g1904 (.Z(w11), .A(w1763), .B(w1713) );
	vdp_and g1905 (.Z(w1805), .A(w1671), .B(w1747) );
	vdp_or g1906 (.Z(w2008), .A(SYSRES), .B(w1748) );
	vdp_not g1907 (.nZ(w1697), .A(w54) );
	vdp_not g1908 (.nZ(w1696), .A(w48) );
	vdp_aon33 g1909 (.Z(w1847), .A3(w1846), .A2(w1959), .A1(w4), .B1(w55), .B3(1'b1), .B2(w1245) );
	vdp_aoi21 g1910 (.Z(w1957), .A1(w1703), .A2(w1713), .B(w1672) );
	vdp_aoi21 g1911 (.Z(w1712), .A1(w1710), .B(w1711), .A2(w1713) );
	vdp_aoi21 g1912 (.Z(w1673), .A1(w40), .A2(w50), .B(w1706) );
	vdp_aoi21 g1913 (.Z(w1739), .A1(w1719), .B(w1981), .A2(w1983) );
	vdp_aoi21 g1914 (.Z(w1978), .A1(w1713), .B(w1977), .A2(w1714) );
	vdp_aoi21 g1915 (.Z(w1771), .B(w1987), .A1(w1713), .A2(w1734) );
	vdp_aoi21 g1916 (.Z(w1958), .A1(w1713), .A2(w1785), .B(w1786) );
	vdp_xor g1917 (.Z(w1769), .B(w1670), .A(w1746) );
	vdp_xor g1918 (.Z(w1817), .A(ODD/EVEN), .B(w1843) );
	vdp_and3 g1919 (.Z(w1672), .A(w1733), .B(w42), .C(w1679) );
	vdp_and3 g1920 (.Z(w2017), .A(w2016), .B(w1870), .C(w1730) );
	vdp_and3 g1921 (.Z(w1711), .A(w1715), .B(w51), .C(w1679) );
	vdp_and3 g1922 (.Z(w1977), .A(w51), .B(w1679), .C(w42) );
	vdp_and3 g1923 (.Z(w1987), .A(w1715), .B(w1733), .C(w1788) );
	vdp_and3 g1924 (.Z(w1786), .A(w42), .B(w1733), .C(w41) );
	vdp_or3 g1925 (.Z(w2009), .A(w1796), .B(w1797), .C(w1795) );
	vdp_and3 g1926 (.Z(w2012), .A(w53), .B(w1722), .C(M5) );
	vdp_and3 g1927 (.Z(w1881), .A(w1719), .B(w53), .C(w1705) );
	vdp_and3 g1928 (.Z(w1681), .A(H40), .B(M5), .C(w1682) );
	vdp_nor4 g1929 (.Z(w1730), .A(w1772), .B(w1808), .C(w1675), .D(w1770) );
	vdp_nor4 g1930 (.Z(w1846), .A(w56), .B(w1849), .D(w1973), .C(SYSRES) );
	vdp_comp_we g1931 (.Z(w1830), .nZ(w1972), .A(w1848) );
	vdp_comp_we g1932 (.Z(w1832), .nZ(w1833), .A(w56) );
	vdp_comp_we g1933 (.Z(w1954), .nZ(w1680), .A(w57) );
	vdp_comp_we g1934 (.Z(w1687), .nZ(w1686), .A(w1671) );
	vdp_and3 g1935 (.Z(w18), .A(w1119), .B(w1943), .C(w31) );
	vdp_or4 g1936 (.Z(w1671), .A(w57), .B(SYSRES), .C(w1881), .D(w2003) );
	vdp_nor3 g1937 (.Z(w1870), .A(w1873), .B(w1731), .C(w1880) );
	vdp_nor3 g1938 (.Z(w1809), .A(w1743), .B(w1855), .C(w1854) );
	vdp_nand g1939 (.Z(w1764), .A(w1765), .B(w1806) );
	vdp_nand g1940 (.Z(w2018), .A(w1726), .B(w2014) );
	vdp_nand g1941 (.Z(w1874), .A(w1979), .B(w1731) );
	vdp_nor3 g1942 (.Z(w1713), .A(w42), .B(w51), .C(w41) );
	vdp_nor g1943 (.Z(w1949), .A(w1843), .B(M5) );
	vdp_nor g1944 (.Z(w1818), .A(ODD/EVEN), .B(w1843) );
	vdp_nor g1945 (.Z(w1946), .A(w1831), .B(w1205) );
	vdp_nor g1946 (.Z(w1976), .A(w1831), .B(w1843) );
	vdp_nor g1947 (.Z(w1981), .A(w1655), .B(SYSRES) );
	vdp_SDELAY8 g1948 (.Q(w1821), .D(w1799), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2), .nC3(nHCLK1), .C3(HCLK1), .nC4(nHCLK2), .C4(HCLK2), .nC5(nHCLK1), .C5(HCLK1), .nC6(nHCLK2), .C6(HCLK2), .nC7(nHCLK1), .C7(HCLK1), .nC8(nHCLK2), .C8(HCLK2), .nC9(nHCLK1), .C9(HCLK1), .nC10(nHCLK2), .C10(HCLK2), .nC11(nHCLK1), .C11(HCLK1), .nC12(nHCLK2), .C12(HCLK2), .nC13(nHCLK1), .C13(HCLK1), .nC14(nHCLK2), .C14(HCLK2), .nC15(nHCLK1), .C15(HCLK1), .nC16(nHCLK2), .C16(HCLK2) );
	vdp_SDELAY7 g1949 (.Q(w1766), .D(w1767), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .nC4(nHCLK2), .C5(HCLK1), .nC5(nHCLK1), .C6(HCLK2), .nC6(nHCLK2), .C7(HCLK1), .nC7(nHCLK1), .C8(HCLK2), .nC8(nHCLK2), .C9(HCLK1), .nC9(nHCLK1), .C10(HCLK2), .nC10(nHCLK2), .C11(HCLK1), .nC11(nHCLK1), .C12(HCLK2), .nC12(nHCLK2), .C13(HCLK1), .nC13(nHCLK1), .C14(HCLK2), .nC14(nHCLK2), .C3(HCLK1) );
	vdp_SDELAY8 g1950 (.Q(w1728), .D(w1769), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2), .C3(HCLK1), .nC4(nHCLK2), .C4(HCLK2), .nC5(nHCLK1), .C5(HCLK1), .nC6(nHCLK2), .C6(HCLK2), .nC7(nHCLK1), .C7(HCLK1), .nC8(nHCLK2), .C8(HCLK2), .nC9(nHCLK1), .C9(HCLK1), .nC10(nHCLK2), .C10(HCLK2), .C11(HCLK1), .nC12(nHCLK2), .C12(HCLK2), .nC13(nHCLK1), .C13(HCLK1), .nC14(nHCLK2), .C14(HCLK2), .nC15(nHCLK1), .C15(HCLK1), .nC16(nHCLK2), .C16(HCLK2), .nC3(nHCLK1), .nC11(nHCLK1) );
	vdp_SDELAY8 g1951 (.Q(w1700), .D(w1698), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2), .C3(HCLK1), .nC4(nHCLK2), .C4(HCLK2), .nC5(nHCLK1), .C5(HCLK1), .nC6(nHCLK2), .C6(HCLK2), .nC7(nHCLK1), .C7(HCLK1), .nC8(nHCLK2), .C8(HCLK2), .nC9(nHCLK1), .C9(HCLK1), .nC10(nHCLK2), .C10(HCLK2), .nC11(nHCLK1), .C11(HCLK1), .nC12(nHCLK2), .C12(HCLK2), .nC13(nHCLK1), .C13(HCLK1), .nC14(nHCLK2), .C14(HCLK2), .nC15(nHCLK1), .C15(HCLK1), .nC16(nHCLK2), .C16(HCLK2), .nC3(nHCLK1) );
	vdp_cnt_bit_load g1952 (.D(w1841), .Q(w1850), .nL(w1972), .L(w1830), .CI(w1939), .nC1(nHCLK1), .CO(w2020), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1953 (.D(w1840), .Q(w1948), .nL(w1972), .L(w1830), .CI(w2020), .nC1(nHCLK1), .CO(w2021), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1954 (.D(w1974), .Q(w1835), .nL(w1972), .L(w1830), .CI(w2021), .nC1(nHCLK1), .CO(w2022), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1955 (.D(w2023), .Q(w1947), .nL(w1972), .L(w1830), .CI(w2022), .nC1(nHCLK1), .CO(w1869), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1956 (.D(w1964), .Q(w1791), .nL(w1972), .L(w1830), .CI(w1869), .nC1(nHCLK1), .CO(w1868), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1957 (.D(w1965), .Q(w1754), .nL(w1972), .L(w1830), .CI(w1868), .nC1(nHCLK1), .CO(w2024), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1958 (.D(w1961), .Q(w1824), .nL(w1972), .L(w1830), .CI(w2024), .nC1(nHCLK1), .CO(w1867), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1959 (.D(w1960), .Q(w1851), .nL(w1972), .L(w1830), .CI(w1867), .nC1(nHCLK1), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1960 (.D(w1822), .Q(w1780), .nL(w1686), .L(w1687), .CI(w1823), .nC1(nHCLK1), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1961 (.D(w1966), .Q(w1752), .nL(w1686), .L(w1687), .CI(w1750), .nC1(nHCLK1), .CO(w1823), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1962 (.D(w1792), .Q(w1927), .nL(w1686), .L(w1687), .CI(w1790), .nC1(nHCLK1), .CO(w1750), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1963 (.D(w1967), .Q(w1775), .nL(w1686), .L(w1687), .CI(w1776), .nC1(nHCLK1), .CO(w1790), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1964 (.D(w2011), .Q(w1742), .nL(w1686), .L(w1687), .CI(w1741), .nC1(nHCLK1), .CO(w1776), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1965 (.D(w1968), .Q(w1694), .nL(w1686), .L(w1687), .CI(w1738), .nC1(nHCLK1), .CO(w1741), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1966 (.D(w1969), .Q(w1695), .nL(w1686), .L(w1687), .CI(w1723), .nC1(nHCLK1), .CO(w1738), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1967 (.D(w1995), .Q(w1690), .nL(w1686), .L(w1687), .CI(w2019), .nC1(nHCLK1), .CO(w1723), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1968 (.D(w1685), .Q(w1951), .nL(w1686), .L(w1687), .CI(w1872), .nC1(nHCLK1), .CO(w2019), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_or8 g1969 (.Z(w1836), .A(w1882), .B(w1883), .C(w1884), .D(w1885), .E(w1887), .F(w1937), .G(w1938), .H(w1887) );
	vdp_or8 g1970 (.Z(w1837), .A(w1888), .B(w1936), .C(w1935), .D(w1920), .E(w1889), .F(w1890), .G(w1891), .H(w1919) );
	vdp_or8 g1971 (.Z(w1838), .A(w1914), .B(w2006), .C(w2007), .D(w1993), .E(w1918), .F(w1916), .G(w1992), .H(w1915) );
	vdp_or5 g1972 (.Z(w1839), .A(w1910), .B(w1911), .C(w1913), .D(w1912), .E(w2025) );
	vdp_or7 g1973 (.Z(w1828), .A(w1903), .B(w1904), .C(w1905), .D(w1906), .E(w1907), .F(w1908), .G(w1909) );
	vdp_or7 g1974 (.Z(w1826), .A(w1892), .B(w1893), .C(w1894), .D(w1895), .E(w1896), .F(w1897), .G(w1898) );
	vdp_nor g1975 (.Z(w1706), .A(w1671), .B(w40) );
	vdp_and g1976 (.Z(w17), .A(w1713), .B(w1732) );
	vdp_not g1977 (.nZ(w1654), .A(w1899) );
	vdp_nor3 g1978 (.Z(w1827), .A(w1902), .B(w1901), .C(w1900) );
	vdp_RS g1979 (.Q(w1635), .S(w1942), .R(w1637) );
	vdp_RS g1980 (.Q(w1633), .S(w1649), .R(w1645) );
	vdp_and g1981 (.Z(w1854), .A(w1624), .B(M5) );
	vdp_nor4 g1982 (.Z(w2016), .A(w1693), .B(w1692), .C(w1691), .D(w1689) );
	vdp_nand3 g1983 (.A(w2146), .B(w2145), .C(w2143), .Z(w2139) );
	vdp_nand3 g1984 (.A(w2143), .B(w2145), .C(w2148), .Z(w2134) );
	vdp_nand3 g1985 (.A(w2143), .B(w2146), .C(w2147), .Z(w2135) );
	vdp_nand3 g1986 (.A(w2147), .B(w2143), .C(w2148), .Z(w2136) );
	vdp_nand3 g1987 (.A(w2147), .B(w2144), .C(w2148), .Z(w2131) );
	vdp_nand3 g1988 (.A(w2144), .B(w2146), .C(w2147), .Z(w2130) );
	vdp_nand3 g1989 (.A(w2145), .B(w2144), .C(w2148), .Z(w2138) );
	vdp_nand3 g1990 (.A(w2146), .B(w2145), .C(w2144), .Z(w2137) );
	vdp_nand3 g1991 (.A(w2119), .B(w2120), .C(w2115), .Z(w2129) );
	vdp_nand3 g1992 (.A(w2115), .B(w2120), .C(w2118), .Z(w2128) );
	vdp_nand3 g1993 (.A(w2117), .B(w2116), .C(w2118), .Z(w2122) );
	vdp_nand3 g1994 (.A(w2116), .B(w2119), .C(w2117), .Z(w2123) );
	vdp_nand3 g1995 (.A(w2120), .B(w2116), .C(w2118), .Z(w2124) );
	vdp_nand3 g1996 (.A(w2119), .B(w2120), .C(w2116), .Z(w2125) );
	vdp_nand3 g1997 (.A(w2117), .B(w2115), .C(w2118), .Z(w2126) );
	vdp_nand3 g1998 (.A(w2115), .B(w2119), .C(w2117), .Z(w2127) );
	vdp_nand3 g1999 (.A(w2107), .B(w2105), .C(w2103), .Z(w2100) );
	vdp_nand3 g2000 (.A(w2103), .B(w2105), .C(w2108), .Z(w2099) );
	vdp_nand3 g2001 (.A(w2106), .B(w2104), .C(w2108), .Z(w2093) );
	vdp_nand3 g2002 (.A(w2104), .B(w2107), .C(w2106), .Z(w2094) );
	vdp_nand3 g2003 (.A(w2105), .B(w2104), .C(w2108), .Z(w2095) );
	vdp_nand3 g2004 (.A(w2107), .B(w2105), .C(w2104), .Z(w2096) );
	vdp_nand3 g2005 (.A(w2106), .B(w2103), .C(w2108), .Z(w2097) );
	vdp_nand3 g2006 (.A(w2103), .B(w2107), .C(w2106), .Z(w2098) );
	vdp_nand3 g2007 (.A(w2046), .B(w2043), .C(w2047), .Z(w2040) );
	vdp_nand3 g2008 (.A(w2047), .B(w2043), .C(w2045), .Z(w2039) );
	vdp_nand3 g2009 (.A(w2044), .B(w2042), .C(w2045), .Z(w2033) );
	vdp_nand3 g2010 (.A(w2042), .B(w2046), .C(w2044), .Z(w2034) );
	vdp_nand3 g2011 (.A(w2043), .B(w2042), .C(w2045), .Z(w2035) );
	vdp_nand3 g2012 (.A(w2046), .B(w2043), .C(w2042), .Z(w2036) );
	vdp_nand3 g2013 (.A(w2044), .B(w2047), .C(w2045), .Z(w2037) );
	vdp_nand3 g2014 (.A(w2047), .B(w2046), .C(w2044), .Z(w2038) );
	vdp_not g2015 (.nZ(w2041), .A(w2028) );
	vdp_not g2016 (.nZ(w2101), .A(w2027) );
	vdp_not g2017 (.nZ(w2109), .A(w2029) );
	vdp_not g2018 (.nZ(w2140), .A(w2026) );
	vdp_nand g2019 (.Z(w2031), .B(w2032), .A(w2041) );
	vdp_nand g2020 (.Z(w2032), .B(w2041), .A(w2048) );
	vdp_nand g2021 (.Z(w2091), .B(w2092), .A(w2101) );
	vdp_nand g2022 (.Z(w2092), .B(w2101), .A(w2052) );
	vdp_comp_we g2023 (.A(w2102), .Z(w2104), .nZ(w2103) );
	vdp_comp_we g2024 (.A(w2162), .Z(w2106), .nZ(w2105) );
	vdp_comp_we g2025 (.A(w2161), .Z(w2108), .nZ(w2107) );
	vdp_comp_we g2026 (.A(w2049), .Z(w2042), .nZ(w2047) );
	vdp_comp_we g2027 (.A(w2050), .Z(w2044), .nZ(w2043) );
	vdp_comp_we g2028 (.A(w2051), .Z(w2045), .nZ(w2046) );
	vdp_nand g2029 (.Z(w2110), .B(w2109), .A(w2113) );
	vdp_comp_we g2030 (.A(w2112), .Z(w2116), .nZ(w2115) );
	vdp_comp_we g2031 (.A(w2114), .Z(w2117), .nZ(w2120) );
	vdp_comp_we g2032 (.A(w2121), .Z(w2118), .nZ(w2119) );
	vdp_nand g2033 (.Z(w2111), .B(w2110), .A(w2109) );
	vdp_nand g2034 (.Z(w2132), .B(w2140), .A(w2141) );
	vdp_comp_we g2035 (.A(w2142), .Z(w2144), .nZ(w2143) );
	vdp_comp_we g2036 (.A(w2149), .Z(w2147), .nZ(w2145) );
	vdp_comp_we g2037 (.A(w2150), .Z(w2148), .nZ(w2146) );
	vdp_nand g2038 (.Z(w2133), .B(w2132), .A(w2140) );
	vdp_comp_str g2039 (.A(w2173), .Z(w2174), .nZ(w2172) );
	vdp_comp_str g2040 (.A(w2190), .Z(w2163), .nZ(w2164) );
	vdp_comp_str g2041 (.A(w2199), .Z(w2154), .nZ(w2153) );
	vdp_comp_str g2042 (.A(w2200), .Z(w2055), .nZ(w2054) );
	vdp_comp_str g2043 (.A(w2063), .Z(w2064), .nZ(w2065) );
	vdp_comp_str g2044 (.A(w2237), .Z(w2423), .nZ(w2300) );
	vdp_comp_str g2045 (.A(w2448), .Z(w2416), .nZ(w2415) );
	vdp_comp_str g2046 (.A(w2419), .Z(w2429), .nZ(w2417) );
	vdp_comp_str g2047 (.A(w2208), .Z(w2420), .nZ(w2418) );
	vdp_comp_str g2048 (.A(w2328), .Z(w2071), .nZ(w2075) );
	vdp_comp_str g2049 (.A(w2449), .Z(w2072), .nZ(w2076) );
	vdp_comp_str g2050 (.A(w2206), .Z(w2074), .nZ(w2077) );
	vdp_dlatch g2051 (.Q(w2433), .C(w2074), .D(w2201), .nC(w2077) );
	vdp_dlatch g2052 (.Q(w2432), .C(w2072), .D(w2201), .nC(w2076) );
	vdp_dlatch g2053 (.Q(w2395), .C(w2074), .D(w2335), .nC(w2077) );
	vdp_dlatch g2054 (.Q(w2431), .C(w2071), .D(w2201), .nC(w2075) );
	vdp_dlatch g2055 (.Q(w2436), .C(w2074), .D(w2336), .nC(w2077) );
	vdp_dlatch g2056 (.Q(w2394), .C(w2071), .D(w2335), .nC(w2075) );
	vdp_dlatch g2057 (.Q(w2396), .C(w2072), .D(w2335), .nC(w2076) );
	vdp_dlatch g2058 (.Q(w2330), .C(w2074), .D(w2338), .nC(w2077) );
	vdp_dlatch g2059 (.Q(w2434), .C(w2071), .D(w2336), .nC(w2075) );
	vdp_dlatch g2060 (.Q(w2435), .C(w2072), .D(w2336), .nC(w2076) );
	vdp_dlatch g2061 (.Q(w2084), .C(w2074), .D(w2073), .nC(w2077) );
	vdp_dlatch g2062 (.Q(w2329), .C(w2071), .D(w2338), .nC(w2075) );
	vdp_dlatch g2063 (.Q(w2331), .C(w2072), .D(w2338), .nC(w2076) );
	vdp_dlatch g2064 (.Q(w2081), .C(w2071), .D(w2073), .nC(w2075) );
	vdp_dlatch g2065 (.Q(w2083), .C(w2072), .D(w2073), .nC(w2076) );
	vdp_dlatch g2066 (.Q(w2078), .C(w2074), .D(w2070), .nC(w2077) );
	vdp_dlatch g2067 (.Q(w2090), .C(w2071), .D(w2070), .nC(w2075) );
	vdp_dlatch g2068 (.Q(w2079), .C(w2072), .D(w2070), .nC(w2076) );
	vdp_dlatch g2069 (.Q(w2409), .C(w2420), .D(w2201), .nC(w2418) );
	vdp_dlatch g2070 (.Q(w2408), .C(w2429), .D(w2201), .nC(w2417) );
	vdp_dlatch g2071 (.Q(w2414), .C(w2420), .D(w2335), .nC(w2418) );
	vdp_dlatch g2072 (.Q(w2410), .C(w2416), .D(w2201), .nC(w2415) );
	vdp_dlatch g2073 (.Q(w2402), .C(w2420), .D(w2336), .nC(w2418) );
	vdp_dlatch g2074 (.Q(w2412), .C(w2416), .D(w2335), .nC(w2415) );
	vdp_dlatch g2075 (.Q(w2413), .C(w2429), .D(w2335), .nC(w2417) );
	vdp_dlatch g2076 (.Q(w2399), .C(w2420), .D(w2338), .nC(w2418) );
	vdp_dlatch g2077 (.Q(w2400), .C(w2416), .D(w2336), .nC(w2415) );
	vdp_dlatch g2078 (.Q(w2401), .C(w2429), .D(w2336), .nC(w2417) );
	vdp_dlatch g2079 (.Q(w2397), .C(w2416), .D(w2338), .nC(w2415) );
	vdp_dlatch g2080 (.Q(w2398), .C(w2429), .D(w2338), .nC(w2417) );
	vdp_dlatch g2081 (.Q(w2284), .C(w2423), .D(w2336), .nC(w2300) );
	vdp_dlatch g2082 (.Q(w2426), .C(w2423), .D(w2335), .nC(w2300) );
	vdp_dlatch g2083 (.Q(w2427), .C(w2423), .D(w2201), .nC(w2300) );
	vdp_and g2084 (.Z(w2244), .A(w2427), .B(w2426) );
	vdp_and g2085 (.Z(w2411), .A(w2426), .B(w2424) );
	vdp_and g2086 (.Z(w2393), .A(w2427), .B(w2425) );
	vdp_and g2087 (.Z(w2339), .A(w2424), .B(w2425) );
	vdp_dlatch g2088 (.Q(w2176), .C(w2174), .D(w2170), .nC(w2172) );
	vdp_or g2089 (.Z(w2150), .A(w2175), .B(w2176) );
	vdp_notif0 g2090 (.A(w2150), .nZ(DB[0]), .nE(w2056) );
	vdp_dlatch g2091 (.Q(w2459), .C(w2174), .D(w2167), .nC(w2172) );
	vdp_or g2092 (.Z(w2149), .A(w2175), .B(w2459) );
	vdp_notif0 g2093 (.A(w2149), .nZ(DB[1]), .nE(w2056) );
	vdp_dlatch g2094 (.Q(w2460), .C(w2174), .D(w2169), .nC(w2172) );
	vdp_or g2095 (.Z(w2142), .A(w2175), .B(w2460) );
	vdp_notif0 g2096 (.A(w2142), .nZ(DB[2]), .nE(w2056) );
	vdp_dlatch g2097 (.Q(w2180), .C(w2174), .D(w2181), .nC(w2172) );
	vdp_or g2098 (.Z(w2141), .A(w2175), .B(w2180) );
	vdp_notif0 g2099 (.A(w2141), .nZ(w156), .nE(w2056) );
	vdp_dlatch g2100 (.Q(w2171), .C(w2163), .D(w2170), .nC(w2164) );
	vdp_or g2101 (.Z(w2121), .A(w2168), .B(w2171) );
	vdp_notif0 g2102 (.A(w2121), .nZ(DB[4]), .nE(w2056) );
	vdp_dlatch g2103 (.Q(w2166), .C(w2163), .D(w2167), .nC(w2164) );
	vdp_or g2104 (.Z(w2114), .A(w2168), .B(w2166) );
	vdp_notif0 g2105 (.A(w2114), .nZ(DB[5]), .nE(w2056) );
	vdp_dlatch g2106 (.Q(w2165), .C(w2163), .D(w2169), .nC(w2164) );
	vdp_or g2107 (.Z(w2112), .A(w2168), .B(w2165) );
	vdp_notif0 g2108 (.A(w2112), .nZ(DB[6]), .nE(w2056) );
	vdp_dlatch g2109 (.Q(w2160), .C(w2163), .D(w2181), .nC(w2164) );
	vdp_or g2110 (.Z(w2113), .A(w2168), .B(w2160) );
	vdp_notif0 g2111 (.A(w2113), .nZ(w160), .nE(w2056) );
	vdp_dlatch g2112 (.Q(w2458), .C(w2154), .D(w2461), .nC(w2153) );
	vdp_or g2113 (.Z(w2161), .A(w2155), .B(w2458) );
	vdp_notif0 g2114 (.A(w2161), .nZ(DB[8]), .nE(w2056) );
	vdp_dlatch g2115 (.Q(w2159), .C(w2154), .D(w2167), .nC(w2153) );
	vdp_or g2116 (.Z(w2162), .A(w2155), .B(w2159) );
	vdp_notif0 g2117 (.A(w2162), .nZ(DB[9]), .nE(w2056) );
	vdp_dlatch g2118 (.Q(w2152), .C(w2154), .D(w2169), .nC(w2153) );
	vdp_or g2119 (.Z(w2102), .A(w2155), .B(w2152) );
	vdp_notif0 g2120 (.A(w2102), .nZ(DB[10]), .nE(w2056) );
	vdp_dlatch g2121 (.Q(w2151), .C(w2154), .D(w2181), .nC(w2153) );
	vdp_or g2122 (.Z(w2052), .A(w2155), .B(w2151) );
	vdp_notif0 g2123 (.A(w2052), .nZ(w170), .nE(w2056) );
	vdp_dlatch g2124 (.Q(w2057), .C(w2055), .D(w2170), .nC(w2054) );
	vdp_or g2125 (.Z(w2051), .A(w2053), .B(w2057) );
	vdp_notif0 g2126 (.A(w2051), .nZ(DB[12]), .nE(w2056) );
	vdp_dlatch g2127 (.Q(w2058), .C(w2055), .D(w2167), .nC(w2054) );
	vdp_or g2128 (.Z(w2050), .A(w2053), .B(w2058) );
	vdp_notif0 g2129 (.A(w2050), .nZ(DB[13]), .nE(w2056) );
	vdp_dlatch g2130 (.Q(w2059), .C(w2055), .D(w2169), .nC(w2054) );
	vdp_or g2131 (.Z(w2049), .A(w2053), .B(w2059) );
	vdp_notif0 g2132 (.A(w2049), .nZ(DB[14]), .nE(w2056) );
	vdp_dlatch g2133 (.Q(w2060), .C(w2055), .D(w2181), .nC(w2054) );
	vdp_or g2134 (.Z(w2048), .A(w2053), .B(w2060) );
	vdp_notif0 g2135 (.A(w2048), .nZ(w358), .nE(w2056) );
	vdp_not g2136 (.A(w1152), .nZ(w2056) );
	vdp_not g2137 (.nZ(w2229), .A(w1061) );
	vdp_clkgen g2138 (.PH(w2229), .CLK1(w2230), .nCLK1(w2231), .CLK2(w2232), .nCLK2(w2233) );
	vdp_comp_dff g2139 (.D(SYSRES), .nC1(w2231), .C1(w2230), .C2(w2232), .nC2(w2233), .Q(w2261) );
	vdp_sr_bit g2140 (.D(w2261), .nC1(w2231), .nC2(w2233), .C1(w2230), .C2(w2232), .Q(w2263) );
	vdp_sr_bit g2141 (.D(w2236), .nC1(w2231), .nC2(w2233), .C1(w2230), .C2(w2232), .Q(w2235) );
	vdp_not g2142 (.nZ(w2262), .A(w2263) );
	vdp_and g2143 (.Z(w2234), .A(w2261), .B(w2262) );
	vdp_nor g2144 (.Z(w2236), .A(w2235), .B(w2234) );
	vdp_cnt_bit g2145 (.CI(w2235), .R(w2234), .C1(w2230), .nC1(w2231), .nC2(w2233), .C2(w2232), .Q(w2260) );
	vdp_dlatch_inv g2146 (.nQ(w2259), .D(w2260), .nC(w2231), .C(w2230) );
	vdp_not g2147 (.nZ(w2258), .A(w2259) );
	vdp_nand g2148 (.Z(w2257), .A(w2235), .B(w2259) );
	vdp_not g2149 (.nZ(w2256), .A(w2257) );
	vdp_not g2150 (.nZ(w2255), .A(w2254) );
	vdp_not g2151 (.nZ(w2212), .A(w2257) );
	vdp_not g2152 (.nZ(w2222), .A(w2256) );
	vdp_not g2153 (.nZ(w2221), .A(w2255) );
	vdp_not g2154 (.nZ(w2211), .A(w2254) );
	vdp_nand g2155 (.Z(w2254), .A(w2235), .B(w2258) );
	vdp_sr_bit g2156 (.D(w2364), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2220) );
	vdp_sr_bit g2157 (.D(w2365), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2364) );
	vdp_sr_bit g2158 (.D(w2363), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2365) );
	vdp_sr_bit g2159 (.D(w2224), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2363) );
	vdp_sr_bit g2160 (.D(w2362), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2223) );
	vdp_sr_bit g2161 (.D(w2361), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2362) );
	vdp_sr_bit g2162 (.D(w2360), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2361) );
	vdp_sr_bit g2163 (.D(w2228), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2360) );
	vdp_sr_bit g2164 (.D(w2359), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2227) );
	vdp_sr_bit g2165 (.D(w2358), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2359) );
	vdp_sr_bit g2166 (.D(w2357), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2358) );
	vdp_sr_bit g2167 (.D(w2290), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2357) );
	vdp_sr_bit g2168 (.D(w2355), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2289) );
	vdp_sr_bit g2169 (.D(w2356), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2355) );
	vdp_sr_bit g2170 (.D(w2354), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2356) );
	vdp_sr_bit g2171 (.D(w2288), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2354) );
	vdp_sr_bit g2172 (.D(w2353), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2287) );
	vdp_sr_bit g2173 (.D(w2352), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2353) );
	vdp_sr_bit g2174 (.D(w2351), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2352) );
	vdp_sr_bit g2175 (.D(w2276), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2351) );
	vdp_sr_bit g2176 (.D(w2350), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2275) );
	vdp_sr_bit g2177 (.D(w2349), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2350) );
	vdp_sr_bit g2178 (.D(w2346), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2349) );
	vdp_sr_bit g2179 (.D(w2273), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2346) );
	vdp_sr_bit g2180 (.D(w2347), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2274) );
	vdp_sr_bit g2181 (.D(w2348), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2347) );
	vdp_sr_bit g2182 (.D(w2374), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2348) );
	vdp_sr_bit g2183 (.D(w2342), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2374) );
	vdp_sr_bit g2184 (.D(w2373), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2343) );
	vdp_sr_bit g2185 (.D(w2375), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2373) );
	vdp_sr_bit g2186 (.D(w2376), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2375) );
	vdp_sr_bit g2187 (.D(w2311), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2376) );
	vdp_sr_bit g2188 (.D(w2301), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2310) );
	vdp_sr_bit g2189 (.D(w2302), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2301) );
	vdp_sr_bit g2190 (.D(w2303), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2302) );
	vdp_sr_bit g2191 (.D(w2312), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2303) );
	vdp_sr_bit g2192 (.D(w2218), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2308) );
	vdp_sr_bit g2193 (.D(w2217), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2218) );
	vdp_sr_bit g2194 (.D(w2216), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2217) );
	vdp_sr_bit g2195 (.D(w2214), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2216) );
	vdp_aon2222 g2196 (.Z(w2086), .D2(1'b0), .C2(w2090), .C1(w2082), .D1(w2089), .B1(w2079), .A2(w2078), .A1(w2080), .B2(w2088) );
	vdp_cgi2a g2197 (.Z(w2428), .A(w2086), .C(w2440), .B(w2220) );
	vdp_aon2222 g2198 (.Z(w2087), .D2(1'b0), .C2(w2081), .C1(w2082), .D1(w2089), .B1(w2083), .A2(w2084), .A1(w2080), .B2(w2088) );
	vdp_cgi2a g2199 (.Z(w2440), .A(w2087), .C(w2439), .B(w2223) );
	vdp_aon2222 g2200 (.Z(w2334), .D2(1'b0), .C2(w2329), .C1(w2082), .D1(w2089), .B1(w2331), .A2(w2330), .A1(w2080), .B2(w2088) );
	vdp_cgi2a g2201 (.Z(w2439), .A(w2334), .C(w2438), .B(w2227) );
	vdp_aon2222 g2202 (.Z(w2333), .D2(w2411), .C2(w2434), .C1(w2082), .D1(w2089), .B1(w2435), .A2(w2436), .A1(w2080), .B2(w2088) );
	vdp_cgi2a g2203 (.Z(w2438), .A(w2333), .C(w2340), .B(w2289) );
	vdp_aon2222 g2204 (.Z(w2332), .D2(w2393), .C2(w2394), .C1(w2082), .D1(w2089), .B1(w2396), .A2(w2395), .A1(w2080), .B2(w2088) );
	vdp_cgi2a g2205 (.Z(w2340), .A(w2332), .C(w2341), .B(w2287) );
	vdp_aon2222 g2206 (.Z(w2404), .D2(w2339), .C2(w2431), .C1(w2082), .D1(w2089), .B1(w2432), .A2(w2433), .A1(w2080), .B2(w2088) );
	vdp_cgi2a g2207 (.Z(w2341), .A(w2404), .C(w2437), .B(w2275) );
	vdp_aon2222 g2208 (.Z(w2403), .D2(1'b0), .C2(w2397), .C1(w2082), .D1(w2089), .B1(w2398), .A2(w2399), .A1(w2080), .B2(w2088) );
	vdp_cgi2a g2209 (.Z(w2437), .A(w2403), .C(w2430), .B(w2274) );
	vdp_aon2222 g2210 (.Z(w2405), .D2(1'b0), .C2(w2400), .C1(w2082), .D1(w2089), .B1(w2401), .A2(w2402), .A1(w2080), .B2(w2088) );
	vdp_cgi2a g2211 (.Z(w2430), .A(w2405), .C(w2304), .B(w2343) );
	vdp_aon2222 g2212 (.Z(w2406), .D2(1'b0), .C2(w2412), .C1(w2082), .D1(w2089), .B1(w2413), .A2(w2414), .A1(w2080), .B2(w2088) );
	vdp_cgi2a g2213 (.Z(w2304), .A(w2406), .C(w2305), .B(w2310) );
	vdp_aon2222 g2214 (.Z(w2307), .D2(1'b0), .C2(w2410), .C1(w2082), .D1(w2089), .B1(w2408), .A2(w2409), .A1(w2080), .B2(w2088) );
	vdp_cgi2a g2215 (.Z(w2305), .A(w2307), .C(1'b1), .B(w2308) );
	vdp_not g2216 (.nZ(w2089), .A(w2407) );
	vdp_sr_bit g2217 (.D(w2388), .C1(w2212), .C2(w2211), .nC1(w2222), .nC2(w2221), .Q(w2309) );
	vdp_nand g2218 (.Z(w2407), .A(w2383), .B(w2309) );
	vdp_not g2219 (.nZ(w2082), .A(w2389) );
	vdp_sr_bit g2220 (.D(w2384), .Q(w2388), .C1(w2212), .C2(w2211), .nC1(w2222), .nC2(w2221) );
	vdp_nand g2221 (.Z(w2389), .A(w2383), .B(w2388) );
	vdp_not g2222 (.nZ(w2088), .A(w2387) );
	vdp_sr_bit g2223 (.D(w2320), .Q(w2384), .C1(w2212), .C2(w2211), .nC1(w2222), .nC2(w2221) );
	vdp_nand g2224 (.Z(w2387), .A(w2383), .B(w2384) );
	vdp_not g2225 (.nZ(w2080), .A(w2385) );
	vdp_sr_bit g2226 (.D(w2386), .Q(w2320), .C1(w2212), .C2(w2211), .nC1(w2222), .nC2(w2221) );
	vdp_nand g2227 (.Z(w2385), .A(w2383), .B(w2320) );
	vdp_sr_bit g2228 (.D(w2210), .Q(w2291), .C1(w2212), .C2(w2211), .nC1(w2222), .nC2(w2221) );
	vdp_sr_bit g2229 (.D(w2392), .Q(w2390), .C1(w2212), .C2(w2211), .nC1(w2222), .nC2(w2221) );
	vdp_sr_bit g2230 (.D(w2391), .Q(w2392), .C1(w2212), .C2(w2211), .nC1(w2222), .nC2(w2221) );
	vdp_sr_bit g2231 (.D(w2319), .Q(w2391), .C1(w2212), .C2(w2211), .nC1(w2222), .nC2(w2221) );
	vdp_sr_bit g2232 (.D(w2428), .Q(w2319), .C1(w2212), .C2(w2211), .nC1(w2222), .nC2(w2221) );
	vdp_not g2233 (.nZ(w2383), .A(w2291) );
	vdp_nor4 g2234 (.Z(w2386), .A(w2388), .B(w2384), .D(w2320), .C(w2210) );
	vdp_nor4 g2235 (.Z(w2281), .A(w2323), .B(w2324), .D(w2321), .C(w2322) );
	vdp_nor4 g2236 (.Z(w2283), .A(w2316), .B(w2317), .D(w2296), .C(w2297) );
	vdp_nor3 g2237 (.Z(w2282), .A(w2292), .B(w2293), .C(w2294) );
	vdp_not g2238 (.nZ(w2068), .A(w2291) );
	vdp_nand4 g2239 (.Z(w2280), .A(w2281), .B(w2283), .D(w2251), .C(w2282) );
	vdp_nand g2240 (.Z(w2285), .A(w2219), .B(w2284) );
	vdp_nand g2241 (.Z(w2286), .A(w2280), .B(w2285) );
	vdp_lfsr_bit g2242 (.Q(w2316), .A(w2286), .C2(w2211), .C1(w2212), .nC2(w2221), .nC1(w2222), .C(w2314), .B(w2315) );
	vdp_lfsr_bit g2243 (.Q(w2317), .A(w2316), .C2(w2211), .C1(w2212), .nC2(w2221), .nC1(w2222), .C(w2314), .B(w2315) );
	vdp_lfsr_bit g2244 (.Q(w2297), .A(w2317), .C2(w2211), .C1(w2212), .nC2(w2221), .nC1(w2222), .C(w2314), .B(w2315) );
	vdp_lfsr_bit g2245 (.Q(w2296), .A(w2297), .C2(w2211), .C1(w2212), .nC2(w2221), .nC1(w2222), .C(w2314), .B(w2315) );
	vdp_lfsr_bit g2246 (.Q(w2292), .A(w2296), .C2(w2211), .C1(w2212), .nC2(w2221), .nC1(w2222), .C(w2314), .B(w2315) );
	vdp_lfsr_bit g2247 (.Q(w2293), .A(w2292), .C2(w2211), .C1(w2212), .nC2(w2221), .nC1(w2222), .C(w2314), .B(w2315) );
	vdp_lfsr_bit g2248 (.Q(w2294), .A(w2293), .C2(w2211), .C1(w2212), .nC2(w2221), .nC1(w2222), .C(w2314), .B(w2315) );
	vdp_lfsr_bit g2249 (.Q(w2321), .A(w2294), .C2(w2211), .C1(w2212), .nC2(w2221), .nC1(w2222), .C(w2314), .B(w2315) );
	vdp_lfsr_bit g2250 (.Q(w2322), .A(w2321), .C2(w2211), .C1(w2212), .nC2(w2221), .nC1(w2222), .C(w2314), .B(w2315) );
	vdp_lfsr_bit g2251 (.Q(w2323), .A(w2322), .C2(w2211), .C1(w2212), .nC2(w2221), .nC1(w2222), .C(w2314), .B(w2315) );
	vdp_lfsr_bit g2252 (.Q(w2324), .A(w2323), .C2(w2211), .C1(w2212), .nC2(w2221), .nC1(w2222), .C(w2314), .B(w2315) );
	vdp_lfsr_bit g2253 (.Q(w2325), .A(w2324), .C2(w2211), .C1(w2212), .nC2(w2221), .nC1(w2222), .C(w2314), .B(w2315) );
	vdp_lfsr_bit g2254 (.Q(w2326), .A(w2325), .C2(w2211), .C1(w2212), .nC2(w2221), .nC1(w2222), .C(w2314), .B(w2315) );
	vdp_lfsr_bit g2255 (.Q(w2313), .A(w2326), .C2(w2212), .C1(w2212), .nC2(w2221), .nC1(w2222), .C(w2314), .B(w2315) );
	vdp_lfsr_bit g2256 (.Q(w2213), .A(w2313), .C2(w2211), .C1(w2212), .nC2(w2221), .nC1(w2222), .C(w2314), .B(w2315) );
	vdp_lfsr_bit g2257 (.Q(w2327), .A(w2213), .C2(w2211), .C1(w2212), .nC2(w2221), .nC1(w2222), .C(w2314), .B(w2315) );
	vdp_xor g2258 (.Z(w2219), .A(w2326), .B(w2327) );
	vdp_and g2259 (.Z(w2372), .A(w2215), .B(w2308) );
	vdp_ha g2260 (.SUM(w2214), .CO(w2270), .B(w2372), .A(1'b1) );
	vdp_and g2261 (.Z(w2345), .A(w2215), .B(w2310) );
	vdp_ha g2262 (.SUM(w2312), .CO(w2269), .B(w2345), .A(w2270) );
	vdp_and g2263 (.Z(w2344), .A(w2215), .B(w2343) );
	vdp_ha g2264 (.SUM(w2311), .CO(w2268), .B(w2344), .A(w2269) );
	vdp_and g2265 (.Z(w2272), .A(w2215), .B(w2274) );
	vdp_ha g2266 (.SUM(w2342), .CO(w2267), .B(w2272), .A(w2268) );
	vdp_and g2267 (.Z(w2371), .A(w2215), .B(w2275) );
	vdp_ha g2268 (.SUM(w2273), .CO(w2266), .B(w2371), .A(w2267) );
	vdp_and g2269 (.Z(w2370), .A(w2215), .B(w2287) );
	vdp_ha g2270 (.SUM(w2276), .CO(w2265), .B(w2370), .A(w2266) );
	vdp_and g2271 (.Z(w2369), .A(w2215), .B(w2289) );
	vdp_ha g2272 (.SUM(w2288), .CO(w2264), .B(w2369), .A(w2265) );
	vdp_and g2273 (.Z(w2368), .A(w2215), .B(w2227) );
	vdp_ha g2274 (.SUM(w2290), .CO(w2226), .B(w2368), .A(w2264) );
	vdp_and g2275 (.Z(w2367), .A(w2215), .B(w2223) );
	vdp_ha g2276 (.SUM(w2228), .CO(w2225), .B(w2367), .A(w2226) );
	vdp_and g2277 (.Z(w2366), .A(w2215), .B(w2220) );
	vdp_ha g2278 (.SUM(w2224), .B(w2366), .A(w2225) );
	vdp_and g2279 (.Z(w2295), .A(w2320), .B(w2390) );
	vdp_cnt_bit g2280 (.CI(w2295), .R(w2291), .C1(w2212), .nC1(w2222), .nC2(w2221), .C2(w2211), .Q(w2421) );
	vdp_and g2281 (.Z(w2299), .A(w2320), .B(w2392) );
	vdp_cnt_bit g2282 (.CI(w2299), .R(w2291), .C1(w2212), .nC1(w2222), .nC2(w2221), .C2(w2211), .Q(w2422) );
	vdp_and g2283 (.Z(w2298), .A(w2320), .B(w2391) );
	vdp_cnt_bit g2284 (.CI(w2298), .R(w2291), .C1(w2212), .nC1(w2222), .nC2(w2221), .C2(w2211), .Q(w2245) );
	vdp_and g2285 (.Z(w2318), .A(w2320), .B(w2319) );
	vdp_cnt_bit g2286 (.CI(w2318), .R(w2291), .C1(w2212), .nC1(w2222), .nC2(w2221), .C2(w2211), .Q(w2238) );
	vdp_nor g2287 (.Z(w2215), .A(w2428), .B(w2291) );
	vdp_dlatch g2288 (.Q(w2069), .C(w2066), .D(w160), .nC(w2067) );
	vdp_comp_str g2289 (.A(w1068), .Z(w2066), .nZ(w2067) );
	vdp_and g2290 (.Z(w2061), .A(w2068), .B(w2069) );
	vdp_and g2291 (.Z(w2063), .A(w2062), .B(w2061) );
	vdp_and g2292 (.Z(w2447), .A(w2068), .B(w2446) );
	vdp_dlatch g2293 (.Q(w2446), .C(w2066), .D(DB[6]), .nC(w2067) );
	vdp_dlatch g2294 (.Q(w2189), .C(w2064), .D(w2447), .nC(w2065) );
	vdp_and g2295 (.Z(w2070), .A(w2068), .B(w2157) );
	vdp_dlatch g2296 (.Q(w2157), .C(w2066), .D(DB[5]), .nC(w2067) );
	vdp_dlatch g2297 (.Q(w2158), .C(w2064), .D(w2070), .nC(w2065) );
	vdp_and g2298 (.Z(w2073), .A(w2068), .B(w2156) );
	vdp_dlatch g2299 (.Q(w2156), .C(w2066), .D(DB[4]), .nC(w2067) );
	vdp_dlatch g2300 (.Q(w2188), .C(w2064), .D(w2073), .nC(w2065) );
	vdp_and g2301 (.Z(w2338), .A(w2068), .B(w2195) );
	vdp_dlatch g2302 (.Q(w2195), .C(w2066), .D(w156), .nC(w2067) );
	vdp_or g2303 (.Z(w2181), .A(w2196), .B(w2338) );
	vdp_and g2304 (.Z(w2336), .A(w2068), .B(w2445) );
	vdp_or g2305 (.Z(w2169), .A(w2196), .B(w2336) );
	vdp_dlatch g2306 (.Q(w2445), .C(w2066), .D(DB[2]), .nC(w2067) );
	vdp_not g2307 (.nZ(w2196), .A(w2068) );
	vdp_and g2308 (.Z(w2335), .A(w2068), .B(w2337) );
	vdp_or g2309 (.Z(w2167), .A(w2196), .B(w2335) );
	vdp_dlatch g2310 (.Q(w2337), .C(w2066), .D(DB[1]), .nC(w2067) );
	vdp_and g2311 (.Z(w2201), .A(w2068), .B(w2202) );
	vdp_or g2312 (.Z(w2461), .A(w2196), .B(w2201) );
	vdp_dlatch g2313 (.Q(w2202), .C(w2066), .D(DB[0]), .nC(w2067) );
	vdp_not g2314 (.nZ(w2200), .A(w2198) );
	vdp_aoi21 g2315 (.Z(w2198), .B(w2210), .A1(w2203), .A2(w2197) );
	vdp_and3 g2316 (.Z(w2197), .A(w2178), .B(w2177), .C(w2188) );
	vdp_not g2317 (.nZ(w2199), .A(w2443) );
	vdp_aoi21 g2318 (.Z(w2443), .B(w2210), .A1(w2203), .A2(w2444) );
	vdp_and3 g2319 (.Z(w2444), .A(w2178), .B(w2158), .C(w2188) );
	vdp_not g2320 (.nZ(w2462), .A(w2442) );
	vdp_aoi21 g2321 (.Z(w2442), .B(w2210), .A1(w2203), .A2(w2441) );
	vdp_and3 g2322 (.Z(w2441), .A(w2189), .B(w2177), .C(w2179) );
	vdp_not g2323 (.nZ(w2207), .A(w2061) );
	vdp_or g2324 (.Z(w2209), .A(w2061), .B(w2210) );
	vdp_and g2325 (.Z(w2448), .A(w2209), .B(w2462) );
	vdp_and g2326 (.Z(w2328), .A(w2207), .B(w2462) );
	vdp_and g2327 (.Z(w2419), .A(w2209), .B(w2194) );
	vdp_and g2328 (.Z(w2449), .A(w2207), .B(w2194) );
	vdp_not g2329 (.nZ(w2194), .A(w2193) );
	vdp_aoi21 g2330 (.Z(w2193), .B(w2210), .A1(w2203), .A2(w2192) );
	vdp_and3 g2331 (.Z(w2192), .A(w2178), .B(w2158), .C(w2179) );
	vdp_not g2332 (.nZ(w2190), .A(w2191) );
	vdp_aoi21 g2333 (.Z(w2191), .B(w2210), .A1(w2203), .A2(w2205) );
	vdp_and3 g2334 (.Z(w2205), .A(w2189), .B(w2177), .C(w2188) );
	vdp_and g2335 (.Z(w2208), .A(w2209), .B(w2204) );
	vdp_and g2336 (.Z(w2206), .A(w2207), .B(w2204) );
	vdp_not g2337 (.nZ(w2204), .A(w2187) );
	vdp_aoi21 g2338 (.Z(w2187), .B(w2210), .A1(w2203), .A2(w2186) );
	vdp_and3 g2339 (.Z(w2186), .A(w2178), .B(w2177), .C(w2179) );
	vdp_and3 g2340 (.Z(w2185), .A(w2189), .B(w2158), .C(w2188) );
	vdp_not g2341 (.nZ(w2173), .A(w2184) );
	vdp_aoi21 g2342 (.Z(w2184), .B(w2210), .A1(w2203), .A2(w2185) );
	vdp_and3 g2343 (.Z(w2182), .A(w2189), .B(w2158), .C(w2179) );
	vdp_not g2344 (.nZ(w2237), .A(w2183) );
	vdp_aoi21 g2345 (.Z(w2183), .B(w2210), .A1(w2203), .A2(w2182) );
	vdp_not g2346 (.nZ(w2424), .A(w2427) );
	vdp_not g2347 (.nZ(w2425), .A(w2426) );
	vdp_not g2348 (.nZ(w2179), .A(w2188) );
	vdp_not g2349 (.nZ(w2177), .A(w2158) );
	vdp_not g2350 (.nZ(w2178), .A(w2189) );
	vdp_nor g2351 (.Z(w2053), .A(w2421), .B(w1165) );
	vdp_nor g2352 (.Z(w2155), .A(w2422), .B(w1165) );
	vdp_nor g2353 (.Z(w2168), .A(w2245), .B(w1165) );
	vdp_nor g2354 (.Z(w2175), .A(w2213), .B(w1165) );
	vdp_aon22 g2355 (.Z(w2240), .A2(w2245), .A1(w2244), .B2(w2239), .B1(w2238) );
	vdp_sr_bit g2356 (.D(w2240), .nC1(w2222), .nC2(w2221), .C1(w2212), .C2(w2211), .Q(w2241) );
	vdp_not g2357 (.nZ(w2239), .A(w2244) );
	vdp_not g2358 (.nZ(w2242), .A(w2241) );
	vdp_not g2359 (.nZ(w2378), .A(w1166) );
	vdp_not g2360 (.nZ(w2377), .A(w1167) );
	vdp_not g2361 (.nZ(w2278), .A(w2277) );
	vdp_sr_bit g2362 (.D(w2062), .nC1(w2231), .nC2(w2233), .C1(w2230), .C2(w2232), .Q(w2203) );
	vdp_nand g2363 (.Z(w2379), .A(w1166), .B(w2377) );
	vdp_nand g2364 (.Z(w2243), .A(w1167), .B(w1166) );
	vdp_nand g2365 (.Z(w2380), .A(w2377), .B(w2378) );
	vdp_nand g2366 (.Z(w2381), .A(w1167), .B(w2378) );
	vdp_and g2367 (.Z(w2247), .A(w2240), .B(w2242) );
	vdp_and g2368 (.Z(w2026), .A(w1165), .B(w2243) );
	vdp_and g2369 (.Z(w2027), .A(w1165), .B(w2379) );
	vdp_and g2370 (.Z(w2028), .A(w1165), .B(w2380) );
	vdp_and g2371 (.Z(w2029), .A(w1165), .B(w2381) );
	vdp_nor4 g2372 (.Z(w2251), .A(w2313), .B(w2326), .D(w2325), .C(w2213) );
	vdp_not g2373 (.nZ(w2248), .A(w2247) );
	vdp_not g2374 (.nZ(w2315), .A(w2249) );
	vdp_not g2375 (.nZ(w2314), .A(w2382) );
	vdp_not g2376 (.nZ(w2210), .A(w2278) );
	vdp_nand g2377 (.Z(w2249), .A(w2246), .B(w2248) );
	vdp_nand g2378 (.Z(w2382), .A(w2246), .B(w2247) );
	vdp_nor g2379 (.Z(w2246), .A(w2210), .B(w2250) );
	vdp_rs_ff g2380 (.S(w2237), .R(w2250), .Q(w2279) );
	vdp_rs_ff g2381 (.S(w2062), .R(w1068), .Q(w2252) );
	vdp_nor g2382 (.Z(w2253), .A(w1068), .B(w2252) );
	vdp_comp_dff g2383 (.D(w2253), .nC1(w2231), .C1(w2230), .C2(w2232), .nC2(w2233), .Q(w2062) );
	vdp_comp_dff g2384 (.D(SYSRES), .nC1(w2222), .C1(w2212), .C2(w2211), .nC2(w2221), .Q(w2277) );
	vdp_comp_dff g2385 (.D(w2279), .nC1(w2222), .C1(w2212), .C2(w2211), .nC2(w2221), .Q(w2250) );
	vdp_sr_bit g2386 (.Q(w2639), .D(w2633), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2387 (.nZ(AD_RD_DIR), .A(w2632) );
	vdp_sr_bit g2388 (.Q(w2640), .D(w2498), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2389 (.Q(w2566), .D(w2511), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2390 (.Q(w2623), .D(w33), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2391 (.Q(w2490), .D(w35), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2392 (.nZ(w2635), .A(w2488) );
	vdp_or g2393 (.Z(w2498), .A(w35), .B(w2490) );
	vdp_sr_bit g2394 (.Q(w2507), .D(w2509), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_sr_bit g2395 (.Q(w2636), .D(w2625), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2396 (.nZ(w2565), .A(w2636) );
	vdp_or g2397 (.Z(w2486), .A(w2490), .B(w2489) );
	vdp_sr_bit g2398 (.Q(w2489), .D(w557), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2399 (.Q(w2487), .D(w32), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2400 (.Q(w2627), .D(w2487), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2401 (.Q(w2626), .D(w2499), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2402 (.Q(w2621), .D(w2623), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2403 (.Q(w2638), .D(w2643), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_not g2404 (.nZ(w2618), .A(w2698) );
	vdp_not g2405 (.nZ(w2510), .A(128k) );
	vdp_sr_bit g2406 (.Q(w2499), .D(VRAM_REFRESH), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2407 (.nZ(w2574), .A(w2485) );
	vdp_not g2408 (.nZ(w2641), .A(w2628) );
	vdp_not g2409 (.nZ(w2505), .A(w2497) );
	vdp_oai21 g2410 (.Z(w2485), .B(w2505), .A1(w2641), .A2(w2629) );
	vdp_or g2411 (.Z(w2497), .A(w2635), .B(w2634) );
	vdp_or g2412 (.Z(w2633), .A(w2489), .B(w557) );
	vdp_not g2413 (.nZ(w2642), .A(w2491) );
	vdp_not g2414 (.nZ(w2690), .A(w2643) );
	vdp_dlatch_inv g2415 (.nQ(w2643), .D(w3), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2416 (.nQ(w2637), .D(w2506), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g2417 (.nQ(w2506), .D(w2638), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g2418 (.nQ(w2488), .D(w2486), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2419 (.nQ(w2634), .D(w2488), .C(HCLK2), .nC(nHCLK2) );
	vdp_dlatch_inv g2420 (.nQ(w2631), .D(w2630), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2421 (.nQ(w2628), .D(w2627), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2422 (.nQ(w2629), .D(w2628), .C(HCLK2), .nC(nHCLK2) );
	vdp_aon22 g2423 (.Z(nCAS1), .A1(w2506), .B1(w2495), .B2(1'b1), .A2(w2636) );
	vdp_and3 g2424 (.Z(nWE1), .A(w2494), .B(w2640), .C(w2495) );
	vdp_and3 g2425 (.Z(nWE0), .A(w2495), .B(w2494), .C(w2639) );
	vdp_aoi222 g2426 (.Z(w2632), .A1(1'b1), .B1(w2492), .B2(1'b1), .A2(w100), .C1(w2497), .C2(w2495) );
	vdp_aon333 g2427 (.Z(nOE1), .A1(w2574), .A2(w2638), .A3(w2495), .B1(w2631), .B2(w2631), .B3(w2642), .C1(w2631), .C2(w2631), .C3(w2492) );
	vdp_or3 g2428 (.Z(w2630), .A(w2625), .B(w2627), .C(w2487) );
	vdp_sr_bit g2429 (.Q(w2492), .D(w2690), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_dlatch_inv g2430 (.nQ(w2494), .D(w2492), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g2431 (.nQ(w2624), .D(w2494), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g2432 (.nQ(w2495), .D(w2493), .C(DCLK1), .nC(nDCLK1) );
	vdp_not g2433 (.nZ(w2493), .A(w2624) );
	vdp_nand g2434 (.Z(w2721), .A(w2624), .B(w2492) );
	vdp_nand g2435 (.Z(w2720), .A(w2492), .B(w2637) );
	vdp_nand g2436 (.Z(w2501), .A(w2638), .B(1'b1) );
	vdp_aoi33 g2437 (.Z(w2704), .A1(w2621), .A2(w34), .A3(w34), .B1(w2512), .B2(w2513), .B3(w3) );
	vdp_and g2438 (.Z(w2508), .A(w2495), .B(w2494) );
	vdp_not g2439 (.nZ(w2502), .A(w2566) );
	vdp_comp_strong g2440 (.nZ(w2519), .Z(w2518), .A(w2525) );
	vdp_comp_strong g2441 (.nZ(w2590), .Z(w2613), .A(w2614) );
	vdp_comp_strong g2442 (.nZ(w2520), .Z(w2567), .A(w2614) );
	vdp_comp_strong g2443 (.nZ(w2572), .Z(w2571), .A(w2525) );
	vdp_comp_strong g2444 (.nZ(w2526), .Z(w2573), .A(w2522) );
	vdp_comp_strong g2445 (.nZ(w2577), .Z(w2619), .A(w2522) );
	vdp_g2446 g2446 (.nZ(w2528), .A(w2492) );
	vdp_g2447 g2447 (.nZ(w2513), .A(w34) );
	vdp_g2448 g2448 (.nZ(w2512), .A(w36) );
	vdp_comp_strong g2449 (.nZ(w2569), .Z(w2570), .A(w2508) );
	vdp_comp_strong g2450 (.nZ(w2503), .Z(w2615), .A(w2508) );
	vdp_or g2451 (.Z(w2625), .A(w2499), .B(w2626) );
	vdp_and g2452 (.Z(w2509), .A(128k), .B(HCLK1) );
	vdp_comp_we g2453 (.nZ(w2616), .Z(w2617), .A(w100) );
	vdp_comp_we g2454 (.nZ(w2521), .Z(w2702), .A(w2529) );
	vdp_not g2455 (.nZ(w2703), .A(w2566) );
	vdp_not g2456 (.nZ(w2524), .A(w2721) );
	vdp_not g2457 (.nZ(w2707), .A(w2720) );
	vdp_not g2458 (.nZ(w2706), .A(w2501) );
	vdp_comp_we g2459 (.nZ(w2554), .Z(w2553), .A(M5) );
	vdp_comp_we g2460 (.nZ(w2576), .Z(w2527), .A(128k) );
	vdp_and g2461 (.Z(w2511), .A(w110), .B(w3) );
	vdp_and g2462 (.Z(w2522), .A(w3), .B(HCLK1) );
	vdp_and g2463 (.Z(w2525), .A(HCLK2), .B(w2622) );
	vdp_and g2464 (.Z(w2614), .A(w3), .B(HCLK1) );
	vdp_oai21 g2465 (.Z(w2698), .A1(HCLK2), .A2(w2510), .B(DCLK1) );
	vdp_notif0 g2466 (.nZ(AD_DATA[0]), .A(w2516), .nE(w2502) );
	vdp_aon22 g2467 (.Z(nYS), .A1(VRAMA[16]), .A2(w2617), .B1(w2616), .B2(w2682) );
	vdp_aon22 g2468 (.Z(w2658), .A1(VRAMA[15]), .B1(w2719), .A2(w2617), .B2(w2597) );
	vdp_aon22 g2469 (.Z(w2656), .A1(VRAMA[14]), .B1(w2719), .A2(w2617), .B2(w2476) );
	vdp_aon22 g2470 (.Z(w2474), .A1(VRAMA[6]), .B1(w2616), .A2(w2617), .B2(w2657) );
	vdp_aon22 g2471 (.Z(w2466), .A1(VRAMA[7]), .B1(w2616), .A2(w2617), .B2(w2465) );
	vdp_aon22 g2472 (.Z(w2686), .A1(VRAMA[13]), .B1(w2719), .A2(w2617), .B2(w2484) );
	vdp_aon22 g2473 (.Z(w2655), .A1(VRAMA[5]), .B1(w2616), .A2(w2617), .B2(w2708) );
	vdp_aon22 g2474 (.Z(w2661), .A1(VRAMA[12]), .B1(w2616), .A2(w2617), .B2(w2556) );
	vdp_aon22 g2475 (.Z(w2482), .A1(VRAMA[4]), .B1(w2616), .A2(w2617), .B2(w2562) );
	vdp_aon22 g2476 (.Z(w2660), .A1(VRAMA[11]), .B1(w2616), .A2(w2617), .B2(w2713) );
	vdp_aon22 g2477 (.Z(w2596), .A1(VRAMA[3]), .B1(w2616), .A2(w2617), .B2(w2709) );
	vdp_aon22 g2478 (.Z(w2688), .A1(VRAMA[10]), .B1(w2616), .A2(w2617), .B2(w2609) );
	vdp_aon22 g2479 (.Z(w2595), .A1(VRAMA[2]), .B1(w2616), .A2(w2617), .B2(w2550) );
	vdp_aon22 g2480 (.Z(w2514), .A1(VRAMA[8]), .B1(w2616), .A2(w2617), .B2(w2517) );
	vdp_aon22 g2481 (.Z(w2711), .A1(VRAMA[0]), .B1(w2616), .A2(w2617), .B2(w2541) );
	vdp_aon22 g2482 (.Z(w2712), .A1(VRAMA[9]), .B1(w2616), .A2(w2617), .B2(w2591) );
	vdp_aon22 g2483 (.Z(w2544), .A1(VRAMA[1]), .B1(w2616), .A2(w2617), .B2(w2546) );
	vdp_notif0 g2484 (.nZ(AD_DATA[1]), .A(w2536), .nE(w2502) );
	vdp_notif0 g2485 (.nZ(AD_DATA[2]), .A(w2593), .nE(w2502) );
	vdp_notif0 g2486 (.nZ(AD_DATA[3]), .A(w2547), .nE(w2502) );
	vdp_notif0 g2487 (.nZ(AD_DATA[5]), .A(w2483), .nE(w2502) );
	vdp_notif0 g2488 (.nZ(AD_DATA[4]), .A(w2568), .nE(w2502) );
	vdp_notif0 g2489 (.nZ(AD_DATA[6]), .A(w2477), .nE(w2502) );
	vdp_notif0 g2490 (.nZ(AD_DATA[7]), .A(w2473), .nE(w2502) );
	vdp_slatch g2491 (.nQ(w2516), .D(w2515), .nC(w2503), .C(w2615) );
	vdp_slatch g2492 (.nQ(w2536), .D(w2535), .nC(w2503), .C(w2615) );
	vdp_slatch g2493 (.nQ(w2593), .D(w2543), .nC(w2503), .C(w2615) );
	vdp_slatch g2494 (.nQ(w2547), .D(w2548), .nC(w2503), .C(w2615) );
	vdp_slatch g2495 (.nQ(w2568), .D(w2500), .nC(w2503), .C(w2615) );
	vdp_slatch g2496 (.nQ(w2483), .D(w2687), .nC(w2503), .C(w2615) );
	vdp_slatch g2497 (.nQ(w2477), .D(w2475), .nC(w2503), .C(w2615) );
	vdp_slatch g2498 (.nQ(w2473), .D(w2659), .nC(w2503), .C(w2615) );
	vdp_slatch g2499 (.nQ(w2468), .D(w2467), .nC(w2569), .C(w2570) );
	vdp_slatch g2500 (.nQ(w2560), .D(w2557), .nC(w2569), .C(w2570) );
	vdp_slatch g2501 (.nQ(w2600), .D(w2699), .nC(w2569), .C(w2570) );
	vdp_slatch g2502 (.nQ(w2601), .D(w2481), .nC(w2569), .C(w2570) );
	vdp_slatch g2503 (.nQ(w2662), .D(w2558), .nC(w2569), .C(w2570) );
	vdp_slatch g2504 (.nQ(w2551), .D(w2549), .nC(w2569), .C(w2570) );
	vdp_slatch g2505 (.nQ(w2545), .D(w2594), .nC(w2569), .C(w2570) );
	vdp_slatch g2506 (.nQ(w2578), .D(w2689), .nC(w2569), .C(w2570) );
	vdp_slatch g2507 (.Q(w2517), .D(w2581), .nC(w2519), .C(w2518) );
	vdp_slatch g2508 (.Q(w2591), .D(w2715), .nC(w2519), .C(w2518) );
	vdp_slatch g2509 (.Q(w2713), .D(w2665), .nC(w2519), .C(w2518) );
	vdp_slatch g2510 (.Q(w2609), .D(w2592), .nC(w2519), .C(w2518) );
	vdp_slatch g2511 (.Q(w2484), .D(w2580), .nC(w2519), .C(w2518) );
	vdp_slatch g2512 (.Q(w2556), .D(w2666), .nC(w2519), .C(w2518) );
	vdp_slatch g2513 (.Q(w2597), .D(w2669), .nC(w2519), .C(w2518) );
	vdp_slatch g2514 (.Q(w2476), .D(w2579), .nC(w2519), .C(w2518) );
	vdp_slatch g2515 (.nQ(w2668), .D(w359), .nC(w2590), .C(w2613) );
	vdp_slatch g2516 (.nQ(w2670), .D(RD_DATA[6]), .nC(w2590), .C(w2613) );
	vdp_slatch g2517 (.nQ(w2667), .D(RD_DATA[5]), .nC(w2590), .C(w2613) );
	vdp_slatch g2518 (.nQ(w2717), .D(RD_DATA[4]), .nC(w2590), .C(w2613) );
	vdp_slatch g2519 (.nQ(w2664), .D(w324), .nC(w2590), .C(w2613) );
	vdp_slatch g2520 (.nQ(w2718), .D(RD_DATA[2]), .nC(w2590), .C(w2613) );
	vdp_slatch g2521 (.nQ(w2716), .D(RD_DATA[0]), .nC(w2590), .C(w2613) );
	vdp_slatch g2522 (.nQ(w2663), .D(RD_DATA[1]), .nC(w2590), .C(w2613) );
	vdp_notif0 g2523 (.nZ(w359), .A(w2468), .nE(w2703) );
	vdp_notif0 g2524 (.nZ(RD_DATA[6]), .A(w2560), .nE(w2703) );
	vdp_notif0 g2525 (.nZ(RD_DATA[5]), .A(w2600), .nE(w2703) );
	vdp_notif0 g2526 (.nZ(RD_DATA[4]), .A(w2601), .nE(w2703) );
	vdp_notif0 g2527 (.nZ(w324), .A(w2662), .nE(w2703) );
	vdp_notif0 g2528 (.nZ(RD_DATA[2]), .A(w2551), .nE(w2703) );
	vdp_notif0 g2529 (.nZ(RD_DATA[1]), .A(w2545), .nE(w2703) );
	vdp_notif0 g2530 (.nZ(RD_DATA[0]), .A(w2578), .nE(w2703) );
	vdp_slatch g2531 (.nQ(w2692), .D(AD_DATA[7]), .nC(w2520), .C(w2567) );
	vdp_slatch g2532 (.nQ(w2691), .D(AD_DATA[6]), .nC(w2520), .C(w2567) );
	vdp_slatch g2533 (.nQ(w2714), .D(AD_DATA[5]), .nC(w2520), .C(w2567) );
	vdp_slatch g2534 (.nQ(w2694), .D(AD_DATA[3]), .nC(w2520), .C(w2567) );
	vdp_slatch g2535 (.nQ(w2695), .D(AD_DATA[2]), .nC(w2520), .C(w2567) );
	vdp_slatch g2536 (.nQ(w2697), .D(AD_DATA[1]), .nC(w2520), .C(w2567) );
	vdp_slatch g2537 (.nQ(w2696), .D(AD_DATA[0]), .nC(w2520), .C(w2567) );
	vdp_slatch g2538 (.Q(w2472), .D(w2589), .nC(w2572), .C(w2571) );
	vdp_slatch g2539 (.Q(w2480), .D(w2588), .nC(w2572), .C(w2571) );
	vdp_slatch g2540 (.Q(w2559), .D(w2587), .nC(w2572), .C(w2571) );
	vdp_slatch g2541 (.Q(w2700), .D(w2584), .nC(w2572), .C(w2571) );
	vdp_slatch g2542 (.Q(w2612), .D(w2585), .nC(w2572), .C(w2571) );
	vdp_slatch g2543 (.Q(w2542), .D(w2583), .nC(w2572), .C(w2571) );
	vdp_slatch g2544 (.Q(w2599), .D(w2471), .nC(w2526), .C(w2573) );
	vdp_slatch g2545 (.Q(w2705), .D(w2479), .nC(w2526), .C(w2573) );
	vdp_slatch g2546 (.Q(w2672), .D(w2534), .nC(w2526), .C(w2573) );
	vdp_slatch g2547 (.Q(w2603), .D(w2533), .nC(w2526), .C(w2573) );
	vdp_slatch g2548 (.Q(w2610), .D(w2611), .nC(w2526), .C(w2573) );
	vdp_slatch g2549 (.Q(w2701), .D(w2539), .nC(w2526), .C(w2573) );
	vdp_slatch g2550 (.Q(w2608), .D(w2504), .nC(w2526), .C(w2573) );
	vdp_slatch g2551 (.Q(w2710), .D(w2540), .nC(w2526), .C(w2573) );
	vdp_slatch g2552 (.Q(w2620), .D(w2538), .nC(w2577), .C(w2619) );
	vdp_slatch g2553 (.Q(w2607), .D(w2726), .nC(w2577), .C(w2619) );
	vdp_slatch g2554 (.Q(w2552), .D(w2532), .nC(w2577), .C(w2619) );
	vdp_slatch g2555 (.Q(w2604), .D(w2722), .nC(w2577), .C(w2619) );
	vdp_slatch g2556 (.Q(w2563), .D(w2478), .nC(w2577), .C(w2619) );
	vdp_slatch g2557 (.Q(w2602), .D(w2530), .nC(w2577), .C(w2619) );
	vdp_slatch g2558 (.Q(w2561), .D(w2470), .nC(w2577), .C(w2619) );
	vdp_slatch g2559 (.Q(w2598), .D(w2469), .nC(w2577), .C(w2619) );
	vdp_sr_bit g2560 (.Q(w2529), .D(w34), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2561 (.nZ(w2733), .A(w111) );
	vdp_not g2562 (.nZ(w2605), .A(w2606) );
	vdp_not g2563 (.nZ(w2531), .A(M5) );
	vdp_not g2564 (.nZ(w2537), .A(w2528) );
	vdp_not g2565 (.nZ(w2491), .A(w2537) );
	vdp_aoi21 g2566 (.Z(w2606), .B(w2673), .A2(VRAMA[9]), .A1(w2531) );
	vdp_aoi22 g2567 (.Z(w2715), .A1(w2545), .B1(w2521), .B2(w2663), .A2(w2702) );
	vdp_aoi22 g2568 (.Z(w2665), .A1(w2662), .B1(w2521), .B2(w2664), .A2(w2702) );
	vdp_aoi22 g2569 (.Z(w2592), .A1(w2551), .B1(w2521), .B2(w2718), .A2(w2702) );
	vdp_aoi22 g2570 (.Z(w2580), .A1(w2600), .B1(w2521), .B2(w2667), .A2(w2702) );
	vdp_aoi22 g2571 (.Z(w2666), .A1(w2601), .B1(w2521), .B2(w2717), .A2(w2702) );
	vdp_aoi22 g2572 (.Z(w2669), .A1(w2468), .B1(w2521), .B2(w2668), .A2(w2702) );
	vdp_aoi22 g2573 (.Z(w2579), .A1(w2560), .B1(w2521), .B2(w2670), .A2(w2702) );
	vdp_slatch g2574 (.Q(w2523), .D(w2582), .nC(w2572), .C(w2571) );
	vdp_slatch g2575 (.nQ(w2693), .D(AD_DATA[4]), .nC(w2520), .C(w2567) );
	vdp_slatch g2576 (.Q(w2555), .D(w2586), .nC(w2572), .C(w2571) );
	vdp_aoi22 g2577 (.Z(w2582), .A1(w2516), .B1(w2521), .B2(w2696), .A2(w2702) );
	vdp_aoi22 g2578 (.Z(w2583), .A1(w2536), .B1(w2521), .B2(w2697), .A2(w2702) );
	vdp_aoi22 g2579 (.Z(w2584), .A1(w2593), .B1(w2521), .B2(w2695), .A2(w2702) );
	vdp_aoi22 g2580 (.Z(w2585), .A1(w2547), .B1(w2521), .B2(w2694), .A2(w2702) );
	vdp_aoi22 g2581 (.Z(w2586), .A1(w2568), .B1(w2521), .B2(w2693), .A2(w2702) );
	vdp_aoi22 g2582 (.Z(w2587), .A1(w2483), .B1(w2521), .B2(w2714), .A2(w2702) );
	vdp_aoi22 g2583 (.Z(w2589), .A1(w2473), .B1(w2521), .B2(w2692), .A2(w2702) );
	vdp_aoi22 g2584 (.Z(w2588), .A1(w2477), .B1(w2521), .B2(w2691), .A2(w2702) );
	vdp_aon22 g2585 (.Z(w2540), .A1(VRAMA[2]), .B1(w2554), .B2(VRAMA[1]), .A2(w2553) );
	vdp_aon22 g2586 (.Z(w2539), .A1(VRAMA[3]), .B1(w2554), .B2(VRAMA[2]), .A2(w2553) );
	vdp_aon22 g2587 (.Z(w2504), .A1(VRAMA[4]), .B1(w2554), .B2(VRAMA[3]), .A2(w2553) );
	vdp_aon22 g2588 (.Z(w2611), .A1(VRAMA[5]), .B1(w2554), .B2(VRAMA[4]), .A2(w2553) );
	vdp_aon22 g2589 (.Z(w2533), .A1(VRAMA[6]), .B1(w2554), .B2(VRAMA[5]), .A2(w2553) );
	vdp_aon22 g2590 (.Z(w2534), .A1(VRAMA[7]), .B1(w2554), .B2(VRAMA[6]), .A2(w2553) );
	vdp_aon22 g2591 (.Z(w2479), .A1(VRAMA[8]), .B1(w2554), .B2(VRAMA[7]), .A2(w2553) );
	vdp_aon22 g2592 (.Z(w2471), .A1(VRAMA[9]), .B1(w2554), .B2(VRAMA[8]), .A2(w2553) );
	vdp_and g2593 (.Z(w2673), .A(VRAMA[1]), .B(M5) );
	vdp_aon22 g2594 (.Z(w2469), .A1(w2671), .B1(w2576), .B2(VRAMA[15]), .A2(w2575) );
	vdp_aon22 g2595 (.Z(w2470), .A1(VRAMA[15]), .B1(w2576), .B2(VRAMA[14]), .A2(w2575) );
	vdp_aon22 g2596 (.Z(w2478), .A1(VRAMA[14]), .B1(w2576), .B2(VRAMA[13]), .A2(w2575) );
	vdp_aon22 g2597 (.Z(w2722), .A1(VRAMA[12]), .B1(w2576), .B2(VRAMA[11]), .A2(w2527) );
	vdp_aon22 g2598 (.Z(w2530), .A1(VRAMA[13]), .B1(w2576), .B2(VRAMA[12]), .A2(w2575) );
	vdp_aon22 g2599 (.Z(w2532), .A1(VRAMA[11]), .B1(w2576), .B2(VRAMA[10]), .A2(w2527) );
	vdp_aon22 g2600 (.Z(w2726), .A1(VRAMA[10]), .B1(w2576), .B2(w2605), .A2(w2527) );
	vdp_aon22 g2601 (.Z(w2538), .A1(w2673), .B1(w2576), .B2(VRAMA[0]), .A2(w2527) );
	vdp_aon22 g2602 (.Z(w2671), .A1(w2733), .B1(w111), .B2(w94), .A2(VRAMA[16]) );
	vdp_aon222 g2603 (.Z(w2541), .A1(w2524), .A2(w2523), .B1(w2707), .B2(w2710), .C1(w2706), .C2(w2620) );
	vdp_aon222 g2604 (.Z(w2546), .A1(w2524), .A2(w2542), .B1(w2707), .B2(w2701), .C1(w2706), .C2(w2607) );
	vdp_aon222 g2605 (.Z(w2550), .A1(w2524), .A2(w2700), .B1(w2707), .B2(w2608), .C1(w2706), .C2(w2552) );
	vdp_aon222 g2606 (.Z(w2709), .A1(w2524), .A2(w2612), .B1(w2707), .B2(w2610), .C1(w2706), .C2(w2604) );
	vdp_aon222 g2607 (.Z(w2562), .A1(w2524), .A2(w2555), .B1(w2707), .B2(w2603), .C1(w2706), .C2(w2602) );
	vdp_aon222 g2608 (.Z(w2708), .A1(w2524), .A2(w2559), .B1(w2707), .B2(w2672), .C1(w2706), .C2(w2563) );
	vdp_aon222 g2609 (.Z(w2657), .A1(w2524), .A2(w2480), .B1(w2707), .B2(w2705), .C1(w2706), .C2(w2561) );
	vdp_aon222 g2610 (.Z(w2465), .A1(w2524), .A2(w2472), .B1(w2707), .B2(w2599), .C1(w2706), .C2(w2598) );
	vdp_dlatch_inv g2611 (.nQ(w2622), .D(w2704), .C(HCLK1), .nC(nHCLK1) );
	vdp_comp_we g2612 (.Z(w2564), .A(w2624) );
	vdp_aon22 g2613 (.Z(nRAS1), .A1(1'b1), .B1(w2565), .B2(w2506), .A2(w2564) );
	vdp_aoi22 g2614 (.Z(w2581), .A1(w2578), .B1(w2521), .B2(w2716), .A2(w2702) );
	vdp_and g2615 (.Z(w2644), .B(w2731), .A(DCLK2) );
	vdp_nor g2616 (.Z(w2727), .A(w2646), .B(RES) );
	vdp_sr_bit g2617 (.Q(w2646), .D(w2727), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_dlatch_inv g2618 (.nQ(w2728), .D(w2647), .C(DCLK1), .nC(nDCLK1) );
	vdp_and g2619 (.Z(w2729), .A(DCLK2), .B(w2728) );
	vdp_dlatch_inv g2620 (.nQ(w2731), .D(w2646), .C(DCLK1), .nC(nDCLK1) );
	vdp_not g2621 (.nZ(w2650), .A(w2652) );
	vdp_not g2622 (.nZ(w2649), .A(w2730) );
	vdp_neg_dff g2623 (.Q(w2652), .C(DCLK1), .D(1'b1), .R(w2644) );
	vdp_not g2624 (.A(w2646), .nZ(w2647) );
	vdp_neg_dff g2625 (.Q(w2730), .R(w2729), .C(DCLK1), .D(1'b1) );
	vdp_sr_bit g2626 (.Q(w2810), .D(w2802), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2627 (.Q(w2806), .D(w2805), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2628 (.Q(w3000), .D(w2806), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2629 (.Q(w2823), .D(w3000), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2630 (.Q(w2778), .D(RD_DATA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2631 (.Q(w2779), .D(RD_DATA[2]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2632 (.Q(w2780), .D(w324), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2633 (.Q(w2981), .D(w3003), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2634 (.Q(w3003), .D(w3004), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2635 (.Q(w3004), .D(w3005), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2636 (.Q(w3005), .D(w3006), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2637 (.Q(w3006), .D(w3007), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2638 (.Q(w3007), .D(w3008), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2639 (.Q(w3008), .D(w3009), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2640 (.Q(w3009), .D(w18), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2641 (.Q(w2788), .D(w2781), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2642 (.Q(w2786), .D(w3012), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2643 (.Q(w3040), .D(w3014), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2644 (.Q(w3014), .D(w2761), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2645 (.Q(w2761), .D(w108), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2646 (.Q(w2736), .D(w2735), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2647 (.Q(w2741), .D(w2884), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2648 (.Q(w2800), .D(w2996), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2649 (.Q(w2804), .D(w3011), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2650 (.Q(w2819), .D(w2812), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2651 (.Q(w2735), .D(w2815), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2652 (.Q(w2840), .D(w2817), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2653 (.Q(w2839), .D(w2885), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2654 (.Q(PLANE_A_PRIO), .D(w2831), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2655 (.Q(PLANE_B_PRIO), .D(w2832), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2656 (.Q(w2796), .D(w2833), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2657 (.Q(w2838), .D(w2837), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2658 (.Q(w2757), .D(w2836), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2659 (.Q(w2836), .D(w130), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2660 (.Q(w2758), .D(w3042), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2661 (.Q(w3042), .D(w129), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2662 (.Q(w2849), .D(w2822), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2663 (.Q(w2835), .D(w2834), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2664 (.Q(SPR_PRIO), .D(w2988), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2665 (.Q(w2846), .D(w175), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2666 (.Q(w2845), .D(w174), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2667 (.Q(w2750), .D(w2766), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2668 (.Q(w2755), .D(w2767), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2669 (.Q(w2752), .D(w2777), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2670 (.Q(w2743), .D(w2768), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2671 (.Q(w2762), .D(w2775), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2672 (.Q(w2742), .D(w2769), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2673 (.Q(w2737), .D(w2872), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2674 (.Q(w2747), .D(w2770), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2675 (.Q(w2753), .D(w2764), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_slatch g2676 (.nQ(w3038), .D(w2766), .C(w2763), .nC(w2760) );
	vdp_slatch g2677 (.nQ(w3039), .D(w2764), .C(w2763), .nC(w2760) );
	vdp_slatch g2678 (.nQ(w3037), .D(w2767), .C(w2763), .nC(w2760) );
	vdp_slatch g2679 (.nQ(w3036), .D(w2777), .C(w2763), .nC(w2760) );
	vdp_slatch g2680 (.nQ(w3035), .D(w2768), .C(w2763), .nC(w2760) );
	vdp_slatch g2681 (.nQ(w3034), .D(w2775), .C(w2763), .nC(w2760) );
	vdp_slatch g2682 (.nQ(w3033), .D(w2769), .C(w2763), .nC(w2760) );
	vdp_slatch g2683 (.nQ(w3032), .D(w2872), .C(w2763), .nC(w2760) );
	vdp_slatch g2684 (.nQ(w3031), .D(w2770), .C(w2763), .nC(w2760) );
	vdp_slatch g2685 (.Q(w2821), .D(w617), .nC(w2799), .C(w2809) );
	vdp_slatch g2686 (.Q(w2818), .D(w681), .nC(w2799), .C(w2809) );
	vdp_slatch g2687 (.Q(w2811), .D(w725), .nC(w2799), .C(w2809) );
	vdp_slatch g2688 (.Q(w2807), .D(w719), .nC(w2799), .C(w2809) );
	vdp_slatch g2689 (.Q(w2803), .D(w698), .nC(w2799), .C(w2809) );
	vdp_slatch g2690 (.Q(w2999), .D(w685), .nC(w2799), .C(w2809) );
	vdp_slatch g2691 (.Q(w2801), .D(w612), .nC(w2799), .C(w2809) );
	vdp_slatch g2692 (.Q(w2974), .D(w661), .nC(w2799), .C(w2809) );
	vdp_aon2222 g2693 (.Z(w2951), .B2(w2890), .B1(w2895), .A2(w3026), .A1(w2890), .D2(w2886), .D1(w2895), .C2(w2895), .C1(w2887) );
	vdp_aon22 g2694 (.Z(w2916), .B2(w2886), .B1(w2900), .A2(w3027), .A1(w2891) );
	vdp_aon22 g2695 (.Z(w2921), .B2(w2886), .B1(w2896), .A2(w3026), .A1(w2891) );
	vdp_not g2696 (.nZ(w2904), .A(w2950) );
	vdp_not g2697 (.nZ(w2898), .A(w2899) );
	vdp_not g2698 (.nZ(w2903), .A(w2902) );
	vdp_not g2699 (.nZ(w2922), .A(w2951) );
	vdp_not g2700 (.nZ(w2915), .A(w2908) );
	vdp_buf g2701 (.Z(w2890), .A(w2786) );
	vdp_not g2702 (.nZ(w2985), .A(w2943) );
	vdp_not g2703 (.nZ(w2946), .A(w2944) );
	vdp_not g2704 (.nZ(w2947), .A(w2948) );
	vdp_not g2705 (.nZ(w2911), .A(w2887) );
	vdp_sr_bit g2706 (.Q(w2910), .D(w2758), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2707 (.Q(w2948), .D(w2756), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2708 (.Q(w2887), .D(w2757), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2709 (.Q(w2943), .D(w2945), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2710 (.Q(w2944), .D(w2782), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g2711 (.Z(w3022), .A(w2947), .B(w2985), .C(w2944) );
	vdp_and3 g2712 (.Z(w3024), .A(w2946), .B(w2948), .C(w2985) );
	vdp_and3 g2713 (.Z(w3023), .A(w2947), .B(w2985), .C(w2946) );
	vdp_and3 g2714 (.Z(w2909), .A(w2985), .B(w2944), .C(w2948) );
	vdp_and3 g2715 (.Z(w2907), .A(w2947), .B(w2943), .C(w2946) );
	vdp_and3 g2716 (.Z(w2905), .A(w2943), .B(w2944), .C(w2948) );
	vdp_and3 g2717 (.Z(w3025), .A(w2947), .B(w2944), .C(w2943) );
	vdp_and3 g2718 (.Z(w2906), .A(w2946), .B(w2948), .C(w2943) );
	vdp_sr_bit g2719 (.Q(w2902), .D(w2949), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2720 (.Q(w2899), .D(w2746), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2721 (.Q(w2950), .D(w2783), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g2722 (.Z(w2901), .A(w2903), .B(w2904), .C(w2898) );
	vdp_and3 g2723 (.Z(w2900), .A(w2898), .B(w2902), .C(w2904) );
	vdp_and3 g2724 (.Z(w3027), .A(w2903), .B(w2904), .C(w2899) );
	vdp_and3 g2725 (.Z(w2896), .A(w2904), .B(w2899), .C(w2902) );
	vdp_and3 g2726 (.Z(w2897), .A(w2898), .B(w2902), .C(w2950) );
	vdp_and3 g2727 (.Z(w2894), .A(w2903), .B(w2950), .C(w2898) );
	vdp_and3 g2728 (.Z(w3026), .A(w2903), .B(w2899), .C(w2950) );
	vdp_and3 g2729 (.Z(w2895), .A(w2950), .B(w2899), .C(w2902) );
	vdp_not g2730 (.nZ(w2984), .A(w3041) );
	vdp_not g2731 (.nZ(w2939), .A(w2941) );
	vdp_not g2732 (.nZ(w2940), .A(w2942) );
	vdp_sr_bit g2733 (.Q(w2941), .D(w2980), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2734 (.Q(w2942), .D(w2978), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2735 (.Q(w3041), .D(w2744), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g2736 (.Z(w2893), .A(w2940), .B(w2984), .C(w2939) );
	vdp_and3 g2737 (.Z(w2892), .A(w2939), .B(w2942), .C(w2984) );
	vdp_and3 g2738 (.A(w2940), .B(w2984), .C(w2941), .Z(w2889) );
	vdp_and3 g2739 (.Z(w3028), .A(w2984), .B(w2941), .C(w2942) );
	vdp_and3 g2740 (.Z(w2888), .A(w2940), .B(w3041), .C(w2939) );
	vdp_and3 g2741 (.Z(w3030), .A(w2939), .B(w2942), .C(w3041) );
	vdp_and3 g2742 (.Z(w2983), .A(w3041), .B(w2941), .C(w2942) );
	vdp_and3 g2743 (.Z(w3029), .A(w2940), .B(w2941), .C(w3041) );
	vdp_aon22 g2744 (.nZ(w2973), .B2(w2886), .B1(w3029), .A2(w3030), .A1(w2887) );
	vdp_aon22 g2745 (.nZ(w2938), .B2(w2886), .B1(w2888), .A2(w2892), .A1(w2887) );
	vdp_aon22 g2746 (.nZ(w2972), .B2(w2887), .B1(w2893), .A2(w2983), .A1(w2891) );
	vdp_and g2747 (.nZ(w2937), .B(w2887), .A(w2888) );
	vdp_and g2748 (.nZ(w2971), .B(w2887), .A(w3029) );
	vdp_and g2749 (.nZ(w2970), .B(w2887), .A(w2889) );
	vdp_aon22 g2750 (.nZ(w2969), .B2(w2890), .B1(w3030), .A2(w2888), .A1(w2890) );
	vdp_aon22 g2751 (.nZ(w2968), .B2(w2886), .B1(w3030), .A2(w3028), .A1(w2887) );
	vdp_aon2222 g2752 (.Z(w2952), .B2(w2890), .B1(w2983), .A2(w3029), .A1(w2890), .D2(w2886), .D1(w2983), .C2(w2983), .C1(w2887) );
	vdp_aon22 g2753 (.Z(w2935), .B2(w2886), .B1(w2892), .A2(w2889), .A1(w2891) );
	vdp_aon22 g2754 (.Z(w2932), .B2(w2886), .B1(w3028), .A2(w3029), .A1(w2891) );
	vdp_and g2755 (.Z(w2936), .B(w3030), .A(w2891) );
	vdp_and g2756 (.Z(w2931), .B(w2891), .A(w3028) );
	vdp_and g2757 (.Z(w2933), .B(w2892), .A(w2891) );
	vdp_aon22 g2758 (.Z(w2930), .B2(w2890), .B1(w3028), .A2(w2889), .A1(w2890) );
	vdp_aon22 g2759 (.Z(w2929), .B2(w2886), .B1(w2889), .A2(w2888), .A1(w2891) );
	vdp_aon2222 g2760 (.Z(w2967), .B2(w2890), .B1(w2892), .A2(w2893), .A1(w2890), .D2(w2886), .D1(w2893), .C2(w2893), .C1(w2891) );
	vdp_not g2761 (.nZ(w2934), .A(w2952) );
	vdp_aon22 g2762 (.nZ(w2966), .B2(w2886), .B1(w3026), .A2(w2897), .A1(w2887) );
	vdp_aon22 g2763 (.nZ(w2965), .B2(w2886), .B1(w2894), .A2(w2900), .A1(w2887) );
	vdp_aon22 g2764 (.nZ(w2928), .B2(w2887), .B1(w2901), .A2(w2895), .A1(w2891) );
	vdp_and g2765 (.nZ(w2927), .B(w2887), .A(w2894) );
	vdp_and g2766 (.nZ(w2926), .B(w2887), .A(w3026) );
	vdp_and g2767 (.nZ(w2925), .B(w2887), .A(w3027) );
	vdp_aon22 g2768 (.nZ(w2924), .B2(w2890), .B1(w2897), .A2(w2894), .A1(w2890) );
	vdp_aon22 g2769 (.nZ(w2923), .B2(w2886), .B1(w2897), .A2(w2896), .A1(w2887) );
	vdp_and g2770 (.Z(w2920), .B(w2897), .A(w2891) );
	vdp_and g2771 (.Z(w3019), .B(w2891), .A(w2896) );
	vdp_and g2772 (.Z(w2919), .B(w2900), .A(w2891) );
	vdp_aon22 g2773 (.Z(w2918), .B2(w2890), .B1(w2896), .A2(w3027), .A1(w2890) );
	vdp_aon22 g2774 (.Z(w2917), .B2(w2886), .B1(w3027), .A2(w2894), .A1(w2891) );
	vdp_aon2222 g2775 (.Z(w3020), .B2(w2890), .B1(w2900), .A2(w2901), .A1(w2890), .D2(w2886), .D1(w2901), .C2(w2901), .C1(w2891) );
	vdp_aon22 g2776 (.nZ(w2914), .B2(w2886), .B1(w3025), .A2(w2906), .A1(w2887) );
	vdp_aon22 g2777 (.nZ(w2964), .B2(w2886), .B1(w2907), .A2(w3024), .A1(w2887) );
	vdp_aon22 g2778 (.nZ(w2960), .B2(w2887), .B1(w3023), .A2(w2905), .A1(w2891) );
	vdp_and g2779 (.nZ(w2961), .B(w2887), .A(w2907) );
	vdp_and g2780 (.nZ(w2962), .B(w2887), .A(w3025) );
	vdp_and g2781 (.nZ(w2959), .B(w2887), .A(w3022) );
	vdp_aon22 g2782 (.nZ(w2963), .B2(w2890), .B1(w2906), .A2(w2907), .A1(w2890) );
	vdp_aon22 g2783 (.nZ(w3021), .B2(w2886), .B1(w2906), .A2(w2909), .A1(w2887) );
	vdp_aon2222 g2784 (.Z(w2908), .B2(w2890), .B1(w2905), .A2(w3025), .A1(w2890), .D2(w2886), .D1(w2905), .C2(w2905), .C1(w2887) );
	vdp_aon22 g2785 (.Z(w2912), .B2(w2886), .B1(w3024), .A2(w3022), .A1(w2891) );
	vdp_aon22 g2786 (.Z(w2913), .B2(w2890), .B1(w2909), .A2(w3022), .A1(w2890) );
	vdp_aon22 g2787 (.Z(w2958), .B2(w2886), .B1(w2909), .A2(w3025), .A1(w2891) );
	vdp_and g2788 (.Z(w2957), .B(w2891), .A(w2909) );
	vdp_and g2789 (.Z(w2956), .B(w3024), .A(w2891) );
	vdp_and g2790 (.Z(w2955), .B(w2891), .A(w2906) );
	vdp_aon22 g2791 (.Z(w2953), .B2(w2886), .B1(w3022), .A2(w2907), .A1(w2891) );
	vdp_aon2222 g2792 (.Z(w2954), .B2(w2890), .B1(w3024), .A2(w3023), .A1(w2890), .D2(w2886), .D1(w3023), .C2(w3023), .C1(w2891) );
	vdp_nor3 g2793 (.Z(w2886), .A(w2890), .B(w2910), .C(w2887) );
	vdp_and g2794 (.Z(w2891), .A(w2910), .B(w2911) );
	vdp_bufif0 g2795 (.A(w2801), .nE(w2808), .Z(COL[0]) );
	vdp_bufif0 g2796 (.A(w2999), .nE(w2808), .Z(COL[1]) );
	vdp_bufif0 g2797 (.A(w2803), .nE(w2808), .Z(COL[2]) );
	vdp_bufif0 g2798 (.A(w2807), .nE(w2808), .Z(COL[3]) );
	vdp_bufif0 g2799 (.A(w2820), .nE(w2808), .Z(COL[4]) );
	vdp_bufif0 g2800 (.A(w2998), .nE(w2808), .Z(COL[5]) );
	vdp_and g2801 (.Z(w2998), .A(M5), .B(w2818) );
	vdp_or g2802 (.Z(w2820), .A(w2791), .B(w2811) );
	vdp_not g2803 (.nZ(w2682), .A(M5) );
	vdp_not g2804 (.nZ(w2789), .A(w2997) );
	vdp_not g2805 (.nZ(w2790), .A(w2792) );
	vdp_not g2806 (.nZ(w2791), .A(M5) );
	vdp_not g2807 (.nZ(w2787), .A(w2793) );
	vdp_not g2808 (.nZ(w2808), .A(w2796) );
	vdp_comp_strong g2809 (.nZ(w2799), .Z(w2809), .A(w73) );
	vdp_not g2810 (.nZ(w2797), .A(w101) );
	vdp_not g2811 (.nZ(w3010), .A(w19) );
	vdp_aon222 g2812 (.Z(w2996), .B2(w2789), .A2(w2790), .A1(VRAMA[0]), .B1(VRAMA[1]), .C2(w2787), .C1(COL[0]) );
	vdp_aon222 g2813 (.Z(w3011), .B2(w2789), .A2(w2790), .A1(VRAMA[1]), .B1(VRAMA[2]), .C2(w2787), .C1(COL[1]) );
	vdp_aon222 g2814 (.Z(w2802), .B2(w2789), .A2(w2790), .A1(VRAMA[2]), .B1(VRAMA[3]), .C2(w2787), .C1(COL[2]) );
	vdp_aon222 g2815 (.Z(w2812), .B2(w2789), .A2(w2790), .A1(VRAMA[3]), .B1(VRAMA[4]), .C2(w2787), .C1(COL[3]) );
	vdp_aon222 g2816 (.Z(w2817), .B2(w2789), .A2(w2790), .A1(VRAMA[4]), .B1(VRAMA[5]), .C2(w2787), .C1(COL[4]) );
	vdp_aon222 g2817 (.Z(w2885), .B2(w2789), .A2(w2790), .A1(1'b0), .B1(VRAMA[6]), .C2(w2787), .C1(COL[5]) );
	vdp_nand g2818 (.Z(w2997), .A(w2793), .B(M5) );
	vdp_nand g2819 (.Z(w2792), .A(w2793), .B(w2791) );
	vdp_and g2820 (.Z(w2822), .A(w2823), .B(w3049) );
	vdp_aon222 g2821 (.Z(w3049), .B2(w3044), .A2(w2828), .A1(w2784), .B1(w2830), .C2(w3043), .C1(w2851) );
	vdp_not g2822 (.nZ(w3044), .A(w2995) );
	vdp_not g2823 (.nZ(w3043), .A(w2785) );
	vdp_not g2824 (.nZ(w2856), .A(w2841) );
	vdp_nor g2825 (.Z(w2830), .A(w2785), .B(w2988) );
	vdp_nor g2826 (.Z(w2995), .A(w2851), .B(w2850) );
	vdp_and g2827 (.Z(w2829), .A(w2824), .B(w2864) );
	vdp_and g2828 (.Z(w2828), .A(w2841), .B(w2855) );
	vdp_and g2829 (.Z(w2858), .A(w2855), .B(w2856) );
	vdp_or g2830 (.Z(w2988), .A(w2859), .B(w2858) );
	vdp_or g2831 (.Z(w2827), .A(w2784), .B(w2785) );
	vdp_and g2832 (.Z(w2798), .A(w2823), .B(w2797) );
	vdp_and g2833 (.Z(w2977), .A(w2824), .B(w2861) );
	vdp_and g2834 (.Z(w2987), .A(w2825), .B(w2863) );
	vdp_not g2835 (.nZ(w2869), .A(w101) );
	vdp_or g2836 (.Z(w2831), .A(w2862), .B(w2848) );
	vdp_not g2837 (.nZ(w3047), .A(w2825) );
	vdp_not g2838 (.nZ(w2975), .A(w2724) );
	vdp_not g2839 (.nZ(w2853), .A(w2842) );
	vdp_not g2840 (.nZ(w2852), .A(w2843) );
	vdp_not g2841 (.nZ(w2857), .A(w2725) );
	vdp_and g2842 (.Z(w2876), .A(w2825), .B(w2860) );
	vdp_and g2843 (.Z(w2854), .A(w2826), .B(w2866) );
	vdp_not g2844 (.nZ(w2986), .A(w98) );
	vdp_not g2845 (.nZ(w2993), .A(w99) );
	vdp_and g2846 (.Z(w2859), .A(w2993), .B(w98) );
	vdp_and g2847 (.Z(w2862), .A(w2986), .B(w99) );
	vdp_and g2848 (.Z(w2875), .A(w98), .B(w99) );
	vdp_or3 g2849 (.Z(w2793), .A(w108), .B(w174), .C(w175) );
	vdp_and3 g2850 (.Z(w2992), .A(w2826), .B(w2825), .C(w2863) );
	vdp_and3 g2851 (.Z(w2861), .A(w2852), .B(w2842), .C(w2725) );
	vdp_and3 g2852 (.Z(w2860), .A(w2853), .B(w2843), .C(w2857) );
	vdp_and3 g2853 (.Z(w2866), .A(w2852), .B(w2842), .C(w2857) );
	vdp_and3 g2854 (.Z(w2863), .A(w2842), .B(w2843), .C(w2857) );
	vdp_and g2855 (.Z(w2982), .A(M5), .B(w89) );
	vdp_or g2856 (.Z(w2824), .A(w2975), .B(w2841) );
	vdp_and3 g2857 (.Z(w2834), .A(w2828), .B(w2785), .C(w2995) );
	vdp_and3 g2858 (.Z(w2991), .A(w2826), .B(w2824), .C(w2861) );
	vdp_and3 g2859 (.Z(w2990), .A(w2826), .B(w2824), .C(w2866) );
	vdp_and3 g2860 (.Z(w2848), .A(w2847), .B(w2798), .C(w3047) );
	vdp_and3 g2861 (.Z(w2841), .A(w2827), .B(w2844), .C(w2982) );
	vdp_and3 g2862 (.Z(w2870), .A(w2825), .B(w2824), .C(w2864) );
	vdp_and3 g2863 (.Z(w3046), .A(w2825), .B(w2824), .C(w2860) );
	vdp_and3 g2864 (.Z(w2867), .A(w2826), .B(w2825), .C(w2824) );
	vdp_and3 g2865 (.Z(w2868), .A(w2798), .B(w2865), .C(w3045) );
	vdp_and g2866 (.Z(w2833), .A(w2976), .B(w2989) );
	vdp_not g2867 (.nZ(w2871), .A(w2798) );
	vdp_not g2868 (.nZ(w3045), .A(w2826) );
	vdp_or g2869 (.Z(w2832), .A(w2875), .B(w2868) );
	vdp_or g2870 (.Z(w2989), .A(w2871), .B(w2867) );
	vdp_not g2871 (.nZ(w3002), .A(M5) );
	vdp_notif0 g2872 (.A(w3039), .nE(w2765), .nZ(w324) );
	vdp_notif0 g2873 (.nZ(RD_DATA[2]), .A(w3038), .nE(w2765) );
	vdp_notif0 g2874 (.nZ(RD_DATA[1]), .A(w3037), .nE(w2765) );
	vdp_notif0 g2875 (.nZ(AD_DATA[7]), .A(w3036), .nE(w2765) );
	vdp_notif0 g2876 (.nZ(AD_DATA[6]), .A(w3035), .nE(w2765) );
	vdp_notif0 g2877 (.nZ(AD_DATA[5]), .A(w3034), .nE(w2765) );
	vdp_notif0 g2878 (.nZ(AD_DATA[3]), .A(w3033), .nE(w2765) );
	vdp_notif0 g2879 (.nZ(AD_DATA[2]), .A(w3032), .nE(w2765) );
	vdp_notif0 g2880 (.nZ(w2734), .A(w3031), .nE(w2765) );
	vdp_notif0 g2881 (.nZ(DB[1]), .A(w2758), .nE(w2749) );
	vdp_notif0 g2882 (.A(w2757), .nE(w2749) );
	vdp_notif0 g2883 (.nZ(DB[2]), .A(w2978), .nE(w2749) );
	vdp_notif0 g2884 (.nZ(DB[5]), .A(w2949), .nE(w2749) );
	vdp_notif0 g2885 (.nZ(DB[8]), .A(w2756), .nE(w2749) );
	vdp_notif0 g2886 (.nZ(DB[10]), .A(w2945), .nE(w2749) );
	vdp_notif0 g2887 (.nZ(DB[9]), .A(w2782), .nE(w2749) );
	vdp_notif0 g2888 (.nZ(w160), .A(w2783), .nE(w2749) );
	vdp_notif0 g2889 (.nZ(DB[6]), .A(w2746), .nE(w2749) );
	vdp_notif0 g2890 (.nZ(DB[4]), .A(w2744), .nE(w2749) );
	vdp_comp_we g2891 (.A(M5), .nZ(w2739), .Z(w2738) );
	vdp_notif0 g2892 (.nZ(w156), .A(w2980), .nE(w2749) );
	vdp_not g2893 (.A(w88), .nZ(w2749) );
	vdp_and g2894 (.Z(w2740), .A(w2741), .B(w2736) );
	vdp_and3 g2895 (.Z(w2980), .A(w97), .B(w2741), .C(w2979) );
	vdp_and3 g2896 (.Z(w2744), .A(w97), .B(w2741), .C(w3013) );
	vdp_and3 g2897 (.Z(w2746), .A(w97), .B(w2741), .C(w2745) );
	vdp_and3 g2898 (.Z(w2783), .A(w97), .B(w2741), .C(w2748) );
	vdp_and3 g2899 (.Z(w2782), .A(w97), .B(w2741), .C(w2751) );
	vdp_and3 g2900 (.Z(w2945), .A(w97), .B(w2741), .C(w2754) );
	vdp_and3 g2901 (.Z(w2756), .A(M5), .B(w2741), .C(w2755) );
	vdp_and3 g2902 (.Z(w2949), .A(M5), .B(w2741), .C(w2762) );
	vdp_and3 g2903 (.Z(w2978), .A(M5), .B(w2741), .C(w2747) );
	vdp_comp_strong g2904 (.nZ(w2760), .A(w2759), .Z(w2763) );
	vdp_and g2905 (.Z(w2759), .A(w2761), .B(HCLK1) );
	vdp_not g2906 (.nZ(w2765), .A(w3040) );
	vdp_aon22 g2907 (.Z(w3001), .B2(FIFOo[5]), .A2(FIFOo[7]), .A1(w2814), .B1(w2813) );
	vdp_aon22 g2908 (.Z(w2776), .B2(FIFOo[4]), .A2(FIFOo[6]), .A1(w2814), .B1(w2813) );
	vdp_aon22 g2909 (.Z(w2774), .B2(FIFOo[3]), .A2(FIFOo[5]), .A1(w2814), .B1(w2813) );
	vdp_aon22 g2910 (.Z(w2773), .B2(FIFOo[2]), .A2(FIFOo[3]), .A1(w2814), .B1(w2813) );
	vdp_aon22 g2911 (.Z(w2772), .B2(FIFOo[1]), .A2(FIFOo[2]), .A1(w2814), .B1(w2813) );
	vdp_aon22 g2912 (.Z(w2771), .B2(FIFOo[0]), .A2(FIFOo[1]), .A1(w2814), .B1(w2813) );
	vdp_comp_we g2913 (.Z(w2814), .nZ(w2813), .A(M5) );
	vdp_aon22 g2914 (.Z(w2805), .B2(w3002), .A2(M5), .A1(w2981), .B1(w18) );
	vdp_aon22 g2915 (.Z(w130), .B2(w2835), .A2(w2821), .A1(w101), .B1(w2869) );
	vdp_aon22 g2916 (.Z(w129), .B2(w2849), .A2(w2974), .A1(w101), .B1(w2869) );
	vdp_and3 g2917 (.Z(w2855), .A(w2798), .B(w2724), .C(w3048) );
	vdp_aon22 g2918 (.Z(w2864), .B2(w2852), .A2(w2843), .A1(w2725), .B1(w2853) );
	vdp_aon22 g2919 (.Z(w2748), .B2(w2762), .A2(w2752), .A1(w2738), .B1(w2739) );
	vdp_aon22 g2920 (.Z(w2745), .B2(w2742), .A2(w2743), .A1(w2738), .B1(w2739) );
	vdp_aon22 g2921 (.Z(w2979), .B2(w2747), .A2(w2737), .A1(w2738), .B1(w2739) );
	vdp_aon22 g2922 (.Z(w3013), .B2(w2737), .A2(w2742), .A1(w2738), .B1(w2739) );
	vdp_aon22 g2923 (.Z(w2751), .B2(w2743), .A2(w2750), .A1(w2738), .B1(w2739) );
	vdp_aon22 g2924 (.Z(w2754), .B2(w2752), .A2(w2753), .A1(w2738), .B1(w2739) );
	vdp_g2925 g2925 (.Z(w2850), .A(w2853), .B(w2725), .C(w2982), .D(w2852) );
	vdp_or5 g2926 (.Z(w2847), .A(w2829), .B(w2860), .C(w2863), .D(w2991), .E(w2990) );
	vdp_or5 g2927 (.Z(w2865), .A(w2870), .B(w2866), .C(w2977), .D(w2987), .E(w3046) );
	vdp_or5 g2928 (.Z(w3048), .A(w2861), .B(w2864), .C(w2876), .D(w2854), .E(w2992) );
	vdp_nor4 g2929 (.Z(w2815), .A(COL[2]), .B(COL[3]), .C(COL[1]), .D(COL[0]) );
	vdp_nor g2930 (.Z(w2976), .A(w98), .B(w99) );
	vdp_nor g2931 (.Z(w2825), .A(w2994), .B(w2874) );
	vdp_nor g2932 (.Z(w2994), .A(w2724), .B(M5) );
	vdp_nand g2933 (.Z(w2826), .A(M5), .B(w2873) );
	vdp_nand g2934 (.Z(w2837), .A(SPR_PRIO), .B(w19) );
	vdp_and4 g2935 (.Z(w2851), .A(w2852), .B(w2982), .C(w2853), .D(w2857) );
	vdp_aoi21 g2936 (.Z(w3012), .B(w2740), .A2(w3010), .A1(w2788) );
	vdp_nor g2937 (.Z(w2884), .A(w21), .B(w20) );
	vdp_g2938 g2938 (.A(w2796), .Z(COL[6]) );
	vdp_slatch g2939 (.Q(w4159), .D(S[3]), .C(w3178), .nC(w3168) );
	vdp_slatch g2940 (.Q(w4161), .D(S[3]), .C(w3159), .nC(w3158) );
	vdp_slatch g2941 (.Q(w4163), .D(S[3]), .C(w3160), .nC(w3156) );
	vdp_slatch g2942 (.Q(w4165), .D(S[3]), .C(w3177), .nC(w3169) );
	vdp_slatch g2943 (.Q(w4167), .D(S[7]), .C(w3178), .nC(w3168) );
	vdp_slatch g2944 (.Q(w4170), .D(S[7]), .C(w3159), .nC(w3158) );
	vdp_slatch g2945 (.Q(w4169), .D(S[7]), .C(w3160), .nC(w3156) );
	vdp_slatch g2946 (.Q(w4174), .D(S[7]), .C(w3177), .nC(w3169) );
	vdp_slatch g2947 (.Q(w4173), .D(S[2]), .C(w3178), .nC(w3168) );
	vdp_slatch g2948 (.Q(w4180), .D(S[2]), .C(w3159), .nC(w3158) );
	vdp_slatch g2949 (.Q(w4179), .D(S[2]), .C(w3160), .nC(w3156) );
	vdp_slatch g2950 (.Q(w4182), .D(S[2]), .C(w3177), .nC(w3169) );
	vdp_slatch g2951 (.Q(w4181), .D(S[6]), .C(w3178), .nC(w3168) );
	vdp_slatch g2952 (.Q(w4186), .D(S[6]), .C(w3159), .nC(w3158) );
	vdp_slatch g2953 (.Q(w4185), .D(S[6]), .C(w3160), .nC(w3156) );
	vdp_slatch g2954 (.Q(w4190), .D(S[6]), .C(w3177), .nC(w3169) );
	vdp_slatch g2955 (.Q(w4189), .D(S[1]), .C(w3178), .nC(w3168) );
	vdp_slatch g2956 (.Q(w4194), .D(S[1]), .C(w3159), .nC(w3158) );
	vdp_slatch g2957 (.Q(w4193), .D(S[1]), .C(w3160), .nC(w3156) );
	vdp_slatch g2958 (.Q(w4198), .D(S[1]), .C(w3177), .nC(w3169) );
	vdp_slatch g2959 (.Q(w4197), .D(S[5]), .C(w3178), .nC(w3168) );
	vdp_slatch g2960 (.Q(w4202), .D(S[5]), .C(w3159), .nC(w3158) );
	vdp_slatch g2961 (.Q(w4201), .D(S[5]), .C(w3160), .nC(w3156) );
	vdp_slatch g2962 (.Q(w4206), .D(S[5]), .C(w3177), .nC(w3169) );
	vdp_slatch g2963 (.Q(w4205), .D(S[0]), .C(w3178), .nC(w3168) );
	vdp_slatch g2964 (.Q(w4210), .D(S[0]), .C(w3159), .nC(w3158) );
	vdp_slatch g2965 (.Q(w4209), .D(S[0]), .C(w3160), .nC(w3156) );
	vdp_slatch g2966 (.Q(w4214), .D(S[0]), .C(w3177), .nC(w3169) );
	vdp_slatch g2967 (.Q(w4213), .D(S[4]), .C(w3178), .nC(w3168) );
	vdp_slatch g2968 (.Q(w4218), .D(S[4]), .C(w3159), .nC(w3158) );
	vdp_slatch g2969 (.Q(w4217), .D(S[4]), .C(w3160), .nC(w3156) );
	vdp_slatch g2970 (.Q(w4221), .D(S[4]), .C(w3177), .nC(w3169) );
	vdp_slatch g2971 (.Q(w4160), .D(w4159), .C(w3148), .nC(w3165) );
	vdp_slatch g2972 (.Q(w4162), .D(w4161), .C(w3166), .nC(w3157) );
	vdp_slatch g2973 (.Q(w4164), .D(w4163), .C(w3167), .nC(w3155) );
	vdp_slatch g2974 (.Q(w4166), .D(w4165), .C(w3163), .nC(w3164) );
	vdp_slatch g2975 (.Q(w4168), .D(w4167), .C(w3148), .nC(w3165) );
	vdp_slatch g2976 (.Q(w4172), .D(w4170), .C(w3166), .nC(w3157) );
	vdp_slatch g2977 (.Q(w4171), .D(w4169), .C(w3167), .nC(w3155) );
	vdp_slatch g2978 (.Q(w4176), .D(w4174), .C(w3163), .nC(w3164) );
	vdp_slatch g2979 (.Q(w4175), .D(w4173), .C(w3148), .nC(w3165) );
	vdp_slatch g2980 (.Q(w4178), .D(w4180), .C(w3166), .nC(w3157) );
	vdp_slatch g2981 (.Q(w4177), .D(w4179), .C(w3167), .nC(w3155) );
	vdp_slatch g2982 (.Q(w4184), .D(w4182), .C(w3163), .nC(w3164) );
	vdp_slatch g2983 (.Q(w4183), .D(w4181), .C(w3148), .nC(w3165) );
	vdp_slatch g2984 (.Q(w4188), .D(w4186), .C(w3166), .nC(w3157) );
	vdp_slatch g2985 (.Q(w4187), .D(w4185), .C(w3167), .nC(w3155) );
	vdp_slatch g2986 (.Q(w4192), .D(w4190), .C(w3163), .nC(w3164) );
	vdp_slatch g2987 (.Q(w4191), .D(w4189), .C(w3148), .nC(w3165) );
	vdp_slatch g2988 (.Q(w4196), .D(w4194), .C(w3166), .nC(w3157) );
	vdp_slatch g2989 (.Q(w4195), .D(w4193), .C(w3167), .nC(w3155) );
	vdp_slatch g2990 (.Q(w4200), .D(w4198), .C(w3163), .nC(w3164) );
	vdp_slatch g2991 (.Q(w4199), .D(w4197), .C(w3148), .nC(w3165) );
	vdp_slatch g2992 (.Q(w4204), .D(w4202), .C(w3166), .nC(w3157) );
	vdp_slatch g2993 (.Q(w4203), .D(w4201), .C(w3167), .nC(w3155) );
	vdp_slatch g2994 (.Q(w4208), .D(w4206), .C(w3163), .nC(w3164) );
	vdp_slatch g2995 (.Q(w4207), .D(w4205), .C(w3148), .nC(w3165) );
	vdp_slatch g2996 (.Q(w4212), .D(w4210), .C(w3166), .nC(w3157) );
	vdp_slatch g2997 (.Q(w4211), .D(w4209), .C(w3167), .nC(w3155) );
	vdp_slatch g2998 (.Q(w4216), .D(w4214), .C(w3163), .nC(w3164) );
	vdp_slatch g2999 (.Q(w4215), .D(w4213), .C(w3148), .nC(w3165) );
	vdp_slatch g3000 (.Q(w4220), .D(w4218), .C(w3166), .nC(w3157) );
	vdp_slatch g3001 (.Q(w4219), .D(w4217), .C(w3167), .nC(w3155) );
	vdp_slatch g3002 (.Q(w4222), .D(w4221), .C(w3163), .nC(w3164) );
	vdp_slatch g3003 (.Q(w3205), .D(w4160), .C(w3170), .nC(w3196) );
	vdp_slatch g3004 (.Q(w3204), .D(w4162), .C(w3149), .nC(w3206) );
	vdp_slatch g3005 (.Q(w3203), .D(w4164), .C(w3161), .nC(w3207) );
	vdp_slatch g3006 (.Q(w3202), .D(w4166), .C(w3162), .nC(w3136) );
	vdp_slatch g3007 (.Q(w3201), .D(w4168), .C(w3170), .nC(w3196) );
	vdp_slatch g3008 (.Q(w3200), .D(w4172), .C(w3149), .nC(w3206) );
	vdp_slatch g3009 (.Q(w3199), .D(w4171), .C(w3161), .nC(w3207) );
	vdp_slatch g3010 (.Q(w3198), .D(w4176), .C(w3162), .nC(w3136) );
	vdp_slatch g3011 (.Q(w3197), .D(w4175), .C(w3170), .nC(w3196) );
	vdp_slatch g3012 (.Q(w3210), .D(w4178), .C(w3149), .nC(w3206) );
	vdp_slatch g3013 (.Q(w3214), .D(w4177), .C(w3161), .nC(w3207) );
	vdp_slatch g3014 (.Q(w3213), .D(w4184), .C(w3162), .nC(w3136) );
	vdp_slatch g3015 (.Q(w3212), .D(w4183), .C(w3170), .nC(w3196) );
	vdp_slatch g3016 (.Q(w3208), .D(w4188), .C(w3149), .nC(w3206) );
	vdp_slatch g3017 (.Q(w3209), .D(w4187), .C(w3161), .nC(w3207) );
	vdp_slatch g3018 (.D(w4192), .Q(w3211), .C(w3162), .nC(w3136) );
	vdp_slatch g3019 (.Q(w3215), .D(w4191), .C(w3170), .nC(w3196) );
	vdp_slatch g3020 (.Q(w3216), .D(w4196), .C(w3149), .nC(w3206) );
	vdp_slatch g3021 (.Q(w3218), .D(w4195), .C(w3161), .nC(w3207) );
	vdp_slatch g3022 (.Q(w3217), .D(w4200), .C(w3162), .nC(w3136) );
	vdp_slatch g3023 (.Q(w3260), .D(w4199), .C(w3170), .nC(w3196) );
	vdp_slatch g3024 (.Q(w3261), .D(w4204), .C(w3149), .nC(w3206) );
	vdp_slatch g3025 (.Q(w3257), .D(w4203), .C(w3161), .nC(w3207) );
	vdp_slatch g3026 (.Q(w3252), .D(w4208), .C(w3162), .nC(w3136) );
	vdp_slatch g3027 (.Q(w3264), .D(w4207), .C(w3170), .nC(w3196) );
	vdp_slatch g3028 (.Q(w3263), .D(w4212), .C(w3149), .nC(w3206) );
	vdp_slatch g3029 (.Q(w3262), .D(w4211), .C(w3161), .nC(w3207) );
	vdp_slatch g3030 (.Q(w3259), .D(w4216), .C(w3162), .nC(w3136) );
	vdp_slatch g3031 (.Q(w3245), .D(w4215), .C(w3170), .nC(w3196) );
	vdp_slatch g3032 (.Q(w3244), .D(w4220), .C(w3149), .nC(w3206) );
	vdp_slatch g3033 (.Q(w3246), .D(w4219), .C(w3161), .nC(w3207) );
	vdp_slatch g3034 (.Q(w3247), .D(w4222), .C(w3162), .nC(w3136) );
	vdp_slatch g3035 (.Q(w3324), .D(w4444), .C(w3321), .nC(w3322) );
	vdp_slatch g3036 (.Q(w3325), .D(w4445), .C(w3320), .nC(w3128) );
	vdp_slatch g3037 (.Q(w3326), .D(w4447), .C(w3319), .nC(w3330) );
	vdp_slatch g3038 (.Q(w3327), .D(w4446), .C(w3318), .nC(w3323) );
	vdp_slatch g3039 (.Q(w3328), .D(w4278), .C(w3321), .nC(w3322) );
	vdp_slatch g3040 (.Q(w3329), .D(w4277), .C(w3320), .nC(w3128) );
	vdp_slatch g3041 (.Q(w3334), .D(w4272), .C(w3319), .nC(w3330) );
	vdp_slatch g3042 (.Q(w3344), .D(w4271), .C(w3318), .nC(w3323) );
	vdp_slatch g3043 (.Q(w3336), .D(w4268), .C(w3321), .nC(w3322) );
	vdp_slatch g3044 (.Q(w3337), .D(w4267), .C(w3320), .nC(w3128) );
	vdp_slatch g3045 (.Q(w3338), .D(w4266), .C(w3319), .nC(w3330) );
	vdp_slatch g3046 (.Q(w3333), .D(w4263), .C(w3318), .nC(w3323) );
	vdp_slatch g3047 (.Q(w3339), .D(w4260), .C(w3321), .nC(w3322) );
	vdp_slatch g3048 (.Q(w3340), .D(w4261), .C(w3320), .nC(w3128) );
	vdp_slatch g3049 (.Q(w3341), .D(w4256), .C(w3319), .nC(w3330) );
	vdp_slatch g3050 (.Q(w3342), .D(w4257), .C(w3318), .nC(w3323) );
	vdp_slatch g3051 (.Q(w3268), .D(w4254), .C(w3321), .nC(w3322) );
	vdp_slatch g3052 (.Q(w4046), .D(w4253), .C(w3320), .nC(w3128) );
	vdp_slatch g3053 (.Q(w3270), .D(w4250), .C(w3319), .nC(w3330) );
	vdp_slatch g3054 (.Q(w3271), .D(w4249), .C(w3318), .nC(w3323) );
	vdp_slatch g3055 (.Q(w3343), .D(w4246), .C(w3321), .nC(w3322) );
	vdp_slatch g3056 (.Q(w3269), .D(w4245), .C(w3320), .nC(w3128) );
	vdp_slatch g3057 (.Q(w3249), .D(w4242), .C(w3319), .nC(w3330) );
	vdp_slatch g3058 (.Q(w3272), .D(w4241), .C(w3318), .nC(w3323) );
	vdp_slatch g3059 (.Q(w3275), .D(w4238), .C(w3321), .nC(w3322) );
	vdp_slatch g3060 (.Q(w3283), .D(w4237), .C(w3320), .nC(w3128) );
	vdp_slatch g3061 (.Q(w3282), .D(w4234), .C(w3319), .nC(w3330) );
	vdp_slatch g3062 (.Q(w3281), .D(w4233), .C(w3318), .nC(w3323) );
	vdp_slatch g3063 (.Q(w3279), .D(w4230), .C(w3321), .nC(w3322) );
	vdp_slatch g3064 (.Q(w3273), .D(w4229), .C(w3320), .nC(w3128) );
	vdp_slatch g3065 (.Q(w3280), .D(w4226), .C(w3319), .nC(w3330) );
	vdp_slatch g3066 (.Q(w3274), .D(w4225), .C(w3318), .nC(w3323) );
	vdp_slatch g3067 (.Q(w4444), .D(w4281), .C(w3314), .nC(w3308) );
	vdp_slatch g3068 (.Q(w4445), .D(w4282), .C(w3127), .nC(w3309) );
	vdp_slatch g3069 (.Q(w4447), .D(w4280), .C(w3316), .nC(w3115) );
	vdp_slatch g3070 (.Q(w4446), .D(w4279), .C(w3317), .nC(w3116) );
	vdp_slatch g3071 (.Q(w4278), .D(w4276), .C(w3314), .nC(w3308) );
	vdp_slatch g3072 (.Q(w4277), .D(w4275), .C(w3127), .nC(w3309) );
	vdp_slatch g3073 (.Q(w4272), .D(w4274), .C(w3316), .nC(w3115) );
	vdp_slatch g3074 (.Q(w4271), .D(w4273), .C(w3317), .nC(w3116) );
	vdp_slatch g3075 (.Q(w4268), .D(w4270), .C(w3314), .nC(w3308) );
	vdp_slatch g3076 (.Q(w4267), .D(w4269), .C(w3127), .nC(w3309) );
	vdp_slatch g3077 (.Q(w4266), .D(w4264), .C(w3316), .nC(w3115) );
	vdp_slatch g3078 (.Q(w4263), .D(w4265), .C(w3317), .nC(w3116) );
	vdp_slatch g3079 (.Q(w4260), .D(w4262), .C(w3314), .nC(w3308) );
	vdp_slatch g3080 (.Q(w4261), .D(w4259), .C(w3127), .nC(w3309) );
	vdp_slatch g3081 (.Q(w4256), .D(w4258), .C(w3316), .nC(w3115) );
	vdp_slatch g3082 (.Q(w4257), .D(w4255), .C(w3317), .nC(w3116) );
	vdp_slatch g3083 (.Q(w4254), .D(w4252), .C(w3314), .nC(w3308) );
	vdp_slatch g3084 (.Q(w4253), .D(w4251), .C(w3127), .nC(w3309) );
	vdp_slatch g3085 (.Q(w4250), .D(w4248), .C(w3316), .nC(w3115) );
	vdp_slatch g3086 (.Q(w4249), .D(w4247), .C(w3317), .nC(w3116) );
	vdp_slatch g3087 (.Q(w4246), .D(w4244), .C(w3314), .nC(w3308) );
	vdp_slatch g3088 (.Q(w4245), .D(w4243), .C(w3127), .nC(w3309) );
	vdp_slatch g3089 (.Q(w4242), .D(w4240), .C(w3316), .nC(w3115) );
	vdp_slatch g3090 (.Q(w4241), .D(w4239), .C(w3317), .nC(w3116) );
	vdp_slatch g3091 (.Q(w4238), .D(w4236), .C(w3314), .nC(w3308) );
	vdp_slatch g3092 (.Q(w4237), .D(w4235), .C(w3127), .nC(w3309) );
	vdp_slatch g3093 (.Q(w4234), .D(w4232), .C(w3316), .nC(w3115) );
	vdp_slatch g3094 (.Q(w4233), .D(w4231), .C(w3317), .nC(w3116) );
	vdp_slatch g3095 (.Q(w4230), .D(w4228), .C(w3314), .nC(w3308) );
	vdp_slatch g3096 (.Q(w4229), .D(w4227), .C(w3127), .nC(w3309) );
	vdp_slatch g3097 (.Q(w4226), .D(w4224), .C(w3316), .nC(w3115) );
	vdp_slatch g3098 (.Q(w4225), .D(w4223), .C(w3317), .nC(w3116) );
	vdp_slatch g3099 (.Q(w4281), .D(S[3]), .C(w3079), .nC(w3113) );
	vdp_slatch g3100 (.Q(w4282), .D(S[3]), .C(w3083), .nC(w3117) );
	vdp_slatch g3101 (.Q(w4280), .D(S[3]), .C(w3086), .nC(w3114) );
	vdp_slatch g3102 (.Q(w4279), .D(S[3]), .C(w3088), .nC(w3112) );
	vdp_slatch g3103 (.Q(w4276), .D(S[7]), .C(w3079), .nC(w3113) );
	vdp_slatch g3104 (.Q(w4275), .D(S[7]), .C(w3083), .nC(w3117) );
	vdp_slatch g3105 (.Q(w4274), .D(S[7]), .C(w3086), .nC(w3114) );
	vdp_slatch g3106 (.Q(w4273), .D(S[7]), .C(w3088), .nC(w3112) );
	vdp_slatch g3107 (.Q(w4270), .D(S[2]), .C(w3079), .nC(w3113) );
	vdp_slatch g3108 (.Q(w4269), .D(S[2]), .C(w3083), .nC(w3117) );
	vdp_slatch g3109 (.Q(w4264), .D(S[2]), .C(w3086), .nC(w3114) );
	vdp_slatch g3110 (.Q(w4265), .D(S[2]), .C(w3088), .nC(w3112) );
	vdp_slatch g3111 (.Q(w4262), .D(S[6]), .C(w3079), .nC(w3113) );
	vdp_slatch g3112 (.Q(w4259), .D(S[6]), .C(w3083), .nC(w3117) );
	vdp_slatch g3113 (.Q(w4258), .D(S[6]), .C(w3086), .nC(w3114) );
	vdp_slatch g3114 (.Q(w4255), .D(S[6]), .C(w3088), .nC(w3112) );
	vdp_slatch g3115 (.Q(w4252), .D(S[1]), .C(w3079), .nC(w3113) );
	vdp_slatch g3116 (.Q(w4251), .D(S[1]), .C(w3083), .nC(w3117) );
	vdp_slatch g3117 (.Q(w4248), .D(S[1]), .C(w3086), .nC(w3114) );
	vdp_slatch g3118 (.Q(w4247), .D(S[1]), .C(w3088), .nC(w3112) );
	vdp_slatch g3119 (.Q(w4244), .D(S[5]), .C(w3079), .nC(w3113) );
	vdp_slatch g3120 (.Q(w4243), .D(S[5]), .C(w3083), .nC(w3117) );
	vdp_slatch g3121 (.Q(w4240), .D(S[5]), .C(w3086), .nC(w3114) );
	vdp_slatch g3122 (.Q(w4239), .D(S[5]), .C(w3088), .nC(w3112) );
	vdp_slatch g3123 (.Q(w4236), .D(S[0]), .C(w3079), .nC(w3113) );
	vdp_slatch g3124 (.Q(w4235), .D(S[0]), .C(w3083), .nC(w3117) );
	vdp_slatch g3125 (.Q(w4232), .D(S[0]), .C(w3086), .nC(w3114) );
	vdp_slatch g3126 (.Q(w4231), .D(S[0]), .C(w3088), .nC(w3112) );
	vdp_slatch g3127 (.Q(w4228), .D(S[4]), .C(w3079), .nC(w3113) );
	vdp_slatch g3128 (.Q(w4227), .D(S[4]), .C(w3083), .nC(w3117) );
	vdp_slatch g3129 (.Q(w4224), .D(S[4]), .C(w3086), .nC(w3114) );
	vdp_slatch g3130 (.Q(w4223), .D(S[4]), .C(w3088), .nC(w3112) );
	vdp_slatch g3131 (.Q(w4286), .D(S[3]), .C(w3080), .nC(w3105) );
	vdp_slatch g3132 (.Q(w4285), .D(S[3]), .C(w3084), .nC(w3110) );
	vdp_slatch g3133 (.Q(w4290), .D(S[3]), .C(w3085), .nC(w3111) );
	vdp_slatch g3134 (.Q(w4289), .D(S[3]), .C(w3087), .nC(w3106) );
	vdp_slatch g3135 (.Q(w4294), .D(S[7]), .C(w3080), .nC(w3105) );
	vdp_slatch g3136 (.Q(w4293), .D(S[7]), .C(w3084), .nC(w3110) );
	vdp_slatch g3137 (.Q(w4298), .D(S[7]), .C(w3085), .nC(w3111) );
	vdp_slatch g3138 (.Q(w4297), .D(S[7]), .C(w3087), .nC(w3106) );
	vdp_slatch g3139 (.Q(w4302), .D(S[2]), .C(w3080), .nC(w3105) );
	vdp_slatch g3140 (.Q(w4301), .D(S[2]), .C(w3084), .nC(w3110) );
	vdp_slatch g3141 (.Q(w4306), .D(S[2]), .C(w3085), .nC(w3111) );
	vdp_slatch g3142 (.Q(w4305), .D(S[2]), .C(w3087), .nC(w3106) );
	vdp_slatch g3143 (.Q(w4308), .D(S[6]), .C(w3080), .nC(w3105) );
	vdp_slatch g3144 (.Q(w4309), .D(S[6]), .C(w3084), .nC(w3110) );
	vdp_slatch g3145 (.Q(w4345), .D(S[6]), .C(w3085), .nC(w3111) );
	vdp_slatch g3146 (.Q(w4344), .D(S[6]), .C(w3087), .nC(w3106) );
	vdp_slatch g3147 (.Q(w4341), .D(S[1]), .C(w3080), .nC(w3105) );
	vdp_slatch g3148 (.Q(w4340), .D(S[1]), .C(w3084), .nC(w3110) );
	vdp_slatch g3149 (.Q(w4337), .D(S[1]), .C(w3085), .nC(w3111) );
	vdp_slatch g3150 (.Q(w4336), .D(S[1]), .C(w3087), .nC(w3106) );
	vdp_slatch g3151 (.Q(w4333), .D(S[5]), .C(w3080), .nC(w3105) );
	vdp_slatch g3152 (.Q(w4332), .D(S[5]), .C(w3084), .nC(w3110) );
	vdp_slatch g3153 (.Q(w4329), .D(S[5]), .C(w3085), .nC(w3111) );
	vdp_slatch g3154 (.Q(w4328), .D(S[5]), .C(w3087), .nC(w3106) );
	vdp_slatch g3155 (.Q(w4325), .D(S[0]), .C(w3080), .nC(w3105) );
	vdp_slatch g3156 (.Q(w4324), .D(S[0]), .C(w3084), .nC(w3110) );
	vdp_slatch g3157 (.Q(w4321), .D(S[0]), .C(w3085), .nC(w3111) );
	vdp_slatch g3158 (.Q(w4320), .D(S[0]), .C(w3087), .nC(w3106) );
	vdp_slatch g3159 (.Q(w4317), .D(S[4]), .C(w3080), .nC(w3105) );
	vdp_slatch g3160 (.Q(w4316), .D(S[4]), .C(w3084), .nC(w3110) );
	vdp_slatch g3161 (.Q(w4313), .D(S[4]), .C(w3085), .nC(w3111) );
	vdp_slatch g3162 (.Q(w4312), .D(S[4]), .C(w3087), .nC(w3106) );
	vdp_slatch g3163 (.Q(w4284), .D(w4286), .C(w3066), .nC(w3107) );
	vdp_slatch g3164 (.Q(w4283), .D(w4285), .C(w3069), .nC(w3108) );
	vdp_slatch g3165 (.Q(w4288), .D(w4290), .C(w3074), .nC(w3109) );
	vdp_slatch g3166 (.Q(w4287), .D(w4289), .C(w3071), .nC(w3077) );
	vdp_slatch g3167 (.Q(w4292), .D(w4294), .C(w3066), .nC(w3107) );
	vdp_slatch g3168 (.Q(w4291), .D(w4293), .C(w3069), .nC(w3108) );
	vdp_slatch g3169 (.Q(w4296), .D(w4298), .C(w3074), .nC(w3109) );
	vdp_slatch g3170 (.Q(w4295), .D(w4297), .C(w3071), .nC(w3077) );
	vdp_slatch g3171 (.Q(w4300), .D(w4302), .C(w3066), .nC(w3107) );
	vdp_slatch g3172 (.Q(w4299), .D(w4301), .C(w3069), .nC(w3108) );
	vdp_slatch g3173 (.Q(w4410), .D(w4306), .C(w3074), .nC(w3109) );
	vdp_slatch g3174 (.Q(w4304), .D(w4305), .C(w3071), .nC(w3077) );
	vdp_slatch g3175 (.Q(w4303), .D(w4308), .C(w3066), .nC(w3107) );
	vdp_slatch g3176 (.Q(w4307), .D(w4309), .C(w3069), .nC(w3108) );
	vdp_slatch g3177 (.Q(w4343), .D(w4345), .C(w3074), .nC(w3109) );
	vdp_slatch g3178 (.Q(w4342), .D(w4344), .C(w3071), .nC(w3077) );
	vdp_slatch g3179 (.Q(w4339), .D(w4341), .C(w3066), .nC(w3107) );
	vdp_slatch g3180 (.Q(w4338), .D(w4340), .C(w3069), .nC(w3108) );
	vdp_slatch g3181 (.Q(w4335), .D(w4337), .C(w3074), .nC(w3109) );
	vdp_slatch g3182 (.Q(w4334), .D(w4336), .C(w3071), .nC(w3077) );
	vdp_slatch g3183 (.Q(w4331), .D(w4333), .C(w3066), .nC(w3107) );
	vdp_slatch g3184 (.Q(w4330), .D(w4332), .C(w3069), .nC(w3108) );
	vdp_slatch g3185 (.Q(w4327), .D(w4329), .C(w3074), .nC(w3109) );
	vdp_slatch g3186 (.Q(w4326), .D(w4328), .C(w3071), .nC(w3077) );
	vdp_slatch g3187 (.D(w4325), .Q(w4323), .C(w3066), .nC(w3107) );
	vdp_slatch g3188 (.Q(w4322), .D(w4324), .C(w3069), .nC(w3108) );
	vdp_slatch g3189 (.Q(w4319), .D(w4321), .C(w3074), .nC(w3109) );
	vdp_slatch g3190 (.Q(w4318), .D(w4320), .C(w3071), .nC(w3077) );
	vdp_slatch g3191 (.Q(w4315), .D(w4317), .C(w3066), .nC(w3107) );
	vdp_slatch g3192 (.Q(w4314), .D(w4316), .C(w3069), .nC(w3108) );
	vdp_slatch g3193 (.Q(w4311), .D(w4313), .C(w3074), .nC(w3109) );
	vdp_slatch g3194 (.Q(w4310), .D(w4312), .C(w3071), .nC(w3077) );
	vdp_slatch g3195 (.Q(w3390), .D(w4284), .C(w3067), .nC(w3068) );
	vdp_slatch g3196 (.Q(w3389), .D(w4283), .C(w3075), .nC(w3076) );
	vdp_slatch g3197 (.Q(w3377), .D(w4288), .C(w3072), .nC(w3073) );
	vdp_slatch g3198 (.Q(w3375), .D(w4287), .C(w3065), .nC(w3064) );
	vdp_slatch g3199 (.Q(w3388), .D(w4292), .C(w3067), .nC(w3068) );
	vdp_slatch g3200 (.Q(w3396), .D(w4291), .C(w3075), .nC(w3076) );
	vdp_slatch g3201 (.D(w4296), .C(w3072), .nC(w3073), .Q(w3386) );
	vdp_slatch g3202 (.Q(w3374), .D(w4295), .C(w3065), .nC(w3064) );
	vdp_slatch g3203 (.Q(w3385), .D(w4300), .C(w3067), .nC(w3068) );
	vdp_slatch g3204 (.Q(w3384), .D(w4299), .C(w3075), .nC(w3076) );
	vdp_slatch g3205 (.Q(w3383), .D(w4410), .C(w3072), .nC(w3073) );
	vdp_slatch g3206 (.Q(w3382), .D(w4304), .C(w3065), .nC(w3064) );
	vdp_slatch g3207 (.Q(w3381), .D(w4303), .C(w3067), .nC(w3068) );
	vdp_slatch g3208 (.Q(w3380), .D(w4307), .C(w3075), .nC(w3076) );
	vdp_slatch g3209 (.Q(w3379), .D(w4343), .C(w3072), .nC(w3073) );
	vdp_slatch g3210 (.Q(w3378), .D(w4342), .C(w3065), .nC(w3064) );
	vdp_slatch g3211 (.Q(w3370), .D(w4339), .C(w3067), .nC(w3068) );
	vdp_slatch g3212 (.Q(w3417), .D(w4338), .C(w3075), .nC(w3076) );
	vdp_slatch g3213 (.Q(w3371), .D(w4335), .C(w3072), .nC(w3073) );
	vdp_slatch g3214 (.Q(w3372), .D(w4334), .C(w3065), .nC(w3064) );
	vdp_slatch g3215 (.Q(w3421), .D(w4331), .C(w3067), .nC(w3068) );
	vdp_slatch g3216 (.Q(w3430), .D(w4330), .C(w3075), .nC(w3076) );
	vdp_slatch g3217 (.Q(w3422), .D(w4327), .C(w3072), .nC(w3073) );
	vdp_slatch g3218 (.Q(w3429), .D(w4326), .nC(w3064), .C(w3065) );
	vdp_slatch g3219 (.Q(w3428), .D(w4323), .C(w3067), .nC(w3068) );
	vdp_slatch g3220 (.Q(w3427), .D(w4322), .C(w3075), .nC(w3076) );
	vdp_slatch g3221 (.Q(w3423), .D(w4319), .C(w3072), .nC(w3073) );
	vdp_slatch g3222 (.Q(w3426), .D(w4318), .C(w3065), .nC(w3064) );
	vdp_slatch g3223 (.Q(w3425), .D(w4315), .C(w3067), .nC(w3068) );
	vdp_slatch g3224 (.Q(w3424), .D(w4314), .C(w3075), .nC(w3070) );
	vdp_slatch g3225 (.Q(w3376), .D(w4311), .C(w3072), .nC(w3073) );
	vdp_slatch g3226 (.Q(w3373), .D(w4310), .C(w3065), .nC(w3064) );
	vdp_slatch g3227 (.Q(w3409), .D(w4349), .nC(w3471), .C(w3470) );
	vdp_slatch g3228 (.Q(w3518), .D(w4348), .nC(w3474), .C(w3475) );
	vdp_slatch g3229 (.Q(w3411), .D(w4353), .nC(w3473), .C(w3472) );
	vdp_slatch g3230 (.Q(w3410), .D(w4352), .nC(w3477), .C(w3476) );
	vdp_slatch g3231 (.Q(w3517), .D(w4357), .nC(w3471), .C(w3470) );
	vdp_slatch g3232 (.Q(w3521), .D(w4356), .nC(w3474), .C(w3475) );
	vdp_slatch g3233 (.Q(w3520), .D(w4361), .nC(w3473), .C(w3472) );
	vdp_slatch g3234 (.Q(w3519), .D(w4360), .nC(w3477), .C(w3476) );
	vdp_slatch g3235 (.Q(w3412), .D(w4365), .nC(w3471), .C(w3470) );
	vdp_slatch g3236 (.Q(w3522), .D(w4364), .nC(w3474), .C(w3475) );
	vdp_slatch g3237 (.Q(w3516), .D(w4369), .nC(w3473), .C(w3472) );
	vdp_slatch g3238 (.Q(w3523), .D(w4368), .nC(w3477), .C(w3476) );
	vdp_slatch g3239 (.Q(w3524), .D(w4373), .nC(w3471), .C(w3470) );
	vdp_slatch g3240 (.Q(w3525), .D(w4372), .nC(w3474), .C(w3475) );
	vdp_slatch g3241 (.Q(w3413), .D(w4377), .nC(w3473), .C(w3472) );
	vdp_slatch g3242 (.Q(w3414), .D(w4376), .nC(w3477), .C(w3476) );
	vdp_slatch g3243 (.Q(w3508), .D(w4381), .nC(w3471), .C(w3470) );
	vdp_slatch g3244 (.Q(w3509), .D(w4380), .nC(w3474), .C(w3475) );
	vdp_slatch g3245 (.Q(w3510), .D(w4385), .nC(w3473), .C(w3472) );
	vdp_slatch g3246 (.Q(w3511), .D(w4384), .nC(w3477), .C(w3476) );
	vdp_slatch g3247 (.Q(w3512), .D(w4389), .nC(w3471), .C(w3470) );
	vdp_slatch g3248 (.Q(w3513), .D(w4388), .nC(w3474), .C(w3475) );
	vdp_slatch g3249 (.Q(w3514), .D(w4393), .nC(w3473), .C(w3472) );
	vdp_slatch g3250 (.Q(w3515), .D(w4392), .nC(w3477), .C(w3476) );
	vdp_slatch g3251 (.Q(w3507), .D(w4397), .nC(w3471), .C(w3470) );
	vdp_slatch g3252 (.Q(w3506), .D(w4396), .nC(w3474), .C(w3475) );
	vdp_slatch g3253 (.Q(w3505), .D(w4401), .nC(w3473), .C(w3472) );
	vdp_slatch g3254 (.Q(w3504), .D(w4400), .nC(w3477), .C(w3476) );
	vdp_slatch g3255 (.Q(w3503), .D(w4405), .nC(w3471), .C(w3470) );
	vdp_slatch g3256 (.Q(w3502), .D(w4404), .nC(w3474), .C(w3475) );
	vdp_slatch g3257 (.Q(w3500), .D(w4409), .nC(w3473), .C(w3472) );
	vdp_slatch g3258 (.Q(w3501), .D(w4408), .nC(w3477), .C(w3476) );
	vdp_slatch g3259 (.Q(w4349), .D(w4347), .C(w3435), .nC(w3469) );
	vdp_slatch g3260 (.Q(w4348), .D(w4346), .C(w3461), .nC(w3463) );
	vdp_slatch g3261 (.Q(w4353), .D(w4351), .C(w3436), .nC(w3464) );
	vdp_slatch g3262 (.Q(w4352), .D(w4350), .C(w3468), .nC(w3467) );
	vdp_slatch g3263 (.Q(w4357), .D(w4355), .C(w3435), .nC(w3469) );
	vdp_slatch g3264 (.Q(w4356), .D(w4354), .C(w3461), .nC(w3463) );
	vdp_slatch g3265 (.Q(w4361), .D(w4359), .C(w3436), .nC(w3464) );
	vdp_slatch g3266 (.Q(w4360), .D(w4358), .C(w3468), .nC(w3467) );
	vdp_slatch g3267 (.Q(w4365), .D(w4363), .C(w3435), .nC(w3469) );
	vdp_slatch g3268 (.Q(w4364), .D(w4362), .C(w3461), .nC(w3463) );
	vdp_slatch g3269 (.Q(w4369), .D(w4367), .C(w3436), .nC(w3464) );
	vdp_slatch g3270 (.Q(w4368), .D(w4366), .C(w3468), .nC(w3467) );
	vdp_slatch g3271 (.Q(w4373), .D(w4371), .C(w3435), .nC(w3469) );
	vdp_slatch g3272 (.Q(w4372), .D(w4370), .C(w3461), .nC(w3463) );
	vdp_slatch g3273 (.Q(w4377), .D(w4375), .C(w3436), .nC(w3464) );
	vdp_slatch g3274 (.Q(w4376), .D(w4374), .C(w3468), .nC(w3467) );
	vdp_slatch g3275 (.Q(w4381), .D(w4379), .C(w3435), .nC(w3469) );
	vdp_slatch g3276 (.Q(w4380), .D(w4378), .C(w3461), .nC(w3463) );
	vdp_slatch g3277 (.Q(w4385), .D(w4383), .C(w3436), .nC(w3464) );
	vdp_slatch g3278 (.Q(w4384), .D(w4382), .C(w3468), .nC(w3467) );
	vdp_slatch g3279 (.Q(w4389), .D(w4387), .C(w3435), .nC(w3469) );
	vdp_slatch g3280 (.Q(w4388), .D(w4386), .C(w3461), .nC(w3463) );
	vdp_slatch g3281 (.Q(w4393), .D(w4391), .C(w3436), .nC(w3464) );
	vdp_slatch g3282 (.Q(w4392), .D(w4390), .C(w3468), .nC(w3467) );
	vdp_slatch g3283 (.Q(w4397), .D(w4395), .C(w3435), .nC(w3469) );
	vdp_slatch g3284 (.Q(w4396), .D(w4394), .C(w3461), .nC(w3463) );
	vdp_slatch g3285 (.Q(w4401), .D(w4399), .C(w3436), .nC(w3464) );
	vdp_slatch g3286 (.Q(w4400), .D(w4398), .C(w3468), .nC(w3467) );
	vdp_slatch g3287 (.Q(w4405), .D(w4403), .C(w3435), .nC(w3469) );
	vdp_slatch g3288 (.Q(w4404), .D(w4402), .C(w3461), .nC(w3463) );
	vdp_slatch g3289 (.Q(w4409), .D(w4407), .C(w3436), .nC(w3464) );
	vdp_slatch g3290 (.Q(w4408), .D(w4406), .C(w3468), .nC(w3467) );
	vdp_slatch g3291 (.Q(w4347), .D(S[3]), .nC(w3462), .C(w3490) );
	vdp_slatch g3292 (.Q(w4346), .D(S[3]), .nC(w3478), .C(w3491) );
	vdp_slatch g3293 (.Q(w4351), .D(S[3]), .nC(w3465), .C(w3489) );
	vdp_slatch g3294 (.Q(w4350), .D(S[3]), .nC(w3466), .C(w3488) );
	vdp_slatch g3295 (.Q(w4355), .D(S[7]), .nC(w3462), .C(w3490) );
	vdp_slatch g3296 (.Q(w4354), .D(S[7]), .nC(w3478), .C(w3491) );
	vdp_slatch g3297 (.Q(w4359), .D(S[7]), .nC(w3465), .C(w3489) );
	vdp_slatch g3298 (.Q(w4358), .D(S[7]), .nC(w3466), .C(w3488) );
	vdp_slatch g3299 (.Q(w4363), .D(S[2]), .nC(w3462), .C(w3490) );
	vdp_slatch g3300 (.Q(w4362), .D(S[2]), .nC(w3478), .C(w3491) );
	vdp_slatch g3301 (.Q(w4367), .D(S[2]), .nC(w3465), .C(w3489) );
	vdp_slatch g3302 (.Q(w4366), .D(S[2]), .nC(w3466), .C(w3488) );
	vdp_slatch g3303 (.Q(w4371), .D(S[6]), .nC(w3462), .C(w3490) );
	vdp_slatch g3304 (.Q(w4370), .D(S[6]), .nC(w3478), .C(w3491) );
	vdp_slatch g3305 (.Q(w4375), .D(S[6]), .nC(w3465), .C(w3489) );
	vdp_slatch g3306 (.Q(w4374), .D(S[6]), .nC(w3466), .C(w3488) );
	vdp_slatch g3307 (.Q(w4379), .D(S[1]), .nC(w3462), .C(w3490) );
	vdp_slatch g3308 (.Q(w4378), .D(S[1]), .nC(w3478), .C(w3491) );
	vdp_slatch g3309 (.Q(w4383), .D(S[1]), .nC(w3465), .C(w3489) );
	vdp_slatch g3310 (.Q(w4382), .D(S[1]), .nC(w3466), .C(w3488) );
	vdp_slatch g3311 (.Q(w4387), .D(S[5]), .nC(w3462), .C(w3490) );
	vdp_slatch g3312 (.Q(w4386), .D(S[5]), .nC(w3478), .C(w3491) );
	vdp_slatch g3313 (.Q(w4391), .D(S[5]), .nC(w3465), .C(w3489) );
	vdp_slatch g3314 (.Q(w4390), .D(S[5]), .nC(w3466), .C(w3488) );
	vdp_slatch g3315 (.Q(w4395), .D(S[0]), .nC(w3462), .C(w3490) );
	vdp_slatch g3316 (.Q(w4394), .D(S[0]), .nC(w3478), .C(w3491) );
	vdp_slatch g3317 (.Q(w4399), .D(S[0]), .nC(w3465), .C(w3489) );
	vdp_slatch g3318 (.Q(w4398), .D(S[0]), .nC(w3466), .C(w3488) );
	vdp_slatch g3319 (.Q(w4403), .D(S[4]), .nC(w3462), .C(w3490) );
	vdp_slatch g3320 (.Q(w4402), .D(S[4]), .nC(w3478), .C(w3491) );
	vdp_slatch g3321 (.Q(w4407), .D(S[4]), .nC(w3465), .C(w3489) );
	vdp_slatch g3322 (.Q(w4406), .D(S[4]), .nC(w3466), .C(w3488) );
	vdp_aon2*8 g3323 (.Z(w4045), .A1(w3205), .B1(w3204), .C1(w3203), .D2(w3202), .A2(w3250), .B2(w3251), .C2(w3256), .D1(w3255), .E2(w3253), .F1(w3254), .E1(w3201), .F2(w3200), .G1(w3199), .H2(w3198), .G2(w3258), .H1(w3248) );
	vdp_aon2*8 g3324 (.Z(w3230), .A1(w3324), .B1(w3251), .C1(w3326), .D2(w3255), .A2(w3250), .B2(w3325), .C2(w3256), .D1(w3327), .E2(w3253), .F1(w3254), .E1(w3328), .F2(w3329), .G1(w3334), .H2(w3335), .G2(w3258), .H1(w3248) );
	vdp_aon2*8 g3325 (.Z(w3233), .A1(w3197), .B1(w3210), .C1(w3214), .D2(w3213), .A2(w3250), .B2(w3251), .C2(w3256), .D1(w3255), .E2(w3253), .F1(w3254), .E1(w3212), .F2(w3208), .G1(w3209), .H2(w3211), .G2(w3258), .H1(w3248) );
	vdp_aon2*8 g3326 (.Z(w3234), .A1(w3336), .B1(w3251), .C1(w3338), .D2(w3255), .A2(w3250), .B2(w3337), .C2(w3256), .D1(w3333), .E2(w3253), .F1(w3254), .E1(w3339), .F2(w3340), .G1(w3341), .H2(w3342), .G2(w3258), .H1(w3248) );
	vdp_aon2*8 g3327 (.Z(w3232), .A1(w3268), .B1(w3251), .C1(w3270), .D2(w3271), .A2(w3250), .B2(w4046), .C2(w3256), .D1(w3255), .E2(w3253), .F1(w3254), .E1(w3343), .F2(w3269), .G1(w3249), .H2(w3272), .G2(w3258), .H1(w3248) );
	vdp_aon2*8 g3328 (.Z(w3235), .A1(w3275), .B1(w3251), .C1(w3282), .D2(w3281), .A2(w3250), .B2(w3283), .C2(w3256), .D1(w3255), .E2(w3253), .F1(w3254), .E1(w3279), .F2(w3273), .G1(w3280), .G2(w3258), .H1(w3248), .H2(w3274) );
	vdp_aon2*8 g3329 (.Z(w3231), .A1(w3215), .B1(w3216), .C1(w3218), .D2(w3217), .A2(w3250), .B2(w3251), .C2(w3256), .D1(w3255), .E2(w3253), .F1(w3254), .E1(w3260), .F2(w3261), .G1(w3257), .H2(w3252), .G2(w3258), .H1(w3248) );
	vdp_aon2*8 g3330 (.Z(w3236), .A1(w3264), .B1(w3263), .C1(w3262), .D2(w3259), .A2(w3250), .B2(w3251), .C2(w3256), .D1(w3255), .E2(w3253), .F1(w3254), .E1(w3245), .F2(w3244), .G1(w3246), .H2(w3247), .G2(w3258), .H1(w3248) );
	vdp_aon2*8 g3331 (.A1(w3390), .B1(w3389), .C1(w3377), .D2(w3375), .A2(w3408), .B2(w3407), .C2(w3406), .D1(w3405), .E2(w3404), .F1(w3403), .E1(w3388), .F2(w3387), .G1(w3386), .H2(w3374), .G2(w3401), .H1(w3402), .Z(w3420) );
	vdp_aon2*8 g3332 (.Z(w3448), .A1(w3385), .B1(w3384), .C1(w3383), .D2(w3382), .A2(w3408), .B2(w3407), .C2(w3406), .D1(w3405), .E2(w3404), .F1(w3403), .E1(w3381), .F2(w3380), .G1(w3379), .H2(w3378), .G2(w3401), .H1(w3402) );
	vdp_aon2*8 g3333 (.Z(w3419), .A1(w3377), .B1(w3386), .C1(w3383), .D2(w3379), .A2(w3403), .B2(w3402), .C2(w3407), .D1(w3405), .E2(w3404), .F1(w3401), .E1(w3371), .F2(w3422), .G1(w3423), .H2(w3376), .G2(w3408), .H1(w3406) );
	vdp_aon2*8 g3334 (.Z(w3451), .A1(w3370), .B1(w3417), .C1(w3371), .D2(w3372), .A2(w3408), .B2(w3407), .C2(w3406), .D1(w3405), .E2(w3404), .F1(w3403), .E1(w3421), .F2(w3430), .G1(w3422), .H2(w3429), .G2(w3401), .H1(w3402) );
	vdp_aon2*8 g3335 (.Z(w3418), .A1(w3428), .B1(w3427), .C1(w3423), .D2(w3426), .A2(w3408), .B2(w3407), .C2(w3406), .D1(w3405), .E2(w3404), .F1(w3403), .E1(w3425), .F2(w3424), .G1(w3376), .H2(w3373), .G2(w3401), .H1(w3402) );
	vdp_aon2*8 g3336 (.Z(w3453), .A1(w3507), .B1(w3407), .C1(w3505), .D2(w3405), .A2(w3408), .B2(w3506), .C2(w3406), .D1(w3504), .E2(w3404), .F1(w3403), .E1(w3503), .F2(w3502), .G1(w3500), .H2(w3501), .G2(w3401), .H1(w3402) );
	vdp_aon2*8 g3337 (.Z(w3454), .A1(w3508), .B1(w3407), .C1(w3510), .D2(w3405), .A2(w3408), .B2(w3509), .C2(w3406), .D1(w3511), .E2(w3404), .F1(w3403), .E1(w3512), .F2(w3513), .G1(w3514), .H2(w3515), .G2(w3401), .H1(w3402) );
	vdp_aon2*8 g3338 (.Z(w3452), .A1(w3375), .B1(w3374), .C1(w3382), .D2(w3378), .A2(w3403), .B2(w3402), .C2(w3407), .D1(w3405), .E2(w3404), .F1(w3401), .E1(w3372), .F2(w3429), .G1(w3426), .H2(w3373), .G2(w3408), .H1(w3406) );
	vdp_aon2*8 g3339 (.Z(w3447), .A1(w3410), .B1(w3402), .C1(w3523), .D2(w3405), .A2(w3403), .B2(w3519), .C2(w3407), .D1(w3414), .E2(w3404), .F1(w3401), .E1(w3511), .F2(w3515), .G1(w3504), .H2(w3501), .G2(w3408), .H1(w3406) );
	vdp_aon2*8 g3340 (.Z(w3450), .A1(w3411), .B1(w3402), .C1(w3516), .D2(w3405), .A2(w3403), .B2(w3520), .C2(w3407), .D1(w3413), .E2(w3404), .F1(w3401), .E1(w3510), .F2(w3514), .G1(w3505), .H2(w3500), .G2(w3408), .H1(w3406) );
	vdp_aon2*8 g3341 (.Z(w3449), .A1(w3412), .B1(w3407), .C1(w3516), .D2(w3405), .A2(w3408), .B2(w3522), .C2(w3406), .D1(w3523), .E2(w3404), .F1(w3403), .E1(w3524), .F2(w3525), .G1(w3413), .H2(w3414), .G2(w3401), .H1(w3402) );
	vdp_aon2*8 g3342 (.A1(w3409), .B1(w3407), .C1(w3411), .D2(w3405), .A2(w3408), .B2(w3518), .C2(w3406), .D1(w3410), .E2(w3404), .F1(w3403), .E1(w3517), .F2(w3521), .G1(w3520), .H2(w3519), .G2(w3401), .H1(w3402), .Z(w3455) );
	vdp_sr_bit g3343 (.Q(w3398), .D(w3553), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3344 (.Q(w3553), .D(w3457), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3345 (.Q(w3458), .D(w3554), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3346 (.Q(w3554), .D(w3460), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3347 (.Q(w3459), .D(w3434), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3348 (.Q(w4076), .D(w3459), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3349 (.Q(w3538), .D(w3456), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3350 (.Q(w3433), .D(w3538), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3351 (.Q(w4078), .D(w3443), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3352 (.Q(w3432), .D(w4078), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3353 (.Q(w3431), .D(w3399), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3354 (.Q(w3399), .D(w3442), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3355 (.Q(w2843), .D(w3444), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3356 (.Q(w3539), .D(w2843), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3357 (.Q(w3221), .D(w3240), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3358 (.Q(w3223), .D(w3221), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3359 (.Q(w3227), .D(w3222), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3360 (.Q(w3222), .D(w3239), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3361 (.Q(w3238), .D(w3219), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3362 (.Q(w3219), .D(w3241), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3363 (.Q(w3220), .D(w3237), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3364 (.Q(w3229), .D(w3220), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3365 (.Q(w3307), .D(w2842), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3366 (.Q(w2842), .D(w3292), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3367 (.Q(w4057), .D(w3242), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3368 (.Q(w3228), .D(w4057), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3369 (.Q(w4056), .D(w3293), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3370 (.Q(w3226), .D(w4056), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3371 (.Q(w3153), .D(VRAMA[1]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3372 (.Q(w3185), .D(VRAMA[2]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3373 (.Q(w3187), .D(VRAMA[3]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3374 (.Q(w3188), .D(VRAMA[4]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3375 (.Q(w3189), .D(VRAMA[5]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3376 (.Q(w3190), .D(VRAMA[6]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3377 (.Q(w4054), .D(w3176), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3378 (.Q(w3540), .D(w4054), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3379 (.Q(w3175), .D(w3541), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3380 (.Q(w3541), .D(w3540), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_dlatch_inv g3381 (.nQ(w3176), .D(w3141), .C(DCLK1), .nC(nDCLK1) );
	vdp_slatch g3382 (.Q(w3301), .D(w4411), .C(w3294), .nC(w3052) );
	vdp_slatch g3383 (.Q(w3300), .D(w4412), .C(w3294), .nC(w3052) );
	vdp_slatch g3384 (.Q(w3299), .D(w4413), .C(w3294), .nC(w3052) );
	vdp_slatch g3385 (.Q(w3298), .D(w4414), .C(w3294), .nC(w3052) );
	vdp_slatch g3386 (.Q(w3297), .D(w4415), .C(w3294), .nC(w3052) );
	vdp_slatch g3387 (.Q(w3296), .D(w4416), .C(w3294), .nC(w3052) );
	vdp_slatch g3388 (.Q(w3295), .D(w4418), .C(w3294), .nC(w3052) );
	vdp_slatch g3389 (.Q(w3053), .D(w4417), .C(w3294), .nC(w3052) );
	vdp_slatch g3390 (.Q(w4411), .D(w3121), .C(w3315), .nC(w3346) );
	vdp_slatch g3391 (.Q(w4412), .D(w3095), .C(w3315), .nC(w3346) );
	vdp_slatch g3392 (.Q(w4413), .D(w3097), .C(w3315), .nC(w3346) );
	vdp_slatch g3393 (.Q(w4414), .D(w3098), .C(w3315), .nC(w3346) );
	vdp_slatch g3394 (.Q(w4415), .D(w3099), .C(w3315), .nC(w3346) );
	vdp_slatch g3395 (.Q(w4416), .D(w3122), .C(w3315), .nC(w3346) );
	vdp_slatch g3396 (.Q(w4418), .D(w3126), .C(w3315), .nC(w3346) );
	vdp_slatch g3397 (.Q(w4417), .D(w3125), .C(w3315), .nC(w3346) );
	vdp_slatch g3398 (.Q(w4419), .D(w3060), .C(w3062), .nC(w3061) );
	vdp_slatch g3399 (.Q(w4420), .D(w3094), .C(w3062), .nC(w3061) );
	vdp_slatch g3400 (.Q(w4421), .D(w3059), .C(w3062), .nC(w3061) );
	vdp_slatch g3401 (.Q(w4422), .D(w4108), .C(w3062), .nC(w3061) );
	vdp_slatch g3402 (.Q(w4423), .D(w3549), .C(w3062), .nC(w3061) );
	vdp_slatch g3403 (.Q(w4424), .D(w3101), .C(w3062), .nC(w3061) );
	vdp_slatch g3404 (.Q(w4425), .D(w3056), .C(w3062), .nC(w3061) );
	vdp_slatch g3405 (.Q(w4426), .D(w3102), .C(w3062), .nC(w3061) );
	vdp_slatch g3406 (.Q(w3355), .D(w4419), .C(w3063), .nC(w3348) );
	vdp_slatch g3407 (.Q(w3354), .D(w4420), .C(w3063), .nC(w3348) );
	vdp_slatch g3408 (.Q(w3353), .D(w4421), .C(w3063), .nC(w3348) );
	vdp_slatch g3409 (.Q(w3352), .D(w4422), .C(w3063), .nC(w3348) );
	vdp_slatch g3410 (.Q(w3351), .D(w4423), .C(w3063), .nC(w3348) );
	vdp_slatch g3411 (.Q(w3350), .D(w4424), .C(w3063), .nC(w3348) );
	vdp_slatch g3412 (.Q(w3349), .D(w4425), .C(w3063), .nC(w3348) );
	vdp_slatch g3413 (.Q(w4452), .D(w4426), .C(w3063), .nC(w3348) );
	vdp_slatch g3414 (.Q(w3492), .D(w3486), .C(w3173), .nC(w3483) );
	vdp_slatch g3415 (.Q(w3485), .D(w3180), .C(w3173), .nC(w3483) );
	vdp_slatch g3416 (.Q(w3887), .D(w3484), .C(w3173), .nC(w3483) );
	vdp_slatch g3417 (.Q(w3479), .D(w3482), .C(w3173), .nC(w3483) );
	vdp_slatch g3418 (.Q(w3060), .D(w3121), .C(w3124), .nC(w3123) );
	vdp_slatch g3419 (.Q(w3094), .D(w3095), .C(w3124), .nC(w3123) );
	vdp_slatch g3420 (.Q(w3059), .D(w3097), .C(w3124), .nC(w3123) );
	vdp_slatch g3421 (.Q(w4108), .D(w3098), .C(w3124), .nC(w3123) );
	vdp_slatch g3422 (.Q(w3549), .D(w3099), .C(w3124), .nC(w3123) );
	vdp_slatch g3423 (.Q(w3101), .D(w3122), .C(w3124), .nC(w3123) );
	vdp_slatch g3424 (.Q(w3056), .D(w3126), .C(w3124), .nC(w3123) );
	vdp_slatch g3425 (.Q(w3102), .D(w3125), .C(w3124), .nC(w3123) );
	vdp_cnt_bit_load g3426 (.D(w3484), .nL(w3145), .L(w3142), .R(1'b0), .Q(w3144), .CI(w3545), .CO(w3546), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3427 (.D(w3180), .nL(w3145), .L(w3142), .R(1'b0), .Q(w4043), .CI(w3546), .CO(w3547), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3428 (.D(w3146), .nL(w3145), .L(w3142), .R(1'b0), .Q(w3130), .CI(w3547), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3429 (.CO(w3545), .CI(1'b1), .D(w3482), .nL(w3145), .L(w3142), .R(1'b0), .Q(w3140), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3430 (.CO(w3544), .CI(1'b1), .D(w3479), .nL(w3481), .L(w3172), .R(1'b0), .Q(w3499), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3431 (.CO(w3543), .CI(w3544), .D(w3887), .nL(w3481), .L(w3172), .R(1'b0), .Q(w3445), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3432 (.CO(w3542), .CI(w3543), .D(w3485), .nL(w3481), .L(w3172), .R(1'b0), .Q(w3487), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3433 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .CI(w3542), .D(w3492), .nL(w3481), .L(w3172), .R(1'b0), .Q(w3397) );
	vdp_xor g3434 (.Z(w3284), .B(w4043), .A(w3139) );
	vdp_xor g3435 (.B(w3144), .A(w3139), .Z(w3131) );
	vdp_xor g3436 (.Z(w3287), .B(w3140), .A(w3139) );
	vdp_sr_bit g3437 (.Q(w3138), .D(w4052), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3438 (.Q(w4051), .D(w3138), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3439 (.Q(w3306), .D(w4051), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3440 (.Q(w4060), .D(w3548), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3441 (.Q(w3548), .D(w4061), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3442 (.Q(w4061), .D(w4062), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3443 (.Q(w3058), .D(w3057), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3444 (.Q(w3057), .D(w3055), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3445 (.Q(w3055), .D(w3054), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3446 (.Q(w4064), .D(w4065), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3447 (.Q(w4031), .D(w4064), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3448 (.Q(w4063), .D(w4031), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3449 (.Q(w4068), .D(w4067), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3450 (.Q(w4069), .D(w4068), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3451 (.Q(w4066), .D(w4069), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3452 (.Q(w3152), .D(w4066), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3453 (.Q(w4151), .D(w4152), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3454 (.Q(w4152), .D(w4071), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_xor g3455 (.Z(w3358), .A(w3441), .B(w3487) );
	vdp_xor g3456 (.Z(w3363), .A(w3441), .B(w3498) );
	vdp_xor g3457 (.Z(w3357), .A(w3441), .B(w3499) );
	vdp_dlatch_inv g3458 (.nQ(w4050), .D(w4049), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g3459 (.nQ(w3054), .D(w3100), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g3460 (.nQ(w4065), .D(w3050), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g3461 (.nQ(w3497), .D(w4072), .nC(nHCLK1), .C(HCLK1) );
	vdp_xor g3462 (.Z(w3498), .A(w3445), .B(M5) );
	vdp_sr_bit g3463 (.Q(w3551), .D(w3446), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_dlatch_inv g3464 (.nQ(w4067), .D(w3150), .nC(nDCLK1), .C(DCLK1) );
	vdp_comp_strong g3465 (.Z(w3067), .nZ(w3068), .A(w3347) );
	vdp_comp_strong g3466 (.Z(w3075), .nZ(w3076), .A(w3347) );
	vdp_comp_strong g3467 (.Z(w3072), .nZ(w3073), .A(w3347) );
	vdp_comp_strong g3468 (.Z(w3065), .nZ(w3064), .A(w3347) );
	vdp_comp_strong g3469 (.Z(w3066), .nZ(w3107), .A(w3103) );
	vdp_comp_strong g3470 (.Z(w3069), .nZ(w3108), .A(w3103) );
	vdp_comp_strong g3471 (.Z(w3074), .nZ(w3109), .A(w3103) );
	vdp_comp_strong g3472 (.Z(w3071), .nZ(w3077), .A(w3103) );
	vdp_comp_strong g3473 (.Z(w3080), .nZ(w3105), .A(w3104) );
	vdp_comp_strong g3474 (.Z(w3084), .nZ(w3110), .A(w3416) );
	vdp_comp_strong g3475 (.Z(w3085), .nZ(w3111), .A(w3415) );
	vdp_comp_strong g3476 (.Z(w3087), .nZ(w3106), .A(w3096) );
	vdp_comp_strong g3477 (.Z(w3079), .nZ(w3113), .A(w4059) );
	vdp_comp_strong g3478 (.Z(w3083), .nZ(w3117), .A(w3118) );
	vdp_comp_strong g3479 (.Z(w3086), .nZ(w3114), .A(w3120) );
	vdp_comp_strong g3480 (.Z(w3088), .nZ(w3112), .A(w3119) );
	vdp_comp_strong g3481 (.Z(w3314), .nZ(w3308), .A(w3051) );
	vdp_comp_strong g3482 (.Z(w3127), .nZ(w3309), .A(w3051) );
	vdp_comp_strong g3483 (.Z(w3316), .nZ(w3115), .A(w3051) );
	vdp_comp_strong g3484 (.Z(w3317), .nZ(w3116), .A(w3051) );
	vdp_comp_strong g3485 (.Z(w3321), .nZ(w3322), .A(w3129) );
	vdp_comp_strong g3486 (.Z(w3320), .nZ(w3128), .A(w3129) );
	vdp_comp_strong g3487 (.Z(w3319), .nZ(w3330), .A(w3129) );
	vdp_comp_strong g3488 (.Z(w3318), .nZ(w3323), .A(w3129) );
	vdp_comp_strong g3489 (.Z(w3170), .nZ(w3196), .A(w3129) );
	vdp_comp_strong g3490 (.Z(w3149), .nZ(w3206), .A(w3129) );
	vdp_comp_strong g3491 (.Z(w3161), .nZ(w3207), .A(w3129) );
	vdp_comp_strong g3492 (.Z(w3162), .nZ(w3136), .A(w3129) );
	vdp_comp_strong g3493 (.Z(w3148), .nZ(w3165), .A(w3051) );
	vdp_comp_strong g3494 (.Z(w3166), .nZ(w3157), .A(w3051) );
	vdp_comp_strong g3495 (.Z(w3167), .nZ(w3155), .A(w3051) );
	vdp_comp_strong g3496 (.Z(w3163), .nZ(w3164), .A(w3051) );
	vdp_comp_strong g3497 (.Z(w3178), .nZ(w3168), .A(w3179) );
	vdp_comp_strong g3498 (.Z(w3159), .nZ(w3158), .A(w3181) );
	vdp_comp_strong g3499 (.Z(w3160), .nZ(w3156), .A(w3182) );
	vdp_comp_strong g3500 (.Z(w3177), .nZ(w3169), .A(w3183) );
	vdp_comp_strong g3501 (.Z(w3490), .nZ(w3462), .A(w3304) );
	vdp_comp_strong g3502 (.Z(w3491), .nZ(w3478), .A(w3493) );
	vdp_comp_strong g3503 (.Z(w3489), .nZ(w3465), .A(w3494) );
	vdp_comp_strong g3504 (.Z(w3488), .nZ(w3466), .A(w3495) );
	vdp_comp_strong g3505 (.Z(w3435), .nZ(w3469), .A(w3103) );
	vdp_comp_strong g3506 (.Z(w3461), .nZ(w3463), .A(w3103) );
	vdp_comp_strong g3507 (.Z(w3436), .nZ(w3464), .A(w3103) );
	vdp_comp_strong g3508 (.Z(w3468), .nZ(w3467), .A(w3103) );
	vdp_comp_strong g3509 (.Z(w3470), .nZ(w3471), .A(w3347) );
	vdp_comp_strong g3510 (.Z(w3475), .nZ(w3474), .A(w3347) );
	vdp_comp_strong g3511 (.Z(w3472), .nZ(w3473), .A(w3347) );
	vdp_comp_strong g3512 (.Z(w3476), .nZ(w3477), .A(w3347) );
	vdp_not g3513 (.nZ(w3146), .A(w3486) );
	vdp_not g3514 (.nZ(w4052), .A(w3265) );
	vdp_not g3515 (.nZ(w3267), .A(w103) );
	vdp_not g3516 (.nZ(w3266), .A(w441) );
	vdp_not g3517 (.nZ(w3132), .A(w3266) );
	vdp_comp_strong g3518 (.Z(w3294), .nZ(w3052), .A(w3129) );
	vdp_comp_strong g3519 (.Z(w3315), .nZ(w3346), .A(w3051) );
	vdp_comp_strong g3520 (.Z(w3124), .nZ(w3123), .A(w3304) );
	vdp_comp_strong g3521 (.Z(w3063), .nZ(w3348), .A(w3347) );
	vdp_comp_strong g3522 (.Z(w3062), .nZ(w3061), .A(w3103) );
	vdp_comp_strong g3523 (.Z(w3173), .nZ(w3483), .A(w3551) );
	vdp_not g3524 (.nZ(w3364), .A(w3357) );
	vdp_not g3525 (.nZ(w3356), .A(w3363) );
	vdp_not g3526 (.nZ(w3367), .A(w3358) );
	vdp_nand3 g3527 (.Z(w3361), .A(w3367), .B(w3363), .C(w3357) );
	vdp_not g3528 (.nZ(w3407), .A(w3360) );
	vdp_nand3 g3529 (.Z(w3360), .A(w3358), .B(w3356), .C(w3357) );
	vdp_nand3 g3530 (.Z(w3359), .A(w3358), .B(w3363), .C(w3357) );
	vdp_nand3 g3531 (.Z(w3365), .A(w3358), .B(w3363), .C(w3364) );
	vdp_nand3 g3532 (.Z(w3362), .A(w3367), .B(w3356), .C(w3357) );
	vdp_nand3 g3533 (.Z(w3368), .A(w3367), .B(w3363), .C(w3364) );
	vdp_nand3 g3534 (.Z(w3366), .A(w3358), .B(w3356), .C(w3364) );
	vdp_nand3 g3535 (.Z(w3369), .A(w3364), .B(w3367), .C(w3356) );
	vdp_not g3536 (.nZ(w3408), .A(w3359) );
	vdp_not g3537 (.nZ(w3406), .A(w3361) );
	vdp_not g3538 (.nZ(w3405), .A(w3362) );
	vdp_not g3539 (.nZ(w3403), .A(w3366) );
	vdp_not g3540 (.nZ(w3404), .A(w3365) );
	vdp_not g3541 (.nZ(w3402), .A(w3369) );
	vdp_not g3542 (.nZ(w3401), .A(w3368) );
	vdp_not g3543 (.nZ(w3277), .A(w3287) );
	vdp_not g3544 (.nZ(w3285), .A(w3137) );
	vdp_not g3545 (.nZ(w3276), .A(w3284) );
	vdp_nand3 g3546 (.Z(w3289), .A(w3276), .B(w3137), .C(w3287) );
	vdp_not g3547 (.nZ(w3251), .A(w3291) );
	vdp_nand3 g3548 (.Z(w3291), .A(w3284), .B(w3285), .C(w3287) );
	vdp_nand3 g3549 (.Z(w3290), .A(w3284), .B(w3137), .C(w3287) );
	vdp_nand3 g3550 (.Z(w4058), .A(w3284), .B(w3137), .C(w3277) );
	vdp_nand3 g3551 (.Z(w3288), .A(w3276), .B(w3285), .C(w3287) );
	vdp_nand3 g3552 (.Z(w3286), .A(w3284), .B(w3285), .C(w3277) );
	vdp_not g3553 (.nZ(w3250), .A(w3290) );
	vdp_not g3554 (.nZ(w3256), .A(w3289) );
	vdp_not g3555 (.nZ(w3255), .A(w3288) );
	vdp_not g3556 (.nZ(w3254), .A(w3286) );
	vdp_not g3557 (.nZ(w3253), .A(w4058) );
	vdp_aon22 g3558 (.Z(w3292), .A1(w3295), .B1(w3302), .A2(w3303), .B2(w3053) );
	vdp_aon22 g3559 (.Z(w3293), .A1(w3297), .B1(w3302), .A2(w3303), .B2(w3296) );
	vdp_aon22 g3560 (.Z(w3242), .A1(w3299), .B1(w3302), .A2(w3303), .B2(w3298) );
	vdp_aon22 g3561 (.Z(w3139), .A1(w3301), .B1(w3302), .A2(w3303), .B2(w3300) );
	vdp_sr_bit g3562 (.Q(w3135), .D(w4053), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3563 (.Q(w4053), .D(w3134), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_xor g3564 (.Z(1'b1), .A(w3137), .B(w3131) );
	vdp_xor g3565 (.A(HPOS[3]), .B(w3154), .Z(w4107) );
	vdp_aon22 g3566 (.Z(w3192), .A1(w3185), .B1(w3186), .A2(w3184), .B2(w4106) );
	vdp_aon22 g3567 (.Z(w3193), .A1(w3187), .B1(w3186), .A2(w3184), .B2(w4105) );
	vdp_aon22 g3568 (.Z(w3195), .A1(w3188), .B1(w3186), .A2(w3184), .B2(w4104) );
	vdp_aon22 g3569 (.Z(w3194), .A1(w3189), .B1(w3186), .A2(w3184), .B2(w4103) );
	vdp_aon22 g3570 (.Z(w3632), .A1(w3190), .B1(w3186), .A2(w3184), .B2(w4102) );
	vdp_aon22 g3571 (.Z(w3237), .A1(w3332), .B1(w4045), .A2(w3230), .B2(w3331) );
	vdp_aon22 g3572 (.Z(w3241), .A1(w3332), .B1(w3231), .A2(w3232), .B2(w3331) );
	vdp_aon22 g3573 (.Z(w3239), .A1(w3332), .B1(w3236), .A2(w3235), .B2(w3331) );
	vdp_aon22 g3574 (.Z(w3240), .A1(w3332), .B1(w3233), .A2(w3234), .B2(w3331) );
	vdp_aon222 g3575 (.Z(w3457), .A1(w3449), .B1(w3448), .C1(w3447), .A2(w3394), .B2(w3395), .C2(w3393) );
	vdp_aon222 g3576 (.Z(w3460), .A1(w3453), .B1(w3418), .C1(w3452), .A2(w3394), .B2(w3395), .C2(w3393) );
	vdp_aon222 g3577 (.Z(w3434), .A1(w3454), .B1(w3451), .C1(w3419), .A2(w3394), .B2(w3395), .C2(w3393) );
	vdp_aon222 g3578 (.A1(w3455), .B1(w3420), .C1(w3450), .A2(w3394), .B2(w3395), .C2(w3393), .Z(w3456) );
	vdp_and5 g3579 (.Z(w3496), .A(w3446), .B(w3492), .C(w3485), .D(w3887), .E(w3479) );
	vdp_aon22 g3580 (.Z(w3443), .A1(w3351), .B1(w3552), .A2(w3171), .B2(w3350) );
	vdp_aon22 g3581 (.Z(w3442), .A1(w3353), .B1(w3552), .A2(w3171), .B2(w3352) );
	vdp_aon22 g3582 (.Z(w3441), .A1(w3355), .B1(w3552), .A2(w3171), .B2(w3354) );
	vdp_aon22 g3583 (.Z(w3444), .A1(w3349), .B1(w3552), .A2(w3171), .B2(w4452) );
	vdp_aon22 g3584 (.Z(w3151), .A1(w3438), .B1(w3175), .A2(w3152), .B2(M5) );
	vdp_and4 g3585 (.Z(w3439), .A(w3499), .B(w3445), .C(w3487), .D(w3440) );
	vdp_comp_we g3586 (.Z(w3171), .nZ(w3552), .A(w3437) );
	vdp_comp_we g3587 (.Z(w3331), .nZ(w3332), .A(w3130) );
	vdp_comp_we g3588 (.Z(w3303), .nZ(w3302), .A(w3130) );
	vdp_comp_we g3589 (.Z(w3142), .nZ(w3145), .A(w3224) );
	vdp_comp_we g3590 (.Z(w3184), .nZ(w3186), .A(w3722) );
	vdp_comp_we g3591 (.Z(w3172), .nZ(w3481), .A(w3446) );
	vdp_not g3592 (.nZ(w4073), .A(M5) );
	vdp_dlatch_inv g3593 (.nQ(w4062), .D(w3147), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g3594 (.Z(w3312), .A(DCLK2), .B(w3055) );
	vdp_and g3595 (.Z(w3313), .A(DCLK2), .B(w3054) );
	vdp_and g3596 (.Z(w3311), .A(DCLK2), .B(w3057) );
	vdp_and g3597 (.Z(w3310), .A(DCLK2), .B(w3058) );
	vdp_and g3598 (.Z(w3119), .A(w4062), .B(DCLK2) );
	vdp_and g3599 (.Z(w3120), .A(w4061), .B(DCLK2) );
	vdp_and g3600 (.Z(w3118), .A(w3548), .B(DCLK2) );
	vdp_and g3601 (.Z(w4059), .A(w4060), .B(DCLK2) );
	vdp_and g3602 (.Z(w3104), .A(DCLK2), .B(w4063) );
	vdp_and g3603 (.Z(w3416), .A(DCLK2), .B(w4031) );
	vdp_and g3604 (.Z(w3415), .A(DCLK2), .B(w4064) );
	vdp_and g3605 (.Z(w3096), .A(DCLK2), .B(w4065) );
	vdp_and g3606 (.Z(w3129), .A(w4050), .B(HCLK2) );
	vdp_and g3607 (.Z(w3305), .A(w3267), .B(w3138) );
	vdp_and g3608 (.Z(w3347), .A(w3497), .B(HCLK2) );
	vdp_or g3609 (.Z(w3440), .A(w4073), .B(w3397) );
	vdp_and g3610 (.Z(w3103), .A(w3151), .B(DCLK2) );
	vdp_and g3611 (.Z(w3495), .A(DCLK2), .B(w4067) );
	vdp_and g3612 (.Z(w3494), .A(DCLK2), .B(w4068) );
	vdp_and g3613 (.Z(w3493), .A(DCLK2), .B(w4069) );
	vdp_and g3614 (.Z(w3304), .A(DCLK2), .B(w4066) );
	vdp_and g3615 (.Z(w3437), .A(M5), .B(w3397) );
	vdp_and g3616 (.Z(w4103), .A(w44), .B(HPOS[7]) );
	vdp_and g3617 (.Z(w4102), .A(w44), .B(HPOS[8]) );
	vdp_and g3618 (.Z(w3183), .A(DCLK2), .B(w3176) );
	vdp_and g3619 (.Z(w4104), .A(w44), .B(HPOS[6]) );
	vdp_and g3620 (.Z(w3182), .A(DCLK2), .B(w4054) );
	vdp_and g3621 (.Z(w3181), .A(DCLK2), .B(w3540) );
	vdp_and g3622 (.Z(w3179), .A(DCLK2), .B(w3541) );
	vdp_and g3623 (.Z(w4105), .A(w44), .B(HPOS[5]) );
	vdp_and g3624 (.Z(w3051), .A(DCLK2), .B(w3175) );
	vdp_and g3625 (.Z(w4106), .A(w44), .B(HPOS[4]) );
	vdp_aon22 g3626 (.Z(w3191), .A1(w3153), .B1(w3186), .A2(w3184), .B2(w4107) );
	vdp_and g3627 (.nZ(w3154), .A(w44), .B(M5) );
	vdp_or4 g3628 (.Z(w2873), .D(w3219), .C(w3220), .B(w3221), .A(w3222) );
	vdp_or g3629 (.Z(w3224), .A(w92), .B(w3225) );
	vdp_or g3630 (.Z(w3446), .A(w10), .B(w90) );
	vdp_or4 g3631 (.Z(w2874), .A(w3554), .B(w3553), .C(w3538), .D(w3459) );
	vdp_not g3632 (.nZ(w4071), .A(w3400) );
	vdp_not g3633 (.nZ(w3134), .A(w3243) );
	vdp_not g3634 (.nZ(w3438), .A(M5) );
	vdp_aoi21 g3635 (.Z(w3400), .A1(w105), .A2(w3132), .B(w17) );
	vdp_aoi21 g3636 (.Z(w3243), .A1(w106), .A2(w3132), .B(w11) );
	vdp_aoi21 g3637 (.Z(w3265), .A1(w103), .A2(w3132), .B(w12) );
	vdp_nand4 g3638 (.D(w3130), .C(w3140), .Z(w4049), .A(w4043), .B(w3144) );
	vdp_nand3 g3639 (.Z(w3278), .A(w3276), .B(w3137), .C(w3277) );
	vdp_not g3640 (.nZ(w3258), .A(w3278) );
	vdp_nand3 g3641 (.Z(w3345), .A(w3277), .B(w3276), .C(w3285) );
	vdp_not g3642 (.nZ(w3248), .A(w3345) );
	vdp_not g3643 (.nZ(w3395), .A(w3391) );
	vdp_not g3644 (.nZ(w3394), .A(w3392) );
	vdp_not g3645 (.nZ(w4048), .A(w3397) );
	vdp_not g3646 (.nZ(w3393), .A(M5) );
	vdp_not g3647 (.nZ(w4077), .A(PLANE_A_PRIO) );
	vdp_not g3648 (.nZ(w4055), .A(PLANE_B_PRIO) );
	vdp_bufif0 g3649 (.Z(COL[5]), .A(w3226), .nE(w4055) );
	vdp_bufif0 g3650 (.Z(COL[6]), .A(w3307), .nE(w4055) );
	vdp_bufif0 g3651 (.Z(COL[4]), .A(w3228), .nE(w4055) );
	vdp_bufif0 g3652 (.Z(COL[3]), .A(w3229), .nE(w4055) );
	vdp_bufif0 g3653 (.Z(COL[2]), .A(w3223), .nE(w4055) );
	vdp_bufif0 g3654 (.Z(COL[1]), .A(w3238), .nE(w4055) );
	vdp_bufif0 g3655 (.Z(COL[0]), .A(w3227), .nE(w4055) );
	vdp_bufif0 g3656 (.Z(COL[5]), .A(w3432), .nE(w4077) );
	vdp_bufif0 g3657 (.Z(COL[6]), .A(w3539), .nE(w4077) );
	vdp_bufif0 g3658 (.Z(COL[4]), .A(w3431), .nE(w4077) );
	vdp_bufif0 g3659 (.Z(COL[3]), .A(w3433), .nE(w4077) );
	vdp_bufif0 g3660 (.Z(COL[2]), .A(w3398), .nE(w4077) );
	vdp_bufif0 g3661 (.Z(COL[1]), .A(w4076), .nE(w4077) );
	vdp_bufif0 g3662 (.Z(COL[0]), .A(w3458), .nE(w4077) );
	vdp_nand g3663 (.Z(w3141), .B(HCLK1), .A(w3135) );
	vdp_nand g3664 (.Z(w3147), .B(HCLK1), .A(w3134) );
	vdp_nand g3665 (.Z(w3100), .A(w3649), .B(HCLK1) );
	vdp_nand g3666 (.Z(w3050), .A(w4071), .B(HCLK1) );
	vdp_nor g3667 (.Z(w4072), .A(w3439), .B(w3496) );
	vdp_nand g3668 (.Z(w3150), .A(w4151), .B(HCLK1) );
	vdp_nand g3669 (.Z(w3392), .A(M5), .B(w3397) );
	vdp_nand g3670 (.Z(w3391), .A(M5), .B(w4048) );
	vdp_xor g3671 (.Z(w3569), .A(w3568), .B(w3567) );
	vdp_aon22 g3672 (.Z(w3567), .A1(w3565), .B1(w3644), .A2(VPOS[3]), .B2(w3566) );
	vdp_xnor g3673 (.Z(w3571), .A(w3568), .B(w3645) );
	vdp_aon22 g3674 (.Z(w3645), .A1(w3565), .B1(w3644), .A2(VPOS[2]), .B2(w3570) );
	vdp_xnor g3675 (.Z(w3573), .A(w3568), .B(w3643) );
	vdp_aon22 g3676 (.Z(w3643), .A1(w3565), .B1(w3644), .A2(VPOS[1]), .B2(w3572) );
	vdp_notif0 g3677 (.nZ(VRAMA[4]), .A(w3571), .nE(w3622) );
	vdp_notif0 g3678 (.nZ(VRAMA[3]), .A(w3573), .nE(w3622) );
	vdp_xnor g3679 (.Z(w3641), .A(w3568), .B(w3642) );
	vdp_aon22 g3680 (.Z(w3642), .A1(w3565), .B1(w3644), .A2(VPOS[0]), .B2(w3574) );
	vdp_notif0 g3681 (.nZ(VRAMA[2]), .A(w3641), .nE(w3622) );
	vdp_notif0 g3682 (.nZ(VRAMA[1]), .A(w3640), .nE(w3622) );
	vdp_notif0 g3683 (.nZ(VRAMA[0]), .A(1'b1), .nE(w3622) );
	vdp_not g3684 (.nZ(w3637), .A(w3648) );
	vdp_not g3685 (.nZ(w3622), .A(w3647) );
	vdp_comp_we g3686 (.Z(w3565), .nZ(w3644), .A(w4145) );
	vdp_comp_we g3687 (.Z(w3575), .nZ(w3639), .A(w1) );
	vdp_notif0 g3688 (.nZ(VRAMA[5]), .A(w3577), .nE(w3637) );
	vdp_aoi22 g3689 (.Z(w3577), .A1(w3569), .B1(w3576), .A2(w3575), .B2(w3639) );
	vdp_notif0 g3690 (.nZ(VRAMA[6]), .A(w3578), .nE(w3637) );
	vdp_aoi22 g3691 (.Z(w3578), .A1(w3576), .B1(w3579), .A2(w3575), .B2(w3639) );
	vdp_notif0 g3692 (.nZ(VRAMA[7]), .A(w3580), .nE(w3637) );
	vdp_aoi22 g3693 (.Z(w3580), .A1(w3579), .B1(w3581), .A2(w3575), .B2(w3639) );
	vdp_notif0 g3694 (.nZ(VRAMA[8]), .A(w3582), .nE(w3637) );
	vdp_aoi22 g3695 (.Z(w3582), .A1(w3581), .B1(w3583), .A2(w3575), .B2(w3639) );
	vdp_notif0 g3696 (.nZ(VRAMA[9]), .A(w4080), .nE(w3637) );
	vdp_aoi22 g3697 (.Z(w4080), .A1(w3583), .B1(w3585), .A2(w3575), .B2(w3639) );
	vdp_notif0 g3698 (.nZ(VRAMA[10]), .A(w3584), .nE(w3637) );
	vdp_aoi22 g3699 (.Z(w3584), .A1(w3585), .B1(w3586), .A2(w3575), .B2(w3639) );
	vdp_notif0 g3700 (.nZ(VRAMA[11]), .A(w4079), .nE(w3637) );
	vdp_aoi22 g3701 (.Z(w4079), .A1(w3586), .B1(w3588), .A2(w3575), .B2(w3639) );
	vdp_notif0 g3702 (.nZ(VRAMA[12]), .A(w3589), .nE(w3637) );
	vdp_aoi22 g3703 (.Z(w3589), .A1(w3588), .B1(w3587), .A2(w3575), .B2(w3639) );
	vdp_notif0 g3704 (.nZ(VRAMA[13]), .A(w3591), .nE(w3637) );
	vdp_aoi22 g3705 (.Z(w3591), .A1(w3587), .B1(w3590), .A2(w3575), .B2(w3639) );
	vdp_not g3706 (.nZ(w3638), .A(w4100) );
	vdp_notif0 g3707 (.nZ(VRAMA[14]), .A(w3593), .nE(w3638) );
	vdp_aoi22 g3708 (.Z(w3593), .A1(w3590), .B1(w3592), .A2(w3575), .B2(w3639) );
	vdp_notif0 g3709 (.nZ(VRAMA[15]), .A(w3595), .nE(w3638) );
	vdp_aoi22 g3710 (.Z(w3595), .A1(w3592), .B1(w3594), .A2(w3575), .B2(w3639) );
	vdp_notif0 g3711 (.nZ(VRAMA[16]), .A(w3597), .nE(w3638) );
	vdp_aoi22 g3712 (.Z(w3597), .A1(w3594), .B1(w3596), .A2(w3575), .B2(w3639) );
	vdp_notif0 g3713 (.nZ(VRAMA[5]), .A(w3600), .nE(w3636) );
	vdp_aoi22 g3714 (.Z(w3600), .A1(w3598), .B1(w3569), .A2(w3599), .B2(w3635) );
	vdp_notif0 g3715 (.nZ(VRAMA[6]), .A(w3602), .nE(w3636) );
	vdp_aoi22 g3716 (.Z(w3602), .A1(w3598), .B1(w3599), .A2(w3601), .B2(w3635) );
	vdp_notif0 g3717 (.nZ(VRAMA[7]), .A(w3603), .nE(w3636) );
	vdp_aoi22 g3718 (.Z(w3603), .A1(w3598), .B1(w3601), .A2(w3621), .B2(w3635) );
	vdp_notif0 g3719 (.nZ(VRAMA[8]), .A(w3604), .nE(w3636) );
	vdp_aoi22 g3720 (.Z(w3604), .A1(w3598), .B1(w3621), .A2(w3605), .B2(w3635) );
	vdp_notif0 g3721 (.nZ(VRAMA[9]), .A(w3606), .nE(w3636) );
	vdp_aoi22 g3722 (.Z(w3606), .A1(w3598), .B1(w3605), .A2(w3607), .B2(w3635) );
	vdp_notif0 g3723 (.nZ(VRAMA[10]), .A(w3609), .nE(w3636) );
	vdp_aoi22 g3724 (.Z(w3609), .A1(w3598), .B1(w3607), .A2(w3608), .B2(w3635) );
	vdp_notif0 g3725 (.nZ(VRAMA[11]), .A(w3611), .nE(w3634) );
	vdp_aoi22 g3726 (.Z(w3611), .A1(w3598), .B1(w3608), .A2(w3610), .B2(w3635) );
	vdp_notif0 g3727 (.nZ(VRAMA[12]), .A(w3613), .nE(w3634) );
	vdp_aoi22 g3728 (.Z(w3613), .A1(w3598), .B1(w3610), .A2(w3612), .B2(w3635) );
	vdp_notif0 g3729 (.nZ(VRAMA[14]), .A(w3616), .nE(w3634) );
	vdp_aoi22 g3730 (.Z(w3616), .A1(w3598), .B1(w3614), .A2(w3617), .B2(w3635) );
	vdp_notif0 g3731 (.nZ(VRAMA[15]), .A(w3619), .nE(w3634) );
	vdp_aoi22 g3732 (.Z(w3619), .A1(w3598), .B1(w3617), .A2(w3618), .B2(w3635) );
	vdp_notif0 g3733 (.nZ(VRAMA[16]), .A(w3620), .nE(w3634) );
	vdp_aoi22 g3734 (.Z(w3620), .A1(w3598), .B1(w3618), .A2(w3596), .B2(w3635) );
	vdp_notif0 g3735 (.nZ(VRAMA[13]), .A(w3615), .nE(w3634) );
	vdp_aoi22 g3736 (.Z(w3615), .A1(w3598), .B1(w3612), .A2(w3614), .B2(w3635) );
	vdp_not g3737 (.nZ(w3636), .A(w3564) );
	vdp_comp_we g3738 (.Z(w3635), .nZ(w3598), .A(w1) );
	vdp_aon22 g3739 (.Z(w3596), .A1(w3559), .B1(w3558), .A2(w3560), .B2(w3631) );
	vdp_not g3740 (.nZ(w3634), .A(w3564) );
	vdp_not g3741 (.nZ(w3560), .A(w3631) );
	vdp_sr_bit g3742 (.Q(w3647), .D(w3662), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3743 (.Q(w3631), .D(HPOS[3]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3744 (.Q(w3640), .D(w3701), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3745 (.Q(w3648), .D(w4153), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3746 (.Q(w3646), .D(w4144), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3747 (.Q(w3666), .D(w4143), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3748 (.Q(w3633), .D(w4142), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3749 (.Q(w4118), .D(w4119), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3750 (.Q(w4120), .D(w4118), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3751 (.Q(w3649), .D(w4120), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3752 (.Q(w3681), .D(w109), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3753 (.Q(w3659), .D(w37), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3754 (.Q(w4121), .D(w38), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3755 (.Q(w3723), .D(w4121), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3756 (.Q(w3724), .D(w3659), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3757 (.Q(w3721), .D(w3681), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3758 (.Q(w3725), .D(w3632), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3759 (.Q(w3726), .D(w3194), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3760 (.Q(w3727), .D(w3195), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3761 (.Q(w3728), .D(w3193), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3762 (.Q(w3756), .D(w3192), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3763 (.Q(w3757), .D(w3191), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3764 (.Q(w3657), .D(w3655), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3765 (.Q(w3658), .D(w3657), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3766 (.Q(w4122), .D(w3658), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_aon22 g3767 (.Z(w3671), .A1(H40), .B1(HPOS[8]), .A2(w3669), .B2(w3668) );
	vdp_aon22 g3768 (.Z(w3753), .A1(w3651), .B1(HPOS[8]), .A2(w3671), .B2(w3661) );
	vdp_aon22 g3769 (.Z(w3716), .A1(w3656), .B1(w3669), .A2(w3671), .B2(w3661) );
	vdp_or3 g3770 (.Z(w3722), .A(w3681), .B(w3659), .C(w4121) );
	vdp_or g3771 (.Z(w3672), .A(M5), .B(w3486) );
	vdp_bufif0 g3772 (.Z(VRAMA[1]), .A(w4117), .nE(w3660) );
	vdp_or g3773 (.Z(w3749), .A(w3671), .B(HPOS[4]) );
	vdp_bufif0 g3774 (.Z(VRAMA[2]), .A(w3674), .nE(w3660) );
	vdp_or g3775 (.Z(w3750), .A(w3671), .B(HPOS[5]) );
	vdp_bufif0 g3776 (.Z(VRAMA[3]), .A(w3675), .nE(w3660) );
	vdp_or g3777 (.Z(w3754), .A(w3671), .B(HPOS[6]) );
	vdp_bufif0 g3778 (.Z(VRAMA[4]), .A(w3676), .nE(w3660) );
	vdp_or g3779 (.Z(w3752), .A(w3671), .B(HPOS[7]) );
	vdp_bufif0 g3780 (.Z(VRAMA[5]), .A(w3677), .nE(w3660) );
	vdp_bufif0 g3781 (.Z(VRAMA[5]), .A(w3650), .nE(w3660) );
	vdp_not g3782 (.nZ(w3665), .A(w3557) );
	vdp_not g3783 (.nZ(w4123), .A(HPOS[3]) );
	vdp_dlatch_inv g3784 (.nQ(w3655), .D(w3654), .C(DCLK1), .nC(nDCLK1) );
	vdp_not g3785 (.nZ(w3669), .A(w4099) );
	vdp_not g3786 (.nZ(w3661), .A(w3671) );
	vdp_not g3787 (.nZ(w3668), .A(H40) );
	vdp_not g3788 (.nZ(w3660), .A(w3667) );
	vdp_bufif0 g3789 (.Z(VRAMA[0]), .A(1'b0), .nE(w3660) );
	vdp_or g3790 (.Z(w3667), .A(w3646), .B(w3666) );
	vdp_or g3791 (.Z(w4119), .A(w3664), .B(w6) );
	vdp_nand3 g3792 (.Z(w3720), .A(M5), .B(w3665), .C(HPOS[3]) );
	vdp_nand3 g3793 (.Z(w3679), .A(M5), .B(w3665), .C(w4123) );
	vdp_and g3794 (.Z(w3680), .A(DCLK2), .B(w4122) );
	vdp_and g3795 (.Z(w3653), .A(w3658), .B(DCLK2) );
	vdp_and g3796 (.Z(w3719), .A(w3657), .B(DCLK2) );
	vdp_and g3797 (.Z(w3652), .A(w3655), .B(DCLK2) );
	vdp_and g3798 (.Z(w4100), .A(M5), .B(w3648) );
	vdp_and g3799 (.Z(w3709), .A(HPOS[3]), .B(w3670) );
	vdp_and g3800 (.Z(w4142), .A(w3557), .B(w6) );
	vdp_and g3801 (.Z(w4143), .A(w3665), .B(w6) );
	vdp_and3 g3802 (.Z(w4144), .A(w3664), .B(M5), .C(w3663) );
	vdp_nor g3803 (.Z(w3670), .A(M5), .B(w3671) );
	vdp_nand g3804 (.Z(w3654), .A(w3306), .B(HCLK1) );
	vdp_oai21 g3805 (.A1(HPOS[6]), .A2(HPOS[7]), .B(HPOS[8]), .Z(w4099) );
	vdp_slatch g3806 (.Q(w3696), .D(w612), .C(w3744), .nC(w3743) );
	vdp_slatch g3807 (.Q(w3692), .D(S[0]), .C(w3739), .nC(w3738) );
	vdp_slatch g3808 (.Q(w3693), .D(S[0]), .C(w3740), .nC(w3737) );
	vdp_slatch g3809 (.Q(w3694), .D(w685), .C(w3744), .nC(w3743) );
	vdp_slatch g3810 (.Q(w3690), .D(S[1]), .C(w3739), .nC(w3738) );
	vdp_slatch g3811 (.Q(w3765), .D(S[1]), .C(w3740), .nC(w3737) );
	vdp_slatch g3812 (.Q(w3766), .D(w698), .C(w3744), .nC(w3743) );
	vdp_slatch g3813 (.Q(w3684), .D(S[2]), .C(w3739), .nC(w3738) );
	vdp_slatch g3814 (.Q(w3767), .D(S[2]), .C(w3740), .nC(w3737) );
	vdp_slatch g3815 (.Q(w3763), .D(w719), .C(w3744), .nC(w3743) );
	vdp_slatch g3816 (.Q(w3762), .D(S[3]), .C(w3739), .nC(w3738) );
	vdp_slatch g3817 (.Q(w4441), .D(S[3]), .C(w3740), .nC(w3737) );
	vdp_slatch g3818 (.Q(w3708), .D(w725), .C(w3744), .nC(w3743) );
	vdp_slatch g3819 (.Q(w3761), .D(S[4]), .C(w3739), .nC(w3738) );
	vdp_slatch g3820 (.Q(w3760), .D(S[4]), .C(w3740), .nC(w3737) );
	vdp_slatch g3821 (.Q(w3759), .D(w681), .C(w3744), .nC(w3743) );
	vdp_slatch g3822 (.Q(w3747), .D(S[5]), .C(w3739), .nC(w3738) );
	vdp_slatch g3823 (.Q(w3746), .D(S[5]), .C(w3740), .nC(w3737) );
	vdp_slatch g3824 (.Q(w3745), .D(w661), .C(w3744), .nC(w3743) );
	vdp_slatch g3825 (.Q(w3741), .D(S[6]), .C(w3739), .nC(w3738) );
	vdp_slatch g3826 (.Q(w3742), .D(S[6]), .C(w3740), .nC(w3737) );
	vdp_slatch g3827 (.Q(w3736), .D(w617), .C(w3744), .nC(w3743) );
	vdp_slatch g3828 (.Q(w3735), .D(S[7]), .C(w3739), .nC(w3738) );
	vdp_slatch g3829 (.Q(w3734), .D(S[7]), .C(w3740), .nC(w3737) );
	vdp_slatch g3830 (.Q(w3732), .D(S[0]), .C(w3712), .nC(w3729) );
	vdp_slatch g3831 (.Q(w3714), .D(S[0]), .C(w3713), .nC(w3733) );
	vdp_slatch g3832 (.Q(w3718), .D(S[1]), .C(w3713), .nC(w3733) );
	vdp_slatch g3833 (.Q(w3717), .D(S[1]), .C(w3712), .nC(w3729) );
	vdp_slatch g3834 (.Q(w3710), .D(w3736), .C(w3689), .nC(w3688) );
	vdp_slatch g3835 (.Q(w3704), .D(w3745), .C(w3689), .nC(w3688) );
	vdp_slatch g3836 (.Q(w3707), .D(w3759), .C(w3689), .nC(w3688) );
	vdp_slatch g3837 (.Q(w3769), .D(w3708), .C(w3689), .nC(w3688) );
	vdp_slatch g3838 (.Q(w3682), .D(w3763), .C(w3689), .nC(w3688) );
	vdp_slatch g3839 (.Q(w3683), .D(w3766), .C(w3689), .nC(w3688) );
	vdp_slatch g3840 (.Q(w3691), .D(w3694), .C(w3689), .nC(w3688) );
	vdp_slatch g3841 (.Q(w3695), .D(w3696), .C(w3689), .nC(w3688) );
	vdp_fa g3842 (.CI(w4097), .SUM(w4042), .B(w3716), .A(w3731) );
	vdp_fa g3843 (.CO(w4097), .CI(w3715), .SUM(w3914), .B(w3753), .A(w3758) );
	vdp_fa g3844 (.CO(w3758), .CI(w3711), .SUM(w3677), .B(w3752), .A(w4096) );
	vdp_fa g3845 (.CO(w4096), .CI(w3705), .SUM(w3676), .B(w3754), .A(w3755) );
	vdp_fa g3846 (.CO(w3755), .CI(w3706), .SUM(w3675), .B(w3750), .A(w3751) );
	vdp_fa g3847 (.CO(w3751), .CI(w3810), .SUM(w3674), .B(w3749), .A(w3748) );
	vdp_fa g3848 (.CO(w3748), .CI(w3672), .SUM(w4117), .B(w3709), .A(1'b1) );
	vdp_aon222 g3849 (.A1(w3686), .B1(w3673), .C1(w3685), .A2(w3717), .B2(w3718), .C2(1'b0), .Z(w3731) );
	vdp_aon222 g3850 (.A1(w3686), .B1(w3673), .C1(w3685), .A2(w3732), .B2(w3714), .C2(1'b0), .Z(w3715) );
	vdp_aon222 g3851 (.A1(w3686), .B1(w3673), .C1(w3685), .A2(w3734), .B2(w3735), .C2(w3710), .Z(w3711) );
	vdp_aon222 g3852 (.A1(w3686), .B1(w3673), .C1(w3685), .A2(w3742), .B2(w3741), .C2(w3704), .Z(w3705) );
	vdp_aon222 g3853 (.A1(w3686), .B1(w3673), .C1(w3685), .A2(w3746), .B2(w3747), .C2(w3707), .Z(w3706) );
	vdp_aon222 g3854 (.A1(w3686), .B1(w3673), .C1(w3685), .A2(w3760), .B2(w3761), .C2(w3769), .Z(w3810) );
	vdp_aon222 g3855 (.A1(w3686), .B1(w3673), .C1(w3685), .A2(w4441), .B2(w3762), .C2(w3682), .Z(w3486) );
	vdp_aon222 g3856 (.A1(w3686), .B1(w3673), .C1(w3685), .A2(w3767), .B2(w3684), .C2(w3683), .Z(w3180) );
	vdp_aon222 g3857 (.A1(w3686), .B1(w3673), .A2(w3765), .B2(w3690), .C2(w3691), .Z(w3484), .C1(w3685) );
	vdp_aon222 g3858 (.A1(w3686), .B1(w3673), .C1(w3685), .A2(w3693), .B2(w3692), .C2(w3695), .Z(w3482) );
	vdp_comp_strong g3859 (.Z(w3712), .nZ(w3729), .A(w3680) );
	vdp_comp_strong g3860 (.Z(w3713), .nZ(w3733), .A(w3719) );
	vdp_not g3861 (.nZ(w3673), .A(w3679) );
	vdp_not g3862 (.nZ(w3686), .A(w3720) );
	vdp_not g3863 (.nZ(w3685), .A(w3764) );
	vdp_not g3864 (.nZ(w3699), .A(w96) );
	vdp_not g3865 (.nZ(w3663), .A(w104) );
	vdp_not g3866 (.nZ(w3700), .A(w3701) );
	vdp_not g3867 (.nZ(w3664), .A(w3702) );
	vdp_not g3868 (.nZ(w3703), .A(M5) );
	vdp_comp_strong g3869 (.Z(w3739), .nZ(w3738), .A(w3652) );
	vdp_comp_strong g3870 (.Z(w3740), .nZ(w3737), .A(w3653) );
	vdp_comp_strong g3871 (.Z(w3744), .nZ(w3743), .A(w86) );
	vdp_comp_strong g3872 (.Z(w3689), .nZ(w3688), .A(w3768) );
	vdp_or g3873 (.Z(w3764), .A(w4101), .B(M5) );
	vdp_or g3874 (.Z(w4153), .A(w13), .B(w3700) );
	vdp_or g3875 (.Z(w3662), .A(w13), .B(w14) );
	vdp_or g3876 (.Z(w3768), .A(w4), .B(w103) );
	vdp_or5 g3877 (.E(w3699), .C(w3698), .D(VPOS[5]), .Z(w4101), .A(w3697), .B(VPOS[4]) );
	vdp_aoi21 g3878 (.Z(w3702), .A1(w104), .A2(w3132), .B(w8) );
	vdp_nand g3879 (.Z(w3701), .A(w14), .B(w3703) );
	vdp_slatch g3880 (.Q(w3805), .D(w4431), .C(w3774), .nC(w3775) );
	vdp_slatch g3881 (.Q(w3780), .D(w4432), .C(w3774), .nC(w3775) );
	vdp_slatch g3882 (.Q(w3781), .D(w4433), .C(w3774), .nC(w3775) );
	vdp_slatch g3883 (.Q(w3782), .D(w4430), .C(w3774), .nC(w3775) );
	vdp_slatch g3884 (.Q(w3785), .D(w4429), .C(w3774), .nC(w3775) );
	vdp_slatch g3885 (.Q(w3784), .D(w4428), .C(w3774), .nC(w3775) );
	vdp_slatch g3886 (.nQ(w3790), .D(w4436), .C(w3776), .nC(w3777) );
	vdp_slatch g3887 (.Q(w3783), .D(w4437), .C(w3776), .nC(w3777) );
	vdp_slatch g3888 (.Q(w3789), .D(w4438), .C(w3776), .nC(w3777) );
	vdp_slatch g3889 (.Q(w3788), .D(w4439), .C(w3776), .nC(w3777) );
	vdp_slatch g3890 (.Q(w3787), .D(w4435), .C(w3776), .nC(w3777) );
	vdp_slatch g3891 (.Q(w3786), .D(w4434), .C(w3776), .nC(w3777) );
	vdp_comp_strong g3892 (.Z(w3774), .nZ(w3775), .A(w3795) );
	vdp_comp_strong g3893 (.Z(w3776), .nZ(w3777), .A(w4124) );
	vdp_cgi2a g3894 (.Z(w4041), .A(w3786), .B(HPOS[4]), .C(1'b1) );
	vdp_cgi2a g3895 (.Z(w4036), .A(w3787), .B(HPOS[5]), .C(w4041) );
	vdp_cgi2a g3896 (.Z(w4035), .A(w3788), .B(HPOS[6]), .C(w4036) );
	vdp_cgi2a g3897 (.Z(w4037), .A(w3789), .B(HPOS[7]), .C(w4035) );
	vdp_cgi2a g3898 (.X(w3791), .A(w3783), .B(HPOS[8]), .C(w4037) );
	vdp_cgi2a g3899 (.Z(w3796), .A(w3793), .B(w3780), .C(w4126) );
	vdp_cgi2a g3900 (.Z(w4126), .A(w3794), .B(w3781), .C(w4038) );
	vdp_cgi2a g3901 (.Z(w4038), .A(w3797), .B(w3782), .C(w4039) );
	vdp_cgi2a g3902 (.Z(w4039), .A(w3800), .B(w3785), .C(w4040) );
	vdp_cgi2a g3903 (.Z(w4040), .A(w3799), .B(w3784), .C(1'b0) );
	vdp_slatch g3904 (.Q(w4431), .D(w617), .C(w3802), .nC(w3779) );
	vdp_slatch g3905 (.Q(w4432), .D(w725), .C(w3802), .nC(w3779) );
	vdp_slatch g3906 (.Q(w4433), .D(w719), .C(w3802), .nC(w3779) );
	vdp_slatch g3907 (.Q(w4430), .D(w698), .C(w3802), .nC(w3779) );
	vdp_slatch g3908 (.Q(w4429), .D(w685), .C(w3802), .nC(w3779) );
	vdp_slatch g3909 (.Q(w4428), .D(w612), .C(w3802), .nC(w3779) );
	vdp_comp_strong g3910 (.Z(w3802), .nZ(w3779), .A(w75) );
	vdp_slatch g3911 (.Q(w4436), .D(w617), .C(w3803), .nC(w3801) );
	vdp_slatch g3912 (.Q(w4437), .D(w725), .C(w3803), .nC(w3801) );
	vdp_slatch g3913 (.Q(w4438), .D(w719), .C(w3803), .nC(w3801) );
	vdp_slatch g3914 (.Q(w4439), .D(w698), .C(w3803), .nC(w3801) );
	vdp_slatch g3915 (.Q(w4435), .D(w685), .C(w3803), .nC(w3801) );
	vdp_slatch g3916 (.Q(w4434), .D(w612), .C(w3803), .nC(w3801) );
	vdp_comp_strong g3917 (.Z(w3803), .nZ(w3801), .A(w74) );
	vdp_xor g3918 (.Z(w3804), .A(w3805), .B(w3796) );
	vdp_xor g3919 (.Z(w3792), .A(w3790), .B(w3791) );
	vdp_aon22 g3920 (.Z(w3793), .A1(w3798), .B1(w3807), .A2(VPOS[8]), .B2(VPOS[7]) );
	vdp_aon22 g3921 (.Z(w3794), .A1(w3798), .B1(w3807), .A2(VPOS[7]), .B2(VPOS[6]) );
	vdp_aon22 g3922 (.Z(w3797), .A1(w3798), .B1(w3807), .A2(VPOS[6]), .B2(VPOS[5]) );
	vdp_aon22 g3923 (.Z(w3800), .A1(w3798), .B1(w3807), .A2(VPOS[5]), .B2(VPOS[4]) );
	vdp_aon22 g3924 (.Z(w3799), .A1(w3798), .B1(w3807), .A2(VPOS[4]), .B2(VPOS[3]) );
	vdp_aon22 g3925 (.Z(w3815), .A1(w3798), .B1(w3807), .A2(VPOS[3]), .B2(VPOS[2]) );
	vdp_aon22 g3926 (.Z(w3814), .A1(w3798), .B1(w3807), .A2(VPOS[2]), .B2(VPOS[1]) );
	vdp_aon22 g3927 (.Z(w3813), .A1(w3798), .B1(w3807), .A2(VPOS[1]), .B2(VPOS[0]) );
	vdp_comp_we g3928 (.Z(w3798), .nZ(w3807), .A(w1) );
	vdp_not g3929 (.nZ(w3557), .A(w4125) );
	vdp_not g3930 (.nZ(w3557), .A(HPOS[3]) );
	vdp_not g3931 (.nZ(w4128), .A(w4127) );
	vdp_or g3932 (.Z(w4124), .A(w103), .B(w4) );
	vdp_or g3933 (.Z(w3795), .A(w103), .B(w4128) );
	vdp_oai21 g3934 (.Z(w4127), .A1(w5), .A2(M5), .B(w4) );
	vdp_and g3935 (.Z(w3806), .A(w3792), .B(w3808) );
	vdp_oai211 g3936 (.Z(w4125), .A1(w3557), .A2(M5), .B(w3806), .C(w3804) );
	vdp_slatch g3937 (.nQ(w3848), .D(w725), .C(w3820), .nC(w3821) );
	vdp_slatch g3938 (.nQ(w3850), .D(w725), .C(w3818), .nC(w3819) );
	vdp_slatch g3939 (.nQ(w3849), .D(w681), .C(w3820), .nC(w3821) );
	vdp_slatch g3940 (.nQ(w3851), .D(w681), .C(w3818), .nC(w3819) );
	vdp_slatch g3941 (.nQ(w3824), .D(w661), .C(w3820), .nC(w3821) );
	vdp_slatch g3942 (.nQ(w3825), .D(w661), .C(w3818), .nC(w3819) );
	vdp_slatch g3943 (.nQ(w4427), .D(w685), .C(w3818), .nC(w3819) );
	vdp_slatch g3944 (.nQ(w3844), .D(w698), .C(w3820), .nC(w3821) );
	vdp_slatch g3945 (.nQ(w3845), .D(w698), .C(w3818), .nC(w3819) );
	vdp_slatch g3946 (.nQ(w3846), .D(w719), .C(w3820), .nC(w3821) );
	vdp_slatch g3947 (.nQ(w3847), .D(w719), .C(w3818), .nC(w3819) );
	vdp_slatch g3948 (.nQ(w3852), .D(w612), .C(w3818), .nC(w3819) );
	vdp_slatch g3949 (.nQ(w3822), .D(w685), .C(w3820), .nC(w3821) );
	vdp_slatch g3950 (.Q(w3559), .D(w612), .C(w3811), .nC(w3812) );
	vdp_slatch g3951 (.Q(w3558), .D(w725), .C(w3811), .nC(w3812) );
	vdp_not g3952 (.nZ(w4130), .A(w3822) );
	vdp_aoi22 g3953 (.Z(w3841), .A1(HPOS[8]), .B1(w3799), .A2(w3817), .B2(w3816) );
	vdp_aoi22 g3954 (.Z(w3842), .A1(w3799), .B1(w3800), .A2(w3817), .B2(w3816) );
	vdp_aoi22 g3955 (.Z(w3829), .A1(w3800), .B1(w3797), .A2(w3817), .B2(w3816) );
	vdp_aoi22 g3956 (.Z(w3854), .A1(w3794), .B1(w3793), .A2(w3817), .B2(w3816) );
	vdp_aoi22 g3957 (.Z(w3843), .A1(w3797), .B1(w3794), .A2(w3817), .B2(w3816) );
	vdp_comp_strong g3958 (.Z(w3811), .nZ(w3812), .A(w85) );
	vdp_comp_strong g3959 (.Z(w3820), .nZ(w3821), .A(w71) );
	vdp_comp_strong g3960 (.Z(w3818), .nZ(w3819), .A(w68) );
	vdp_aoi22 g3961 (.Z(w3853), .A1(w3793), .B1(w3816), .A2(w3817), .B2(w4130) );
	vdp_nand g3962 (.Z(w3855), .A(w3793), .B(w93) );
	vdp_nand g3963 (.Z(w3828), .A(w3794), .B(w93) );
	vdp_nand g3964 (.Z(w3856), .A(w3800), .B(w93) );
	vdp_nand g3965 (.Z(w3830), .A(w3797), .B(w93) );
	vdp_nand g3966 (.Z(w3840), .A(w3799), .B(w93) );
	vdp_nand g3967 (.Z(w4129), .A(w3815), .B(w91) );
	vdp_nand g3968 (.Z(w4154), .A(w3814), .B(w91) );
	vdp_nand g3969 (.Z(w3836), .A(w3813), .B(w91) );
	vdp_nand g3970 (.Z(w3808), .A(HPOS[7]), .B(HPOS[8]) );
	vdp_comp_we g3971 (.Z(w3817), .nZ(w3816), .A(H40) );
	vdp_notif0 g3972 (.nZ(VRAMA[16]), .A(w3825), .nE(w3823) );
	vdp_notif0 g3973 (.nZ(VRAMA[16]), .A(w3824), .nE(w3827) );
	vdp_notif0 g3974 (.nZ(VRAMA[15]), .A(w3851), .nE(w3823) );
	vdp_notif0 g3975 (.nZ(VRAMA[15]), .A(w3849), .nE(w3827) );
	vdp_notif0 g3976 (.nZ(VRAMA[14]), .A(w3850), .nE(w3823) );
	vdp_notif0 g3977 (.nZ(VRAMA[14]), .A(w3848), .nE(w3827) );
	vdp_notif0 g3978 (.nZ(VRAMA[13]), .A(w3847), .nE(w3823) );
	vdp_notif0 g3979 (.nZ(VRAMA[13]), .A(w3846), .nE(w3827) );
	vdp_notif0 g3980 (.nZ(VRAMA[12]), .A(w3845), .nE(w3823) );
	vdp_notif0 g3981 (.nZ(VRAMA[12]), .A(w3844), .nE(w3827) );
	vdp_notif0 g3982 (.nZ(VRAMA[11]), .A(w4427), .nE(w3823) );
	vdp_notif0 g3983 (.nZ(VRAMA[11]), .A(w3853), .nE(w3827) );
	vdp_notif0 g3984 (.nZ(VRAMA[10]), .A(w3852), .nE(w3823) );
	vdp_notif0 g3985 (.nZ(VRAMA[10]), .A(w3854), .nE(w3827) );
	vdp_notif0 g3986 (.nZ(VRAMA[9]), .A(w3855), .nE(w3826) );
	vdp_notif0 g3987 (.nZ(VRAMA[9]), .A(w3843), .nE(w3827) );
	vdp_notif0 g3988 (.nZ(VRAMA[6]), .A(w3856), .nE(w3826) );
	vdp_notif0 g3989 (.nZ(VRAMA[6]), .A(w3841), .nE(w3831) );
	vdp_notif0 g3990 (.nZ(VRAMA[5]), .A(w3840), .nE(w3826) );
	vdp_notif0 g3991 (.nZ(VRAMA[5]), .A(w3839), .nE(w3831) );
	vdp_notif0 g3992 (.nZ(VRAMA[4]), .A(w4129), .nE(w3826) );
	vdp_notif0 g3993 (.nZ(VRAMA[4]), .A(w3838), .nE(w3831) );
	vdp_notif0 g3994 (.nZ(VRAMA[3]), .A(w4154), .nE(w3826) );
	vdp_notif0 g3995 (.nZ(VRAMA[3]), .A(w3837), .nE(w3831) );
	vdp_notif0 g3996 (.nZ(VRAMA[2]), .A(w3836), .nE(w3826) );
	vdp_notif0 g3997 (.nZ(VRAMA[2]), .A(w3835), .nE(w3831) );
	vdp_notif0 g3998 (.A(1'b1), .nE(w3826) );
	vdp_notif0 g3999 (.A(1'b1), .nE(w3831) );
	vdp_notif0 g4000 (.A(w3833), .nE(w3826) );
	vdp_notif0 g4001 (.A(w3833), .nE(w3831) );
	vdp_notif0 g4002 (.nZ(VRAMA[8]), .A(w3828), .nE(w3826) );
	vdp_notif0 g4003 (.nZ(VRAMA[8]), .A(w3829), .nE(w3831) );
	vdp_notif0 g4004 (.nZ(VRAMA[7]), .A(w3830), .nE(w3826) );
	vdp_notif0 g4005 (.nZ(VRAMA[7]), .A(w3842), .nE(w3831) );
	vdp_not g4006 (.nZ(w3833), .A(1'b0) );
	vdp_not g4007 (.nZ(w3835), .A(HPOS[4]) );
	vdp_not g4008 (.nZ(w3837), .A(HPOS[5]) );
	vdp_not g4009 (.nZ(w3838), .A(HPOS[6]) );
	vdp_not g4010 (.nZ(w3839), .A(HPOS[7]) );
	vdp_not g4011 (.nZ(w3826), .A(w3305) );
	vdp_not g4012 (.nZ(w3823), .A(w3305) );
	vdp_not g4013 (.nZ(w3831), .A(w3633) );
	vdp_not g4014 (.nZ(w3827), .A(w3633) );
	vdp_not g4015 (.nZ(w3865), .A(w4034) );
	vdp_comp_strong g4016 (.Z(w3859), .nZ(w3860), .A(w70) );
	vdp_comp_we g4017 (.Z(w3864), .nZ(w3863), .A(w3646) );
	vdp_comp_strong g4018 (.Z(w3862), .nZ(w3861), .A(w72) );
	vdp_slatch g4019 (.Q(w3885), .D(w661), .C(w3859), .nC(w3860) );
	vdp_slatch g4020 (.Q(w4139), .D(w719), .C(w3862), .nC(w3861) );
	vdp_slatch g4021 (.Q(w3884), .D(w681), .C(w3859), .nC(w3860) );
	vdp_slatch g4022 (.Q(w3882), .D(w698), .C(w3862), .nC(w3861) );
	vdp_slatch g4023 (.Q(w3868), .D(w725), .C(w3859), .nC(w3860) );
	vdp_slatch g4024 (.Q(w4442), .D(w685), .C(w3862), .nC(w3861) );
	vdp_slatch g4025 (.Q(w3871), .D(w719), .C(w3859), .nC(w3860) );
	vdp_slatch g4026 (.Q(w4140), .D(w612), .C(w3862), .nC(w3861) );
	vdp_slatch g4027 (.Q(w3879), .D(w685), .C(w3859), .nC(w3860) );
	vdp_slatch g4028 (.Q(w3876), .D(w698), .C(w3859), .nC(w3860) );
	vdp_bufif0 g4029 (.Z(VRAMA[11]), .A(w3878), .nE(w3867) );
	vdp_bufif0 g4030 (.Z(VRAMA[10]), .A(w3872), .nE(w3867) );
	vdp_bufif0 g4031 (.Z(VRAMA[13]), .A(w3880), .nE(w3867) );
	vdp_bufif0 g4032 (.Z(VRAMA[9]), .A(w3870), .nE(w3867) );
	vdp_bufif0 g4033 (.Z(VRAMA[8]), .A(w3869), .nE(w3867) );
	vdp_bufif0 g4034 (.Z(VRAMA[14]), .A(w3881), .nE(w3865) );
	vdp_bufif0 g4035 (.Z(VRAMA[7]), .A(w3866), .nE(w3867) );
	vdp_bufif0 g4036 (.Z(VRAMA[15]), .A(w4098), .nE(w3865) );
	vdp_bufif0 g4037 (.Z(VRAMA[16]), .A(w3883), .nE(w3865) );
	vdp_aon22 g4038 (.Z(w3883), .A1(w3863), .B1(w3864), .A2(w3885), .B2(w4139) );
	vdp_aon22 g4039 (.Z(w4098), .A1(w3863), .B1(w3864), .A2(w3884), .B2(w3882) );
	vdp_aon22 g4040 (.Z(w3881), .A1(w3863), .B1(w3864), .A2(w3868), .B2(w4442) );
	vdp_aon22 g4041 (.Z(w3880), .A1(w3863), .B1(w3864), .A2(w3871), .B2(w4140) );
	vdp_aon22 g4042 (.Z(w3878), .A1(w3874), .B1(w3877), .A2(w3879), .B2(w3875) );
	vdp_aon22 g4043 (.Z(w3873), .A1(w3874), .B1(w3888), .A2(w3876), .B2(w3875) );
	vdp_bufif0 g4044 (.Z(VRAMA[12]), .A(w3873), .nE(w3867) );
	vdp_not g4045 (.nZ(w3867), .A(w3667) );
	vdp_and g4046 (.Z(w4034), .A(w3667), .B(M5) );
	vdp_comp_we g4047 (.Z(w3875), .nZ(w3874), .A(M5) );
	vdp_fa g4048 (.CO(w3903), .CI(w4087), .SUM(w3923), .B(VPOS[6]), .A(w4086) );
	vdp_fa g4049 (.CO(w4086), .CI(w4089), .SUM(w3904), .B(VPOS[5]), .A(w4088) );
	vdp_fa g4050 (.CO(w4088), .CI(w4091), .SUM(w3905), .B(VPOS[4]), .A(w4090) );
	vdp_fa g4051 (.CO(w4090), .CI(w3971), .SUM(w3566), .B(VPOS[3]), .A(w4092) );
	vdp_fa g4052 (.CO(w4092), .CI(w4094), .SUM(w3570), .B(VPOS[2]), .A(w4093) );
	vdp_fa g4053 (.CO(w4093), .CI(w4029), .SUM(w3572), .B(VPOS[1]), .A(w4095) );
	vdp_fa g4054 (.CO(w4095), .CI(w3984), .SUM(w3574), .B(VPOS[0]), .A(1'b0) );
	vdp_fa g4055 (.CO(w3922), .CI(w4085), .SUM(w3920), .B(VPOS[7]), .A(w3903) );
	vdp_fa g4056 (.CO(w3902), .CI(w3957), .SUM(w3931), .B(VPOS[8]), .A(w3922) );
	vdp_fa g4057 (.CO(w3930), .CI(w3958), .SUM(w3897), .B(1'b0), .A(w3902) );
	vdp_fa g4058 (.CI(w3942), .SUM(w3898), .B(1'b0), .A(w3930) );
	vdp_aon22 g4059 (.Z(w3942), .A1(w3940), .B1(w3941), .A2(w3901), .B2(w3900) );
	vdp_aon22 g4060 (.Z(w3958), .A1(w4032), .B1(w3945), .A2(w3901), .B2(w3900) );
	vdp_aon22 g4061 (.Z(w3957), .A1(w3946), .B1(w3947), .A2(w3901), .B2(w3900) );
	vdp_aon22 g4062 (.Z(w4085), .A1(w3949), .B1(w3950), .A2(w3901), .B2(w3900) );
	vdp_aon22 g4063 (.Z(w4087), .A1(w3956), .B1(w3953), .A2(w3901), .B2(w3900) );
	vdp_aon22 g4064 (.Z(w4089), .A1(w3961), .B1(w3960), .A2(w3901), .B2(w3900) );
	vdp_aon22 g4065 (.Z(w4091), .A1(w3965), .B1(w3966), .A2(w3901), .B2(w3900) );
	vdp_aon22 g4066 (.Z(w3971), .A1(w3970), .B1(w3969), .A2(w3901), .B2(w3900) );
	vdp_aon22 g4067 (.Z(w4094), .A1(w3972), .B1(w3973), .A2(w3901), .B2(w3900) );
	vdp_aon22 g4068 (.Z(w4029), .A1(w3976), .B1(w4033), .A2(w3901), .B2(w3900) );
	vdp_aon22 g4069 (.Z(w3984), .A1(w3978), .B1(w3977), .A2(w3901), .B2(w3900) );
	vdp_comp_we g4070 (.Z(w3901), .nZ(w3900), .A(w3909) );
	vdp_comp_strong g4071 (.Z(w3911), .nZ(w3906), .A(w69) );
	vdp_sr_bit g4072 (.Q(w3932), .D(RD_DATA[1]), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4073 (.Q(w3907), .D(RD_DATA[2]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4074 (.Q(w3981), .D(w3932), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4075 (.Q(w3999), .D(w3907), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4076 (.Q(w3980), .D(HPOS[3]), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4077 (.Q(w3651), .D(w612), .C(w3911), .nC(w3906) );
	vdp_slatch g4078 (.Q(w3656), .D(w685), .C(w3911), .nC(w3906) );
	vdp_slatch g4079 (.Q(w3927), .D(w681), .C(w3911), .nC(w3906) );
	vdp_slatch g4080 (.Q(w3926), .D(w725), .C(w3911), .nC(w3906) );
	vdp_slatch g4081 (.Q(w3978), .D(w3982), .C(w3933), .nC(w3937) );
	vdp_slatch g4082 (.Q(w4150), .D(w3983), .C(w3939), .nC(w3934) );
	vdp_slatch g4083 (.Q(w3976), .D(w3975), .C(w3933), .nC(w3937) );
	vdp_slatch g4084 (.Q(w4149), .D(w3974), .C(w3939), .nC(w3934) );
	vdp_slatch g4085 (.Q(w3972), .D(w4001), .C(w3933), .nC(w3937) );
	vdp_slatch g4086 (.Q(w4148), .D(w3968), .C(w3939), .nC(w3934) );
	vdp_slatch g4087 (.Q(w3970), .D(w3967), .C(w3933), .nC(w3937) );
	vdp_slatch g4088 (.Q(w4147), .D(w3964), .C(w3939), .nC(w3934) );
	vdp_slatch g4089 (.Q(w3965), .D(w3963), .C(w3933), .nC(w3937) );
	vdp_slatch g4090 (.Q(w4146), .D(w3962), .C(w3939), .nC(w3934) );
	vdp_slatch g4091 (.Q(w3961), .D(w3955), .C(w3933), .nC(w3937) );
	vdp_slatch g4092 (.Q(w4157), .D(w3954), .C(w3939), .nC(w3934) );
	vdp_slatch g4093 (.Q(w3956), .D(w3951), .C(w3933), .nC(w3937) );
	vdp_slatch g4094 (.Q(w4158), .D(w3952), .C(w3939), .nC(w3934) );
	vdp_slatch g4095 (.Q(w3949), .D(w3948), .C(w3933), .nC(w3937) );
	vdp_slatch g4096 (.Q(w3947), .D(w3959), .C(w3939), .nC(w3934) );
	vdp_slatch g4097 (.Q(w3946), .D(w4006), .C(w3933), .nC(w3937) );
	vdp_slatch g4098 (.Q(w3945), .D(w3944), .C(w3939), .nC(w3934) );
	vdp_slatch g4099 (.Q(w4032), .D(w3943), .C(w3933), .nC(w3937) );
	vdp_slatch g4100 (.Q(w3941), .D(w4021), .C(w3939), .nC(w3934) );
	vdp_slatch g4101 (.Q(w3940), .D(w3938), .C(w3933), .nC(w3937) );
	vdp_slatch g4102 (.Q(w4133), .D(w612), .C(w3990), .nC(w3989) );
	vdp_aon22 g4103 (.Z(w3979), .A1(w3982), .B1(w3998), .A2(w4000), .B2(w4133) );
	vdp_slatch g4104 (.Q(w4002), .D(w685), .C(w3990), .nC(w3989) );
	vdp_aon22 g4105 (.Z(w3983), .A1(w3975), .B1(w3998), .A2(w4000), .B2(w4002) );
	vdp_slatch g4106 (.Q(w4132), .D(w698), .C(w3990), .nC(w3989) );
	vdp_aon22 g4107 (.Z(w3974), .A1(w4001), .B1(w3998), .A2(w4000), .B2(w4132) );
	vdp_slatch g4108 (.Q(w4003), .D(w719), .C(w3990), .nC(w3989) );
	vdp_aon22 g4109 (.Z(w3968), .A1(w3967), .B1(w3998), .A2(w4000), .B2(w4003) );
	vdp_slatch g4110 (.Q(w4004), .D(w725), .C(w3990), .nC(w3989) );
	vdp_aon22 g4111 (.Z(w3964), .A1(w3963), .B1(w3998), .A2(w4000), .B2(w4004) );
	vdp_slatch g4112 (.Q(w4030), .D(w681), .C(w3990), .nC(w3989) );
	vdp_aon22 g4113 (.Z(w3962), .A1(w3955), .B1(w3998), .A2(w4000), .B2(w4030) );
	vdp_slatch g4114 (.Q(w4131), .D(w661), .C(w3990), .nC(w3989) );
	vdp_aon22 g4115 (.Z(w3954), .A1(w3951), .B1(w3998), .A2(w4000), .B2(w4131) );
	vdp_slatch g4116 (.Q(w4005), .D(w617), .C(w3990), .nC(w3989) );
	vdp_aon22 g4117 (.Z(w3952), .A1(w3948), .B1(w3998), .A2(w4000), .B2(w4005) );
	vdp_aon22 g4118 (.Z(w3959), .A1(w4006), .B1(w3998), .A2(w4000), .B2(1'b0) );
	vdp_aon22 g4119 (.Z(w3944), .A1(w3943), .B1(w3998), .A2(w4000), .B2(1'b0) );
	vdp_aon22 g4120 (.Z(w4021), .A1(w3938), .B1(w3998), .A2(w4000), .B2(1'b0) );
	vdp_notif0 g4121 (.nZ(RD_DATA[2]), .A(w4022), .nE(w3994) );
	vdp_slatch g4122 (.nQ(w4022), .D(w3938), .C(w3993), .nC(w3992) );
	vdp_notif0 g4123 (.nZ(RD_DATA[1]), .A(w4007), .nE(w3994) );
	vdp_slatch g4124 (.nQ(w4007), .D(w3943), .C(w3993), .nC(w3992) );
	vdp_notif0 g4125 (.nZ(RD_DATA[0]), .A(w4156), .nE(w3994) );
	vdp_slatch g4126 (.nQ(w4156), .D(w4006), .C(w3993), .nC(w3992) );
	vdp_notif0 g4127 (.nZ(AD_DATA[7]), .A(w4451), .nE(w3994) );
	vdp_slatch g4128 (.nQ(w4451), .D(w3948), .C(w3993), .nC(w3992) );
	vdp_notif0 g4129 (.nZ(AD_DATA[6]), .A(w4008), .nE(w3994) );
	vdp_slatch g4130 (.nQ(w4008), .D(w3951), .C(w3993), .nC(w3992) );
	vdp_notif0 g4131 (.nZ(AD_DATA[5]), .A(w4009), .nE(w3994) );
	vdp_slatch g4132 (.nQ(w4009), .D(w3955), .C(w3993), .nC(w3992) );
	vdp_notif0 g4133 (.nZ(AD_DATA[4]), .A(w4010), .nE(w3994) );
	vdp_slatch g4134 (.nQ(w4010), .D(w3963), .C(w3993), .nC(w3992) );
	vdp_notif0 g4135 (.nZ(AD_DATA[3]), .A(w4019), .nE(w3994) );
	vdp_slatch g4136 (.nQ(w4019), .D(w3967), .C(w3993), .nC(w3992) );
	vdp_notif0 g4137 (.nZ(AD_DATA[2]), .A(w4017), .nE(w3994) );
	vdp_slatch g4138 (.nQ(w4017), .D(w4001), .C(w3993), .nC(w3992) );
	vdp_notif0 g4139 (.nZ(AD_DATA[1]), .A(w4012), .nE(w3994) );
	vdp_slatch g4140 (.nQ(w4012), .D(w3975), .C(w3993), .nC(w3992) );
	vdp_notif0 g4141 (.nZ(AD_DATA[0]), .A(w4016), .nE(w3994) );
	vdp_slatch g4142 (.nQ(w4016), .D(w3982), .C(w3993), .nC(w3992) );
	vdp_sr_bit g4143 (.Q(w4015), .D(w3721), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4144 (.Q(w4023), .D(w4027), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4145 (.Q(w4027), .D(RD_DATA[0]), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4146 (.Q(w4155), .D(w3979), .C(w3939), .nC(w3934) );
	vdp_comp_strong g4147 (.Z(w3939), .nZ(w3934), .A(w3997) );
	vdp_comp_strong g4148 (.Z(w3933), .nZ(w3937), .A(w3995) );
	vdp_comp_strong g4149 (.Z(w3990), .nZ(w3989), .A(w87) );
	vdp_sr_bit g4150 (.Q(w3935), .D(w4136), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_comp_strong g4151 (.Z(w3993), .nZ(w3992), .A(w4014) );
	vdp_not g4152 (.nZ(w3994), .A(w4015) );
	vdp_and g4153 (.Z(w4014), .A(w3721), .B(HCLK1) );
	vdp_and g4154 (.Z(w3950), .A(w4158), .B(w3935) );
	vdp_and g4155 (.Z(w3953), .A(w4157), .B(w3935) );
	vdp_and g4156 (.Z(w3960), .A(w4146), .B(w3935) );
	vdp_and g4157 (.Z(w3966), .A(w4147), .B(w3935) );
	vdp_and g4158 (.Z(w3969), .A(w4148), .B(w3935) );
	vdp_and g4159 (.Z(w3973), .A(w4149), .B(w3935) );
	vdp_and g4160 (.Z(w4033), .A(w4150), .B(w3935) );
	vdp_and g4161 (.Z(w3977), .A(w4155), .B(w3935) );
	vdp_not g4162 (.nZ(w4135), .A(w4134) );
	vdp_not g4163 (.nZ(w3995), .A(w3996) );
	vdp_not g4164 (.nZ(w3909), .A(w3908) );
	vdp_not g4165 (.nZ(w3913), .A(w3651) );
	vdp_not g4166 (.nZ(w3912), .A(w3656) );
	vdp_not g4167 (.nZ(w3890), .A(w4137) );
	vdp_not g4168 (.nZ(w3889), .A(w4138) );
	vdp_not g4169 (.nZ(w3891), .A(w4141) );
	vdp_not g4170 (.nZ(w4084), .A(M5) );
	vdp_not g4171 (.nZ(w3929), .A(w4083) );
	vdp_aon22 g4172 (.Z(w3917), .A1(w3896), .B1(w3904), .A2(w3923), .B2(w3899) );
	vdp_aon22 g4173 (.Z(w3921), .A1(w3896), .B1(w3923), .A2(w3920), .B2(w3899) );
	vdp_ha g4174 (.CO(w3925), .SUM(w3895), .B(w3924), .A(w3921) );
	vdp_aon222 g4175 (.A1(w3891), .B1(w3889), .C1(w3890), .A2(w3919), .B2(w3918), .C2(w3895), .Z(w3870) );
	vdp_aon22 g4176 (.Z(w4082), .A1(w3896), .B1(w3920), .A2(w3931), .B2(w3899) );
	vdp_ha g4177 (.SUM(w3894), .B(w3925), .A(w4082) );
	vdp_aon222 g4178 (.A1(w3891), .B1(w3889), .C1(w3890), .A2(w3918), .B2(w3895), .C2(w3894), .Z(w3872) );
	vdp_ha g4179 (.CO(w3924), .SUM(w3918), .B(w3917), .A(w3928) );
	vdp_aon222 g4180 (.A1(w3891), .B1(w3889), .C1(w3890), .A2(w3915), .B2(w3919), .C2(w3918), .Z(w3869) );
	vdp_aon22 g4181 (.Z(w3919), .A1(w3896), .B1(w3905), .A2(w3904), .B2(w3899) );
	vdp_aon222 g4182 (.A1(w3891), .B1(w3889), .C1(w3890), .A2(w4042), .B2(w3915), .C2(w3919), .Z(w3866) );
	vdp_aon222 g4183 (.A1(w3891), .B1(w3889), .C1(w3890), .A2(w3914), .B2(w3914), .C2(w3915), .Z(w3650) );
	vdp_aon22 g4184 (.Z(w3915), .A1(w3896), .B1(w3566), .A2(w3905), .B2(w3899) );
	vdp_comp_we g4185 (.Z(w4000), .nZ(w3998), .A(M5) );
	vdp_comp_we g4186 (.Z(w3896), .nZ(w3899), .A(w1) );
	vdp_and g4187 (.Z(w3928), .A(w3929), .B(w4084) );
	vdp_aon222 g4188 (.A1(w3891), .B1(w3889), .C1(w3890), .A2(w3895), .B2(w3894), .C2(w3892), .Z(w3877) );
	vdp_aon222 g4189 (.A1(w3891), .B1(w3889), .C1(w3890), .A2(w3894), .B2(w3892), .C2(w4081), .Z(w3888) );
	vdp_aon22 g4190 (.Z(w3893), .A1(w3896), .B1(w3897), .A2(w3898), .B2(w3899) );
	vdp_aon22 g4191 (.Z(w3916), .A1(w3896), .B1(w3931), .A2(w3897), .B2(w3899) );
	vdp_and g4192 (.Z(w3892), .B(w3916), .A(w3926) );
	vdp_and g4193 (.Z(w4081), .B(w3893), .A(w3927) );
	vdp_oai21 g4194 (.Z(w3908), .A1(w44), .A2(w3980), .B(M5) );
	vdp_aoi21 g4195 (.Z(w3996), .A1(HCLK1), .A2(w16), .B(w103) );
	vdp_oai211 g4196 (.Z(w4134), .A1(HCLK1), .A2(w4), .B(w5), .C(M5) );
	vdp_or g4197 (.Z(w3997), .A(w103), .B(w4135) );
	vdp_nand3 g4198 (.Z(w4136), .A(w95), .B(HPOS[6]), .C(HPOS[7]) );
	vdp_nand g4199 (.Z(w4141), .A(w3656), .B(w3651) );
	vdp_nand g4200 (.Z(w4138), .A(w3651), .B(w3912) );
	vdp_nand g4201 (.Z(w4137), .A(w3912), .B(w3913) );
	vdp_aoi31 g4202 (.Z(w4083), .B3(w4082), .B2(w3921), .B1(w3917), .A(w3916) );
	vdp_slatch g4203 (.Q(w3599), .D(S[0]), .C(w3561), .nC(w3174) );
	vdp_slatch g4204 (.Q(w3601), .D(S[1]), .C(w3561), .nC(w3174) );
	vdp_slatch g4205 (.Q(w3621), .D(S[2]), .C(w3561), .nC(w3174) );
	vdp_slatch g4206 (.Q(w3605), .D(S[3]), .C(w3561), .nC(w3174) );
	vdp_slatch g4207 (.Q(w3607), .D(S[4]), .C(w3561), .nC(w3174) );
	vdp_slatch g4208 (.Q(w3608), .D(S[5]), .C(w3561), .nC(w3174) );
	vdp_slatch g4209 (.Q(w3610), .D(S[6]), .C(w3561), .nC(w3174) );
	vdp_slatch g4210 (.Q(w3612), .D(S[7]), .C(w3561), .nC(w3174) );
	vdp_slatch g4211 (.Q(w3614), .D(S[0]), .C(w3556), .nC(w3555) );
	vdp_slatch g4212 (.Q(w3617), .D(S[1]), .C(w3556), .nC(w3555) );
	vdp_slatch g4213 (.Q(w3618), .D(S[2]), .C(w3556), .nC(w3555) );
	vdp_slatch g4214 (.Q(w3121), .D(S[3]), .C(w3556), .nC(w3555) );
	vdp_slatch g4215 (.Q(w3625), .D(S[4]), .C(w3556), .nC(w3555) );
	vdp_slatch g4216 (.Q(w3097), .D(S[5]), .C(w3556), .nC(w3555) );
	vdp_slatch g4217 (.Q(w3099), .D(S[6]), .C(w3556), .nC(w3555) );
	vdp_slatch g4218 (.Q(w3126), .D(S[7]), .C(w3556), .nC(w3555) );
	vdp_comp_strong g4219 (.Z(w3556), .nZ(w3555), .A(w3310) );
	vdp_comp_strong g4220 (.Z(w3561), .nZ(w3174), .A(w3311) );
	vdp_comp_strong g4221 (.Z(w3562), .nZ(w3623), .A(w3312) );
	vdp_slatch g4222 (.Q(w4116), .D(S[7]), .C(w3562), .nC(w3623) );
	vdp_slatch g4223 (.Q(w4115), .D(S[6]), .C(w3562), .nC(w3623) );
	vdp_slatch g4224 (.Q(w4114), .D(S[5]), .C(w3562), .nC(w3623) );
	vdp_slatch g4225 (.Q(w3628), .D(S[4]), .C(w3562), .nC(w3623) );
	vdp_slatch g4226 (.Q(w3629), .D(S[3]), .C(w3562), .nC(w3623) );
	vdp_slatch g4227 (.Q(w3594), .D(S[2]), .C(w3562), .nC(w3623) );
	vdp_slatch g4228 (.Q(w3592), .D(S[1]), .C(w3562), .nC(w3623) );
	vdp_slatch g4229 (.Q(w3590), .D(S[0]), .C(w3562), .nC(w3623) );
	vdp_slatch g4230 (.Q(w3587), .D(S[7]), .C(w3563), .nC(w3624) );
	vdp_slatch g4231 (.Q(w3588), .D(S[6]), .C(w3563), .nC(w3624) );
	vdp_slatch g4232 (.Q(w3586), .D(S[5]), .C(w3563), .nC(w3624) );
	vdp_slatch g4233 (.Q(w3585), .D(S[4]), .C(w3563), .nC(w3624) );
	vdp_slatch g4234 (.Q(w3583), .D(S[3]), .C(w3563), .nC(w3624) );
	vdp_slatch g4235 (.Q(w3581), .D(S[2]), .C(w3563), .nC(w3624) );
	vdp_slatch g4236 (.Q(w3579), .D(S[1]), .C(w3563), .nC(w3624) );
	vdp_slatch g4237 (.Q(w3576), .D(S[0]), .C(w3563), .nC(w3624) );
	vdp_sr_bit g4238 (.Q(w4145), .D(w3557), .C1(HCLK2), .C2(HCLK1), .nC2(nHCLK1), .nC1(nHCLK2) );
	vdp_sr_bit g4239 (.Q(w3564), .D(w4113), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and g4240 (.Z(w4113), .A(w14), .B(M5) );
	vdp_not g4241 (.nZ(w4111), .A(w3564) );
	vdp_aon22 g4242 (.Z(w3125), .A1(w4116), .B1(w3628), .A2(w3627), .B2(w4074) );
	vdp_aon22 g4243 (.Z(w3122), .A1(w4115), .B1(1'b0), .A2(w3627), .B2(w4074) );
	vdp_aon22 g4244 (.Z(w3626), .A1(w3628), .B1(w3594), .A2(w3627), .B2(w4074) );
	vdp_aon22 g4245 (.Z(w3095), .A1(w3629), .B1(w3592), .A2(w3627), .B2(w4074) );
	vdp_aon22 g4246 (.Z(w3098), .A1(w4114), .B1(w3629), .A2(w3627), .B2(w4074) );
	vdp_comp_strong g4247 (.Z(w3563), .nZ(w3624), .A(w3313) );
	vdp_comp_we g4248 (.Z(w3627), .nZ(w4074), .A(M5) );
	vdp_aon22 g4249 (.Z(w3568), .A1(w3625), .B1(w3626), .A2(w3564), .B2(w4111) );
	vdp_sr_bit g4250 (.Q(w4024), .D(FIFOo[0]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4251 (.Q(w4028), .D(FIFOo[1]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4252 (.Q(w4026), .D(FIFOo[2]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4253 (.Q(w4025), .D(FIFOo[3]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4254 (.Q(w4013), .D(FIFOo[4]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4255 (.Q(w4011), .D(FIFOo[5]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4256 (.Q(w4018), .D(FIFOo[6]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4257 (.Q(w4020), .D(FIFOo[7]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_aon22 g4258 (.Z(w1413), .B1(w4494), .A1(w1441), .B2(w4512), .A2(w43) );
	vdp_not g4259 (.nZ(w4512), .A(w43) );
	vdp_not g4260 (.nZ(w4484), .A(w4471) );
	vdp_not g4261 (.nZ(w4483), .A(w4484) );
	vdp_not g4262 (.nZ(w4482), .A(w4483) );
	vdp_not g4263 (.nZ(w4481), .A(w4482) );
	vdp_and g4264 (.Z(w4494), .B(w4485), .A(w4489) );
	vdp_not g4265 (.nZ(w4485), .A(w4488) );
	vdp_not g4266 (.nZ(w4488), .A(w4487) );
	vdp_not g4267 (.nZ(w4487), .A(w4486) );
	vdp_not g4268 (.nZ(w4486), .A(w4489) );
	vdp_or g4269 (.Z(w4489), .B(w4469), .A(w4468) );
	vdp_dff g4270 (.Q(w4469), .R(w4458), .D(w4468), .C(w4467) );
	vdp_not g4271 (.nZ(w4467), .A(w4490) );
	vdp_nor g4272 (.Z(w4466), .B(w4491), .A(w4468) );
	vdp_dff g4273 (.Q(w4468), .R(w4458), .D(w4491), .C(w4490) );
	vdp_dff g4274 (.Q(w4491), .R(w4458), .D(w4466), .C(w4490) );
	vdp_not g4275 (.nZ(w4490), .A(w4477) );
	vdp_not g4276 (.nZ(w4464), .A(w4477) );
	vdp_dff g4277 (.Q(w4461), .R(w4458), .D(w4492), .C(w4460) );
	vdp_dff g4278 (.Q(w4492), .R(w4458), .D(w4459), .C(w4457) );
	vdp_not g4279 (.nZ(w4457), .A(w4500) );
	vdp_dff g4280 (.Q(w4459), .R(w4458), .D(w4478), .C(w4457) );
	vdp_not g4281 (.nZ(w4460), .A(w4457) );
	vdp_nor g4282 (.Z(w4519), .B(w4495), .A(w4496) );
	vdp_nor g4283 (.Z(w4497), .B(w4495), .A(H40) );
	vdp_not g4284 (.nZ(w4496), .A(H40) );
	vdp_not g4285 (.nZ(w4472), .A(w1205) );
	vdp_AOI222 g4286 (.Z(w4465), .B1(w4499), .A1(w4498), .B2(w4519), .A2(w4495), .C1(w4464), .C2(w4497) );
	vdp_not g4287 (.nZ(EDCLK_O), .A(w4465) );
	vdp_or g4288 (.Z(w4493), .B(w4461), .A(w4492) );
	vdp_nor g4289 (.Z(w4478), .B(w4459), .A(w4492) );
	vdp_not g4290 (.nZ(w4454), .A(w4518) );
	vdp_nand g4291 (.Z(w4473), .B(w4454), .A(w4453) );
	vdp_SR_bit g4292 (.Q(w4518), .D(w4453), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_not g4293 (.nZ(w4517), .A(w4503) );
	vdp_not g4294 (.nZ(w1170), .A(w4516) );
	vdp_not g4295 (.nZ(SYSRES), .A(w4517) );
	vdp_comp_DFF g4296 (.Q(w4453), .D(w4503), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_not g4297 (.nZ(w4513), .A(w4514) );
	vdp_not g4298 (.nZ(w4458), .A(w4515) );
	vdp_not g4299 (.nZ(w4502), .A(w4501) );
	vdp_nand g4300 (.Z(w4515), .B(w4502), .A(w4456) );
	vdp_not g4301 (.nZ(w4500), .A(w4504) );
	vdp_nand g4302 (.Z(w4507), .B(w4506), .A(w4505) );
	vdp_not g4303 (.nZ(w4477), .A(w4462) );
	vdp_nand g4304 (.Z(w4510), .B(w4509), .A(w4508) );
	vdp_not g4305 (.nZ(w4471), .A(w4476) );
	vdp_not g4306 (.nZ(RES), .A(w4473) );
	vdp_dff g4307 (.Q(w4456), .R(1'b0), .D(w4503), .C(w4474) );
	vdp_dff g4308 (.Q(w4501), .R(1'b0), .D(w4456), .C(w4474) );
	vdp_dff g4309 (.Q(w4514), .R(w4458), .D(w4504), .C(w4474) );
	vdp_dff g4310 (.Q(w4504), .R(w4458), .D(w4513), .C(w4474) );
	vdp_dff g4311 (.Q(w4505), .R(w4458), .D(w4462), .C(w4474) );
	vdp_dff g4312 (.Q(w4506), .R(w4458), .D(w4505), .C(w4474) );
	vdp_dff g4313 (.Q(w4462), .R(w4458), .D(w4507), .C(w4474) );
	vdp_dff g4314 (.Q(w4508), .R(w4458), .D(w4476), .C(w4474) );
	vdp_dff g4315 (.Q(w4509), .R(w4458), .D(w4508), .C(w4474) );
	vdp_dff g4316 (.Q(w4511), .R(w4458), .D(w4510), .C(w4474) );
	vdp_dff g4317 (.Q(w4476), .R(w4458), .D(w4511), .C(w4474) );
	vdp_not g4318 (.nZ(w4499), .A(w4500) );
	vdp_nand g4319 (.Z(w4503), .B(w1442), .A(w4516) );
	vdp_not g4320 (.nZ(68K CPU CLOCK), .A(w4470) );
	vdp_or g4321 (.Z(w4495), .B(w43), .A(w1151) );
	vdp_aon22 g4322 (.Z(w4463), .B1(w4493), .A1(w4494), .B2(w1205), .A2(w4472) );
	vdp_or g4323 (.Z(w4470), .B(w4481), .A(w4471) );
	vdp_comp_we g4324 (.A(w2650), .nZ(nHCLK2), .Z(HCLK2) );
	vdp_comp_we g4325 (.A(w2649), .nZ(nHCLK1), .Z(HCLK1) );
	vdp_comp_we g4326 (.A(w4527), .nZ(nDCLK2), .Z(DCLK2) );
	vdp_comp_we g4327 (.A(EDCLK_O), .nZ(nDCLK1), .Z(DCLK1) );
	vdp_not g4328 (.nZ(w4527), .A(EDCLK_O) );
	vdp_sr_bit g4329 (.Q(w4625), .D(w4624), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4330 (.Q(w4643), .D(w4620), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4331 (.Q(w4620), .D(w4605), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4332 (.Q(w4605), .D(w4597), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4333 (.Q(w4600), .D(w6578), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4334 (.Q(w6578), .D(w6579), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4335 (.Q(w6579), .D(w6581), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4336 (.Q(w6581), .D(w6580), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4337 (.Q(w6580), .D(w6582), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4338 (.Q(w6582), .D(w6583), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4339 (.Q(w6583), .D(w6585), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4340 (.Q(w6585), .D(w6584), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4341 (.Q(w6584), .D(w6412), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4342 (.Q(w6412), .D(w4543), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4343 (.Q(w4581), .D(w4582), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4344 (.Q(w4582), .D(w24), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4345 (.Q(w4579), .D(w6586), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4346 (.Q(w4548), .D(w4578), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4347 (.Q(w4547), .D(w6574), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4348 (.Q(w6274), .D(w4627), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4349 (.Q(w4626), .D(w6587), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4350 (.Q(w4628), .D(w4618), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4351 (.Q(w6576), .D(w4), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4352 (.Q(w4568), .D(w4590), .nC(w4593), .C(w4594) );
	vdp_slatch g4353 (.Q(w4572), .D(w4591), .nC(w4593), .C(w4594) );
	vdp_slatch g4354 (.Q(w4560), .D(w4592), .nC(w4593), .C(w4594) );
	vdp_slatch g4355 (.Q(w4551), .D(w4598), .nC(w4593), .C(w4594) );
	vdp_slatch g4356 (.Q(w4550), .D(w4589), .nC(w4593), .C(w4594) );
	vdp_slatch g4357 (.Q(w4549), .D(w4588), .nC(w4593), .C(w4594) );
	vdp_slatch g4358 (.Q(w4602), .D(w4587), .nC(w4593), .C(w4594) );
	vdp_slatch g4359 (.Q(w4552), .D(w4585), .nC(w4593), .C(w4594) );
	vdp_slatch g4360 (.Q(w4556), .D(w4586), .nC(w4593), .C(w4594) );
	vdp_slatch g4361 (.Q(w4557), .D(w4584), .nC(w4593), .C(w4594) );
	vdp_comp_str g4362 (.nZ(w4593), .A(w4599), .Z(w4594) );
	vdp_sr_bit g4363 (.Q(w4621), .D(w4644), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4364 (.Q(w6260), .D(w7), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_xor g4365 (.Z(w4566), .B(w4558), .A(w4569) );
	vdp_xor g4366 (.Z(w4561), .B(w4559), .A(w4567) );
	vdp_xor g4367 (.Z(w4563), .B(w4545), .A(w4560) );
	vdp_xor g4368 (.Z(w6363), .B(w4545), .A(w4551) );
	vdp_xor g4369 (.Z(w6364), .B(w4545), .A(w4550) );
	vdp_xor g4370 (.Z(w6359), .B(w4545), .A(w4549) );
	vdp_aon22 g4371 (.Z(w6360), .B2(w4573), .B1(w4568), .A1(w4566), .A2(w4562) );
	vdp_aon22 g4372 (.Z(w6361), .B2(w4573), .B1(w4566), .A1(w4561), .A2(w4562) );
	vdp_aon22 g4373 (.Z(w6362), .B2(w4573), .B1(w4561), .A1(w4563), .A2(w4562) );
	vdp_aon22 g4374 (.Z(w4564), .B2(w4555), .B1(w4560), .A1(w4572), .A2(w4565) );
	vdp_aon22 g4375 (.Z(w4570), .B2(w4555), .B1(w4572), .A1(w4568), .A2(w4565) );
	vdp_aon22 g4376 (.Z(w4636), .B2(w4629), .B1(w4632), .A1(w4633), .A2(w80) );
	vdp_aon22 g4377 (.Z(w4637), .B2(w4631), .B1(w4632), .A1(w4633), .A2(w79) );
	vdp_aon22 g4378 (.Z(w4638), .B2(w4630), .B1(w4632), .A1(w4633), .A2(w78) );
	vdp_aon22 g4379 (.Z(w4639), .B2(w4634), .B1(w4632), .A1(w4633), .A2(w77) );
	vdp_aon22 g4380 (.Z(w4640), .B2(w4635), .B1(w4632), .A1(w4633), .A2(w76) );
	vdp_not g4381 (.nZ(w4606), .A(w4543) );
	vdp_not g4382 (.nZ(w4576), .A(w4610) );
	vdp_not g4383 (.nZ(w4609), .A(w125) );
	vdp_not g4384 (.nZ(w4614), .A(w4612) );
	vdp_not g4385 (.nZ(w4601), .A(M5) );
	vdp_not g4386 (.nZ(w4642), .A(w81) );
	vdp_not g4387 (.nZ(w4641), .A(w82) );
	vdp_not g4388 (.nZ(w4616), .A(1'b0) );
	vdp_not g4389 (.nZ(w4617), .A(M5) );
	vdp_not g4390 (.nZ(w4542), .A(w4543) );
	vdp_not g4391 (.nZ(w4546), .A(w4577) );
	vdp_not g4392 (.nZ(w4553), .A(w4557) );
	vdp_not g4393 (.nZ(w4559), .A(w4596) );
	vdp_and g4394 (.Z(w4597), .B(w4606), .A(w4607) );
	vdp_and g4395 (.Z(w4611), .B(w4609), .A(w4620) );
	vdp_or g4396 (.Z(w4608), .B(w4611), .A(w4623) );
	vdp_or g4397 (.Z(w4604), .B(w4646), .A(w4611) );
	vdp_and g4398 (.Z(w4622), .B(w4615), .A(1'b0) );
	vdp_and g4399 (.Z(w4645), .B(w4615), .A(w4616) );
	vdp_or g4400 (.Z(w4644), .B(w7), .A(w27) );
	vdp_and g4401 (.Z(w127), .B(w6735), .A(w4) );
	vdp_and g4402 (.Z(w6574), .B(w4542), .A(w4544) );
	vdp_or g4403 (.Z(w4595), .B(w4548), .A(w4547) );
	vdp_and g4404 (.Z(w4558), .B(w4552), .A(w4545) );
	vdp_comp_we g4405 (.nZ(w4555), .A(w1), .Z(w4565) );
	vdp_comp_we g4406 (.nZ(w4573), .A(w1), .Z(w4562) );
	vdp_comp_we g4407 (.nZ(w4632), .A(w125), .Z(w4633) );
	vdp_not g4408 (.nZ(w4654), .A(w4624) );
	vdp_rs_FF g4409 (.Q(w6575), .R(w6576), .S(w4595) );
	vdp_rs_FF g4410 (.Q(w6735), .R(w6576), .S(w4547) );
	vdp_ha g4411 (.SUM(w4569), .B(w4570), .A(w4571) );
	vdp_ha g4412 (.SUM(w4567), .B(w4564), .A(w4554), .CO(w4571) );
	vdp_not g4413 (.nZ(w4580), .A(w4541) );
	vdp_and g4414 (.Z(w4583), .B(w4543), .A(w4544) );
	vdp_and3 g4415 (.Z(w4554), .B(w4552), .A(w4545), .C(w4553) );
	vdp_and3 g4416 (.Z(w4627), .B(w4625), .A(M5), .C(w4654) );
	vdp_and3 g4417 (.Z(w6587), .B(w4630), .A(w4629), .C(w4628) );
	vdp_and3 g4418 (.Z(w4646), .B(w82), .A(w4642), .C(w118) );
	vdp_and3 g4419 (.Z(w6577), .B(w81), .A(w4641), .C(w118) );
	vdp_and3 g4420 (.Z(w4623), .B(w4642), .A(w4641), .C(w118) );
	vdp_or3 g4421 (.Z(w4603), .B(w6577), .A(w4611), .C(w4614) );
	vdp_and3 g4422 (.Z(w4599), .B(HCLK1), .A(w4581), .C(DCLK1) );
	vdp_or3 g4423 (.Z(w4615), .B(w4618), .A(w4643), .C(w4617) );
	vdp_oai21 g4424 (.Z(w4596), .B(w4545), .A1(w4552), .A2(w4557) );
	vdp_nor g4425 (.Z(w4541), .B(w4583), .A(w4582) );
	vdp_nor g4426 (.Z(w6586), .B(w4546), .A(w6575) );
	vdp_nand g4427 (.Z(w4619), .B(w4601), .A(w4600) );
	vdp_nand g4428 (.Z(w4575), .B(w4642), .A(w4641) );
	vdp_nand g4429 (.Z(w4610), .B(w81), .A(w4641) );
	vdp_nand g4430 (.Z(w4574), .B(w82), .A(w4642) );
	vdp_nor g4431 (.Z(w4624), .B(w4626), .A(w4539) );
	vdp_cnt_bit_rev g4432 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4629), .CI(w4658), .B(w4621), .A(w4622) );
	vdp_cnt_bit_rev g4433 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4631), .CI(w4657), .B(w4621), .A(w4622), .CO(w4658) );
	vdp_cnt_bit_rev g4434 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4630), .CI(w4656), .B(w4621), .A(w4622), .CO(w4657) );
	vdp_cnt_bit_rev g4435 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4634), .CI(w4655), .B(w4621), .A(w4622), .CO(w4656) );
	vdp_cnt_bit_rev g4436 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4635), .CI(w4645), .B(w4621), .A(w4622), .CO(w4655) );
	vdp_cnt_bit_load g4437 (.Q(w4665), .D(w4705), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4667), .CI(w6638), .L(w4706), .nL(w4671) );
	vdp_cnt_bit_load g4438 (.Q(w4668), .D(w4710), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4667), .CI(w6637), .L(w4706), .nL(w4671), .CO(w6638) );
	vdp_cnt_bit_load g4439 (.Q(w4670), .D(w4711), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4667), .CI(w6636), .L(w4706), .nL(w4671), .CO(w6637) );
	vdp_cnt_bit_load g4440 (.Q(w4672), .D(w4735), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4667), .CI(w6635), .L(w4706), .nL(w4671), .CO(w6636) );
	vdp_cnt_bit_load g4441 (.Q(w4676), .D(w4736), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4667), .CI(w6634), .L(w4706), .nL(w4671), .CO(w6635) );
	vdp_cnt_bit_load g4442 (.Q(w4673), .D(w4737), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4667), .CI(w6633), .L(w4706), .nL(w4671), .CO(w6634) );
	vdp_cnt_bit_load g4443 (.Q(w4669), .D(w4738), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4667), .CI(w4666), .L(w4706), .nL(w4671), .CO(w6633) );
	vdp_fa g4444 (.SUM(w4813), .CO(w6648), .CI(1'b1), .A(w4867), .B(w4816) );
	vdp_fa g4445 (.SUM(w4815), .CO(w6649), .CI(w6648), .A(w4866), .B(w4820) );
	vdp_fa g4446 (.SUM(w4821), .CO(w6650), .CI(w6649), .A(w4865), .B(w4824) );
	vdp_fa g4447 (.SUM(w4823), .CO(w6651), .CI(w6650), .A(w4864), .B(w4826) );
	vdp_fa g4448 (.SUM(w4828), .CO(w6652), .CI(w6651), .A(w4863), .B(w4830) );
	vdp_fa g4449 (.SUM(w4834), .CO(w6653), .CI(w6652), .A(w4862), .B(w4858) );
	vdp_fa g4450 (.SUM(w4837), .CO(w6654), .CI(w6653), .A(w4860), .B(w4836) );
	vdp_fa g4451 (.SUM(w4841), .CO(w6655), .CI(w6654), .A(w4872), .B(w4840) );
	vdp_fa g4452 (.SUM(w4843), .CO(w6656), .CI(w6655), .A(w4873), .B(w4842) );
	vdp_fa g4453 (.SUM(w4856), .CI(w6656), .A(w4877), .B(w4855) );
	vdp_fa g4454 (.SUM(w4867), .CO(w6639), .CI(1'b0), .A(VPOS[0]), .B(w4868) );
	vdp_fa g4455 (.SUM(w4866), .CO(w6640), .CI(w6639), .A(VPOS[1]), .B(w1) );
	vdp_fa g4456 (.SUM(w4865), .CO(w6641), .CI(w6640), .A(VPOS[2]), .B(1'b0) );
	vdp_fa g4457 (.SUM(w4864), .CO(w6642), .CI(w6641), .A(VPOS[3]), .B(1'b0) );
	vdp_fa g4458 (.SUM(w4863), .CO(w6643), .CI(w6642), .A(VPOS[4]), .B(1'b0) );
	vdp_fa g4459 (.SUM(w4862), .CO(w6644), .CI(w6643), .A(VPOS[5]), .B(1'b0) );
	vdp_fa g4460 (.SUM(w4860), .CO(w6645), .CI(w6644), .A(VPOS[6]), .B(1'b0) );
	vdp_fa g4461 (.SUM(w4872), .CO(w6646), .CI(w6645), .A(VPOS[7]), .B(w4868) );
	vdp_fa g4462 (.SUM(w4873), .CO(w6647), .CI(w6646), .A(VPOS[8]), .B(w1) );
	vdp_fa g4463 (.SUM(w4877), .CI(w6647), .A(VPOS[9]), .B(1'b0) );
	vdp_slatch g4464 (.nC(w4761), .C(w4760), .Q(w4807), .D(S[0]) );
	vdp_dlatch_inv g4465 (.nQ(w4806), .D(w4774), .nC(nHCLK2), .C(HCLK2) );
	vdp_slatch g4466 (.nC(w4746), .C(w4745), .Q(w4774), .D(w4763) );
	vdp_slatch g4467 (.nC(w4761), .C(w4760), .Q(w4804), .D(S[1]) );
	vdp_slatch g4468 (.nC(w4746), .C(w4745), .Q(w6678), .D(w4765) );
	vdp_slatch g4469 (.nC(w4761), .C(w4760), .Q(w4802), .D(S[2]) );
	vdp_slatch g4470 (.nC(w4746), .C(w4745), .Q(w6679), .D(w4756) );
	vdp_slatch g4471 (.nC(w4761), .C(w4760), .Q(w4800), .D(S[3]) );
	vdp_slatch g4472 (.nC(w4746), .C(w4745), .Q(w6680), .D(w4752) );
	vdp_slatch g4473 (.nC(w4761), .C(w4760), .Q(w4796), .D(S[4]) );
	vdp_slatch g4474 (.nC(w4746), .C(w4745), .Q(w6681), .D(w4748) );
	vdp_slatch g4475 (.nC(w4761), .C(w4760), .Q(w4795), .D(S[5]) );
	vdp_slatch g4476 (.nC(w4746), .C(w4745), .Q(w6682), .D(w4744) );
	vdp_slatch g4477 (.nC(w4761), .C(w4760), .Q(w4792), .D(S[6]) );
	vdp_slatch g4478 (.nC(w4746), .C(w4745), .Q(w6683), .D(w6625) );
	vdp_slatch g4479 (.nC(w4761), .C(w4760), .Q(w6684), .D(S[7]) );
	vdp_slatch g4480 (.nC(w4746), .C(w4745), .Q(w6685), .D(w4776) );
	vdp_slatch g4481 (.nC(w4746), .C(w4745), .Q(w4777), .D(w4778) );
	vdp_slatch g4482 (.nC(w4746), .C(w4745), .Q(w6686), .D(w4780) );
	vdp_dlatch_inv g4483 (.nQ(w4803), .D(w6678), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4484 (.nQ(w4801), .D(w6679), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4485 (.nQ(w4798), .D(w6680), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4486 (.nQ(w4797), .D(w6681), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4487 (.nQ(w4794), .D(w6682), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4488 (.nQ(w4791), .D(w6683), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4489 (.nQ(w4790), .D(w6685), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4490 (.nQ(w4789), .D(w4777), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4491 (.nQ(w4779), .D(w6686), .nC(nHCLK2), .C(HCLK2) );
	vdp_sr_bit g4492 (.Q(w4731), .D(w4662), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4493 (.Z(w4577), .B2(w4727), .B1(w4733), .A1(M5), .A2(w4732) );
	vdp_sr_bit g4494 (.Q(w4662), .D(w4728), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4495 (.Q(w6624), .D(w4729), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4496 (.Q(w4729), .D(w4707), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4497 (.Q(w4768), .D(w4770), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4498 (.Q(w4759), .D(w4773), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4499 (.Q(w4755), .D(w4766), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4500 (.Q(w4751), .D(w4767), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4501 (.Q(w4747), .D(w4749), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4502 (.Q(w4743), .D(w4741), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4503 (.Q(w4775), .D(w4742), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4504 (.Q(w6687), .D(w4740), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4505 (.Q(w4689), .D(w4739), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4506 (.Q(w4696), .D(w4734), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4507 (.Q(w4730), .D(w4663), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4508 (.Q(w4663), .D(w4685), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4509 (.Q(w4913), .D(w131), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4510 (.Q(w4915), .D(VRAMA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4511 (.Q(w4685), .D(w9), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4512 (.Q(w4916), .D(w6632), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4513 (.Q(w6632), .D(w4913), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4514 (.Q(w6676), .D(w4899), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4515 (.Q(w6674), .D(w4902), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4516 (.Q(w6672), .D(w4917), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4517 (.Q(w6670), .D(w4879), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4518 (.Q(w6668), .D(w4705), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4519 (.Q(w6666), .D(w4710), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4520 (.Q(w6664), .D(w4711), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4521 (.Q(w6662), .D(w4735), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4522 (.Q(w6660), .D(w4736), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4523 (.Q(w6658), .D(w4737), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4524 (.Q(w4897), .D(w4738), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4525 (.Q(w4889), .D(w6657), .nC(w4888), .C(w4880) );
	vdp_dlatch_inv g4526 (.nQ(w6657), .D(w4897), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4527 (.Q(w4890), .D(w6659), .nC(w4888), .C(w4880) );
	vdp_dlatch_inv g4528 (.nQ(w6659), .D(w6658), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4529 (.Q(w4891), .D(w6661), .nC(w4888), .C(w4880) );
	vdp_dlatch_inv g4530 (.nQ(w6661), .D(w6660), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4531 (.Q(w4892), .D(w6663), .nC(w4888), .C(w4880) );
	vdp_dlatch_inv g4532 (.nQ(w6663), .D(w6662), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4533 (.Q(w4893), .D(w6665), .nC(w4888), .C(w4880) );
	vdp_dlatch_inv g4534 (.nQ(w6665), .D(w6664), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4535 (.Q(w6631), .D(w6667), .nC(w4888), .C(w4880) );
	vdp_dlatch_inv g4536 (.nQ(w6667), .D(w6666), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4537 (.Q(w4894), .D(w6669), .nC(w4888), .C(w4880) );
	vdp_dlatch_inv g4538 (.nQ(w6669), .D(w6668), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4539 (.Q(w4884), .D(w6671), .nC(w4888), .C(w4880) );
	vdp_dlatch_inv g4540 (.nQ(w6671), .D(w6670), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4541 (.Q(w4887), .D(w6673), .nC(w4888), .C(w4880) );
	vdp_dlatch_inv g4542 (.nQ(w6673), .D(w6672), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4543 (.Q(w4885), .D(w6675), .nC(w4888), .C(w4880) );
	vdp_dlatch_inv g4544 (.nQ(w6675), .D(w6674), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4545 (.Q(w4886), .D(w6677), .nC(w4888), .C(w4880) );
	vdp_dlatch_inv g4546 (.nQ(w6677), .D(w6676), .nC(nHCLK1), .C(HCLK1) );
	vdp_aon22 g4547 (.Z(w6431), .B2(w4715), .B1(w4665), .A1(w4664), .A2(w6409) );
	vdp_aon22 g4548 (.Z(w6432), .B2(w4715), .B1(w4668), .A1(w4664), .A2(w4720) );
	vdp_aon22 g4549 (.Z(w6433), .B2(w4715), .B1(w4670), .A1(w4664), .A2(w4719) );
	vdp_aon22 g4550 (.Z(w6434), .B2(w4715), .B1(w4672), .A1(w4664), .A2(w4718) );
	vdp_aon22 g4551 (.Z(w6435), .B2(w4715), .B1(w4676), .A1(w4664), .A2(w4717) );
	vdp_aon22 g4552 (.Z(w6437), .B2(w4715), .B1(w4673), .A1(w4664), .A2(w4716) );
	vdp_aon22 g4553 (.Z(w6436), .B2(w4715), .B1(w4669), .A1(w4664), .A2(w4714) );
	vdp_aon22 g4554 (.Z(w4938), .B2(w4678), .B1(w3), .A1(w4674), .A2(w4669) );
	vdp_aon22 g4555 (.Z(w4827), .B2(w4787), .B1(w4796), .A1(w4797), .A2(w4811) );
	vdp_2x_sr_bit g4556 (.Q(w4726), .D(w4669), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4557 (.Z(w6410), .B2(w4678), .B1(w4726), .A1(w4674), .A2(w4673) );
	vdp_2x_sr_bit g4558 (.Q(w4675), .D(w4673), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4559 (.Z(w4998), .B2(w4678), .B1(w4675), .A1(w4674), .A2(w4676) );
	vdp_2x_sr_bit g4560 (.Q(w4713), .D(w4676), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4561 (.Z(w5004), .B2(w4678), .B1(w4713), .A1(w4674), .A2(w4672) );
	vdp_2x_sr_bit g4562 (.Q(w4677), .D(w4672), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4563 (.Z(w5056), .B2(w4678), .B1(w4677), .A1(w4674), .A2(w4670) );
	vdp_2x_sr_bit g4564 (.Q(w4680), .D(w4670), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4565 (.Z(w5108), .B2(w4678), .B1(w4680), .A1(w4674), .A2(w4668) );
	vdp_aon22 g4566 (.Z(w5123), .B2(w4678), .B1(1'b1), .A1(w4674), .A2(w4665) );
	vdp_aon22 g4567 (.Z(w4763), .B2(w4688), .B1(w4764), .A1(w4691), .A2(w4762) );
	vdp_dlatch_inv g4568 (.nQ(w4762), .D(w4768), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4569 (.nZ(w4764), .A(S[0]) );
	vdp_aon22 g4570 (.Z(w4765), .B2(w4688), .B1(w4758), .A1(w4691), .A2(w4757) );
	vdp_dlatch_inv g4571 (.nQ(w4757), .D(w4759), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4572 (.nZ(w4758), .A(S[1]) );
	vdp_aon22 g4573 (.Z(w4756), .B2(w4688), .B1(w4754), .A1(w4691), .A2(w4753) );
	vdp_dlatch_inv g4574 (.nQ(w4753), .D(w4755), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4575 (.nZ(w4754), .A(S[2]) );
	vdp_aon22 g4576 (.Z(w4752), .B2(w4688), .B1(w4712), .A1(w4691), .A2(w4750) );
	vdp_dlatch_inv g4577 (.nQ(w4750), .D(w4751), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4578 (.nZ(w4712), .A(S[3]) );
	vdp_aon22 g4579 (.Z(w4748), .B2(w4688), .B1(w4708), .A1(w4691), .A2(w4709) );
	vdp_dlatch_inv g4580 (.nQ(w4709), .D(w4747), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4581 (.nZ(w4708), .A(S[4]) );
	vdp_aon22 g4582 (.Z(w4744), .B2(w4688), .B1(w4704), .A1(w4691), .A2(w4703) );
	vdp_dlatch_inv g4583 (.nQ(w4703), .D(w4743), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4584 (.nZ(w4704), .A(S[5]) );
	vdp_aon22 g4585 (.Z(w6625), .B2(w4688), .B1(w4699), .A1(w4691), .A2(w4698) );
	vdp_dlatch_inv g4586 (.nQ(w4698), .D(w4775), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4587 (.nZ(w4699), .A(S[6]) );
	vdp_aon22 g4588 (.Z(w4776), .B2(w4688), .B1(w4692), .A1(w4691), .A2(w4690) );
	vdp_dlatch_inv g4589 (.nQ(w4690), .D(w6687), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4590 (.nZ(w4692), .A(S[7]) );
	vdp_aon22 g4591 (.Z(w4778), .B2(w4688), .B1(w4933), .A1(w4691), .A2(1'b1) );
	vdp_dlatch_inv g4592 (.nQ(w4933), .D(w4689), .nC(nHCLK1), .C(HCLK1) );
	vdp_aon22 g4593 (.Z(w4780), .B2(w4688), .B1(1'b1), .A1(w4691), .A2(w4697) );
	vdp_dlatch_inv g4594 (.nQ(w4697), .D(w4696), .nC(nHCLK1), .C(HCLK1) );
	vdp_sr_bit g4595 (.Q(w4667), .D(w6604), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4596 (.Q(w4679), .D(w30), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4597 (.Q(w4700), .D(w4679), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4598 (.Q(w4684), .D(w5), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4599 (.Q(w4694), .D(w4684), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4600 (.Q(w4707), .D(w6603), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_not g4601 (.nZ(w4702), .A(w4701) );
	vdp_not g4602 (.nZ(w4695), .A(M5) );
	vdp_not g4603 (.nZ(w6604), .A(w4693) );
	vdp_not g4604 (.nZ(w4683), .A(w4694) );
	vdp_not g4605 (.nZ(w6603), .A(w4686) );
	vdp_not g4606 (.nZ(w4681), .A(w4666) );
	vdp_aon22 g4607 (.Z(w4786), .B2(w4782), .B1(w4592), .A1(w4781), .A2(w4591) );
	vdp_aon22 g4608 (.Z(w4785), .B2(w4782), .B1(w4591), .A1(w4781), .A2(w4590) );
	vdp_aon22 g4609 (.Z(w4784), .B2(w4782), .B1(w4590), .A1(w4781), .A2(1'b0) );
	vdp_slatch g4610 (.nQ(w6696), .D(w4912), .nC(w4896), .C(w4901) );
	vdp_aon22 g4611 (.Z(w4912), .B2(w4895), .B1(w4770), .A1(w4900), .A2(w4738) );
	vdp_notif0 g4612 (.A(w6696), .nZ(AD_DATA[0]), .nE(w4906) );
	vdp_slatch g4613 (.nQ(w6695), .D(w4911), .nC(w4896), .C(w4901) );
	vdp_aon22 g4614 (.Z(w4911), .B2(w4895), .B1(w4773), .A1(w4900), .A2(w4737) );
	vdp_notif0 g4615 (.A(w6695), .nZ(AD_DATA[1]), .nE(w4906) );
	vdp_slatch g4616 (.nQ(w6694), .D(w4910), .nC(w4896), .C(w4901) );
	vdp_aon22 g4617 (.Z(w4910), .B2(w4895), .B1(w4766), .A1(w4900), .A2(w4736) );
	vdp_notif0 g4618 (.A(w6694), .nZ(AD_DATA[2]), .nE(w4906) );
	vdp_slatch g4619 (.nQ(w6693), .D(w6629), .nC(w4896), .C(w4901) );
	vdp_aon22 g4620 (.Z(w6629), .B2(w4895), .B1(w4767), .A1(w4900), .A2(w4735) );
	vdp_notif0 g4621 (.A(w6693), .nZ(AD_DATA[3]), .nE(w4906) );
	vdp_slatch g4622 (.nQ(w6692), .D(w6628), .nC(w4896), .C(w4901) );
	vdp_aon22 g4623 (.Z(w6628), .B2(w4895), .B1(w4749), .A1(w4900), .A2(w4711) );
	vdp_notif0 g4624 (.A(w6692), .nZ(AD_DATA[4]), .nE(w4906) );
	vdp_slatch g4625 (.nQ(w6691), .D(w6627), .nC(w4896), .C(w4901) );
	vdp_aon22 g4626 (.Z(w6627), .B2(w4895), .B1(w4741), .A1(w4900), .A2(w4710) );
	vdp_notif0 g4627 (.A(w6691), .nZ(AD_DATA[5]), .nE(w4906) );
	vdp_slatch g4628 (.nQ(w6690), .D(w4909), .nC(w4896), .C(w4901) );
	vdp_aon22 g4629 (.Z(w4909), .B2(w4895), .B1(w4742), .A1(w4900), .A2(w4705) );
	vdp_notif0 g4630 (.A(w6690), .nZ(AD_DATA[6]), .nE(w4906) );
	vdp_slatch g4631 (.nQ(w6689), .D(w4918), .nC(w4896), .C(w4901) );
	vdp_aon22 g4632 (.Z(w4918), .B2(w4895), .B1(w4740), .A1(w4900), .A2(w4879) );
	vdp_notif0 g4633 (.A(w6689), .nZ(AD_DATA[7]), .nE(w4906) );
	vdp_slatch g4634 (.nQ(w4908), .D(w4907), .nC(w4896), .C(w4901) );
	vdp_aon22 g4635 (.Z(w4907), .B2(w4895), .B1(w4739), .A1(w4900), .A2(w4917) );
	vdp_notif0 g4636 (.A(w4908), .nZ(RD_DATA[0]), .nE(w4906) );
	vdp_slatch g4637 (.nQ(w4905), .D(w4904), .nC(w4896), .C(w4901) );
	vdp_aon22 g4638 (.Z(w4904), .B2(w4895), .B1(w4734), .A1(w4900), .A2(w4902) );
	vdp_notif0 g4639 (.A(w4905), .nZ(RD_DATA[1]), .nE(w4906) );
	vdp_slatch g4640 (.nQ(w4903), .D(w4898), .nC(w4896), .C(w4901) );
	vdp_aon22 g4641 (.Z(w4898), .B2(w4895), .B1(1'b0), .A1(w4900), .A2(w4899) );
	vdp_notif0 g4642 (.A(w4903), .nZ(RD_DATA[2]), .nE(w4906) );
	vdp_not g4643 (.nZ(w4906), .A(w4916) );
	vdp_sr_bit g4644 (.Q(w4585), .D(w6700), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4645 (.Q(w4586), .D(w4875), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4646 (.Q(w4871), .D(w4869), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_dlatch_inv g4647 (.nQ(w4870), .D(w4772), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4648 (.nQ(w4869), .D(w4810), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g4649 (.nQ(w4816), .D(w4812), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4650 (.nQ(w6626), .D(w4813), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4651 (.nQ(w4820), .D(w4814), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4652 (.nQ(w4818), .D(w4815), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4653 (.nQ(w4824), .D(w4819), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4654 (.nQ(w4822), .D(w4821), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4655 (.nQ(w4826), .D(w4825), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4656 (.nQ(w4835), .D(w4823), .nC(nHCLK2), .C(HCLK2) );
	vdp_aon22 g4657 (.Z(w4825), .B2(w4787), .B1(w4800), .A1(w4798), .A2(w4811) );
	vdp_aon22 g4658 (.Z(w4819), .B2(w4787), .B1(w4802), .A1(w4801), .A2(w4811) );
	vdp_aon22 g4659 (.Z(w4814), .B2(w4787), .B1(w4804), .A1(w4803), .A2(w4811) );
	vdp_aon22 g4660 (.Z(w4812), .B2(w4787), .B1(w4807), .A1(w4806), .A2(w4811) );
	vdp_not g4661 (.nZ(w4809), .A(w4772) );
	vdp_not g4662 (.nZ(w4588), .A(w6626) );
	vdp_not g4663 (.nZ(w4589), .A(w4818) );
	vdp_not g4664 (.nZ(w4598), .A(w4822) );
	vdp_not g4665 (.nZ(w4592), .A(w4835) );
	vdp_not g4666 (.nZ(w4831), .A(w4827) );
	vdp_not g4667 (.nZ(w4591), .A(w4829) );
	vdp_dlatch_inv g4668 (.nQ(w4830), .D(w4827), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4669 (.nQ(w4829), .D(w4828), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g4670 (.nZ(w4590), .A(w4838) );
	vdp_dlatch_inv g4671 (.nQ(w4858), .D(w4793), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4672 (.nQ(w4838), .D(w4834), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g4673 (.nZ(w4839), .A(w4859) );
	vdp_dlatch_inv g4674 (.nQ(w4836), .D(w4859), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4675 (.nQ(w4848), .D(w4837), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g4676 (.nZ(w4833), .A(w4844) );
	vdp_dlatch_inv g4677 (.nQ(w4840), .D(w4844), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4678 (.nQ(w4849), .D(w4841), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4679 (.nQ(w4842), .D(w4832), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4680 (.nQ(w4846), .D(w4843), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4681 (.nQ(w4855), .D(w4845), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4682 (.nQ(w4857), .D(w4856), .nC(nHCLK2), .C(HCLK2) );
	vdp_sr_bit g4683 (.Q(w4584), .D(w6688), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4684 (.Z(w4845), .B2(w4787), .B1(1'b0), .A1(w4779), .A2(w4811) );
	vdp_aon22 g4685 (.Z(w4832), .B2(w4787), .B1(1'b0), .A1(w4789), .A2(w4811) );
	vdp_aon22 g4686 (.Z(w6688), .B2(w4883), .B1(M5), .A1(w132), .A2(w4929) );
	vdp_not g4687 (.nZ(w4874), .A(w1) );
	vdp_not g4688 (.nZ(w4932), .A(w4886) );
	vdp_not g4689 (.nZ(w4875), .A(w4885) );
	vdp_not g4690 (.nZ(w4930), .A(w4887) );
	vdp_not g4691 (.nZ(w4883), .A(w4884) );
	vdp_not g4692 (.nZ(w4929), .A(M5) );
	vdp_not g4693 (.nZ(w4578), .A(w4881) );
	vdp_not g4694 (.nZ(w4876), .A(w4584) );
	vdp_not g4695 (.nZ(w6697), .A(w4585) );
	vdp_not g4696 (.nZ(w4931), .A(M5) );
	vdp_not g4697 (.nZ(w4847), .A(w1) );
	vdp_not g4698 (.nZ(w4851), .A(w4784) );
	vdp_bufif0 g4699 (.A(1'b0), .Z(VRAMA[0]), .nE(w4681) );
	vdp_bufif0 g4700 (.A(w4669), .Z(VRAMA[1]), .nE(w4681) );
	vdp_bufif0 g4701 (.A(w4673), .Z(VRAMA[2]), .nE(w4681) );
	vdp_bufif0 g4702 (.A(w4676), .Z(VRAMA[3]), .nE(w4681) );
	vdp_bufif0 g4703 (.A(w4672), .Z(VRAMA[4]), .nE(w4681) );
	vdp_bufif0 g4704 (.A(w4670), .Z(VRAMA[5]), .nE(w4681) );
	vdp_bufif0 g4705 (.A(1'b0), .Z(VRAMA[6]), .nE(w4681) );
	vdp_bufif0 g4706 (.A(1'b0), .Z(VRAMA[7]), .nE(w4681) );
	vdp_aon22 g4707 (.Z(w4844), .B2(w4787), .B1(w6684), .A1(w4790), .A2(w4811) );
	vdp_aon22 g4708 (.Z(w4859), .B2(w4787), .B1(w4792), .A1(w4791), .A2(w4811) );
	vdp_aon22 g4709 (.Z(w4793), .B2(w4787), .B1(w4795), .A1(w4794), .A2(w4811) );
	vdp_comp_str g4710 (.A(w4808), .nZ(w4746), .Z(w4745) );
	vdp_and g4711 (.Z(w4771), .B(w4731), .A(w4727) );
	vdp_comp_we g4712 (.A(w4771), .nZ(w4811), .Z(w4787) );
	vdp_comp_str g4713 (.A(w4805), .nZ(w4761), .Z(w4760) );
	vdp_not g4714 (.nZ(w4727), .A(M5) );
	vdp_comp_str g4715 (.A(w4878), .nZ(w4888), .Z(w4880) );
	vdp_comp_str g4716 (.A(w4914), .nZ(w4896), .Z(w4901) );
	vdp_comp_we g4717 (.A(M5), .nZ(w4688), .Z(w4691) );
	vdp_comp_we g4718 (.A(w4723), .nZ(w4715), .Z(w4664) );
	vdp_comp_we g4719 (.A(w4702), .nZ(w4671), .Z(w4706) );
	vdp_comp_we g4720 (.A(M5), .nZ(w4678), .Z(w4674) );
	vdp_comp_we g4721 (.A(w1), .nZ(w4782), .Z(w4781) );
	vdp_comp_we g4722 (.nZ(w4895), .A(w4915), .Z(w4900) );
	vdp_and g4723 (.Z(w4808), .B(w4869), .A(DCLK2) );
	vdp_and g4724 (.Z(w4805), .B(w4871), .A(DCLK2) );
	vdp_and g4725 (.Z(w4868), .B(M5), .A(w4874) );
	vdp_and g4726 (.Z(w6700), .B(w4930), .A(M5) );
	vdp_and g4727 (.Z(w6699), .B(w4876), .A(w4585) );
	vdp_and g4728 (.Z(w4914), .B(w4913), .A(HCLK1) );
	vdp_or g4729 (.Z(w4850), .B(w4847), .A(w4857) );
	vdp_or g4730 (.Z(w6701), .B(w4931), .A(w4846) );
	vdp_and g4731 (.Z(w4666), .B(w4695), .A(w4679) );
	vdp_and g4732 (.Z(w4724), .B(w4660), .A(w4722) );
	vdp_and g4733 (.Z(w6428), .B(w4722), .A(w4661) );
	vdp_and g4734 (.Z(w6429), .B(w4659), .A(w4661) );
	vdp_and g4735 (.Z(w6430), .B(w4660), .A(w4659) );
	vdp_and g4736 (.Z(w6403), .B(H40), .A(VRAMA[9]) );
	vdp_or g4737 (.Z(w4733), .B(w4662), .A(w4731) );
	vdp_or g4738 (.Z(w4732), .B(w4662), .A(w4728) );
	vdp_not g4739 (.nZ(w4659), .A(w4722) );
	vdp_oai21 g4740 (.Z(w4686), .B(w30), .A1(w31), .A2(w5) );
	vdp_oai21 g4741 (.Z(w4881), .B(w4577), .A1(w4799), .A2(w4882) );
	vdp_aoi22 g4742 (.Z(w4772), .B2(w4727), .B1(w4728), .A1(M5), .A2(w4769) );
	vdp_or3 g4743 (.Z(w4769), .B(w6624), .A(w4729), .C(w4730) );
	vdp_and3 g4744 (.Z(w4878), .B(DCLK1), .A(HCLK2), .C(w4870) );
	vdp_oai21 g4745 (.Z(w4701), .B(M5), .A1(w4679), .A2(w4700) );
	vdp_2a3oi g4746 (.Z(w4693), .B(w4684), .A1(w4683), .A2(w4), .C(SYSRES) );
	vdp_or8 g4747 (.Z(w4882), .B(w4894), .A(M5), .C(w6631), .D(w4893), .F(w4891), .E(w4892), .G(w4890), .H(w4889) );
	vdp_and9 g4748 (.Z(w4544), .B(w4852), .A(w4854), .C(w4853), .D(w4851), .F(w4849), .E(w4850), .G(w4848), .H(w4579), .I(w6701) );
	vdp_nor12 g4749 (.Z(w4799), .B(w4793), .A(1'b0), .C(w4833), .D(M5), .F(w4845), .E(w4832), .G(w4839), .H(w4831), .J(w4814), .I(w4819), .K(w4812), .L(w4825) );
	vdp_or4 g4750 (.Z(w4723), .B(w4661), .A(w4660), .C(w4721), .D(w4663) );
	vdp_nand g4751 (.Z(w4810), .B(w4809), .A(HCLK1) );
	vdp_nand g4752 (.Z(w4854), .B(w4786), .A(w6698) );
	vdp_nand g4753 (.Z(w4853), .B(w4785), .A(w6697) );
	vdp_nor g4754 (.Z(w6698), .B(w4584), .A(w4585) );
	vdp_nand3 g4755 (.Z(w4852), .B(w4785), .A(w6699), .C(w4786) );
	vdp_sr_bit g4756 (.Q(w4587), .D(w4932), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4757 (.Q(w4940), .D(w4941), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4758 (.Q(w4607), .D(w6605), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4759 (.Q(w4939), .D(w6589), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4760 (.Q(w6589), .D(w6590), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4761 (.Q(w6590), .D(w4938), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4762 (.Z(w4946), .B2(w4939), .B1(w4944), .A1(DB[4]), .A2(w4943) );
	vdp_noif0 g4763 (.A(HPOS[1]), .nZ(VRAMA[1]), .nE(w5166) );
	vdp_aon22 g4764 (.Z(w6605), .B2(w4937), .B1(w4940), .A1(M5), .A2(w4941) );
	vdp_not g4765 (.nZ(w4937), .A(M5) );
	vdp_lfsr_bit g4766 (.Q(w4947), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6622), .A1(w4946), .A2(w6621) );
	vdp_lfsr_bit g4767 (.Q(w4950), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5307), .A1(w4947), .A2(w6620) );
	vdp_lfsr_bit g4768 (.Q(w4952), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5308), .A1(w4950), .A2(w6619) );
	vdp_lfsr_bit g4769 (.Q(w4953), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5309), .A1(w4952), .A2(w6618) );
	vdp_lfsr_bit g4770 (.Q(w4957), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5310), .A1(w4953), .A2(w6617) );
	vdp_lfsr_bit g4771 (.Q(w4955), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5311), .A1(w4957), .A2(w6616) );
	vdp_lfsr_bit g4772 (.Q(w4959), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5312), .A1(w4955), .A2(w6615) );
	vdp_lfsr_bit g4773 (.Q(w4936), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5313), .A1(w4959), .A2(w6614) );
	vdp_lfsr_bit g4774 (.Q(w4963), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5026), .A1(w4936), .A2(w6613) );
	vdp_lfsr_bit g4775 (.Q(w4965), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5316), .A1(w4963), .A2(w5317) );
	vdp_lfsr_bit g4776 (.Q(w4969), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5192), .A1(w4965), .A2(w5193) );
	vdp_lfsr_bit g4777 (.Q(w4966), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5189), .A1(w4969), .A2(w5190) );
	vdp_lfsr_bit g4778 (.Q(w4968), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5187), .A1(w4966), .A2(w5188) );
	vdp_lfsr_bit g4779 (.Q(w4972), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6612), .A1(w4968), .A2(w5186) );
	vdp_lfsr_bit g4780 (.Q(w4973), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5183), .A1(w4972), .A2(w5184) );
	vdp_lfsr_bit g4781 (.Q(w4977), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6610), .A1(w4973), .A2(w6611) );
	vdp_lfsr_bit g4782 (.Q(w4976), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6609), .A1(w4977), .A2(w6608) );
	vdp_lfsr_bit g4783 (.Q(w4981), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5180), .A1(w4976), .A2(w5181) );
	vdp_lfsr_bit g4784 (.Q(w4983), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5179), .A1(w4981), .A2(w5178) );
	vdp_lfsr_bit g4785 (.Q(w4935), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5176), .A1(w4983), .A2(w5177) );
	vdp_bufif0 g4786 (.A(w4936), .Z(VRAMA[1]), .nE(w6607) );
	vdp_bufif0 g4787 (.A(1'b0), .Z(VRAMA[1]), .nE(w5200) );
	vdp_noif0 g4788 (.A(w4935), .nZ(DB[4]), .nE(w5318) );
	vdp_sr_bit g4789 (.Q(w4991), .D(w6592), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4790 (.Q(w6592), .D(w6591), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4791 (.Q(w6591), .D(w6410), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4792 (.Z(w4945), .B2(w4991), .B1(w4944), .A1(DB[5]), .A2(w4943) );
	vdp_noif0 g4793 (.A(w5000), .nZ(VRAMA[2]), .nE(w5166) );
	vdp_lfsr_bit g4794 (.Q(w4948), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6622), .A1(w4945), .A2(w6621) );
	vdp_lfsr_bit g4795 (.Q(w4949), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5307), .A1(w4948), .A2(w6620) );
	vdp_lfsr_bit g4796 (.Q(w4951), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5308), .A1(w4949), .A2(w6619) );
	vdp_lfsr_bit g4797 (.Q(w4954), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5309), .A1(w4951), .A2(w6618) );
	vdp_lfsr_bit g4798 (.Q(w4958), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5310), .A1(w4954), .A2(w6617) );
	vdp_lfsr_bit g4799 (.Q(w4956), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5311), .A1(w4958), .A2(w6616) );
	vdp_lfsr_bit g4800 (.Q(w4960), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5312), .A1(w4956), .A2(w6615) );
	vdp_lfsr_bit g4801 (.Q(w4961), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5313), .A1(w4960), .A2(w6614) );
	vdp_lfsr_bit g4802 (.Q(w4964), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5026), .A1(w4961), .A2(w6613) );
	vdp_lfsr_bit g4803 (.Q(w4962), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5316), .A1(w4964), .A2(w5317) );
	vdp_lfsr_bit g4804 (.Q(w4970), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5192), .A1(w4962), .A2(w5193) );
	vdp_lfsr_bit g4805 (.Q(w4967), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5189), .A1(w4970), .A2(w5190) );
	vdp_lfsr_bit g4806 (.Q(w4971), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5187), .A1(w4967), .A2(w5188) );
	vdp_lfsr_bit g4807 (.Q(w4975), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6612), .A1(w4971), .A2(w5186) );
	vdp_lfsr_bit g4808 (.Q(w4974), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5183), .A1(w4975), .A2(w5184) );
	vdp_lfsr_bit g4809 (.Q(w4978), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6610), .A1(w4974), .A2(w6611) );
	vdp_lfsr_bit g4810 (.Q(w4979), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6609), .A1(w4978), .A2(w6608) );
	vdp_lfsr_bit g4811 (.Q(w4980), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5180), .A1(w4979), .A2(w5181) );
	vdp_lfsr_bit g4812 (.Q(w4984), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5179), .A1(w4980), .A2(w5178) );
	vdp_lfsr_bit g4813 (.Q(w4988), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5176), .A1(w4984), .A2(w5177) );
	vdp_bufif0 g4814 (.A(w4961), .Z(VRAMA[2]), .nE(w6607) );
	vdp_bufif0 g4815 (.A(1'b1), .Z(VRAMA[2]), .nE(w5200) );
	vdp_noif0 g4816 (.A(w4988), .nZ(DB[5]), .nE(w5318) );
	vdp_aon22 g4817 (.Z(w4987), .B2(w4977), .B1(w5050), .A1(w4989), .A2(w4935) );
	vdp_dlatch_inv g4818 (.nQ(w5001), .D(w4994), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g4819 (.nQ(w4996), .D(w4942), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g4820 (.Z(w4995), .B(w4996), .A(DCLK2) );
	vdp_nand g4821 (.Z(w4994), .B(HCLK1), .A(w4607) );
	vdp_nand g4822 (.Z(w4942), .B(HCLK1), .A(w4941) );
	vdp_sr_bit g4823 (.Q(w4993), .D(w6594), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4824 (.Q(w6594), .D(w6593), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4825 (.Q(w6593), .D(w4998), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4826 (.Z(w5009), .B2(w4993), .B1(w4944), .A1(DB[6]), .A2(w4992) );
	vdp_noif0 g4827 (.A(w5007), .nZ(w6411), .nE(w5166) );
	vdp_lfsr_bit g4828 (.Q(w5011), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6622), .A1(w5009), .A2(w6621) );
	vdp_lfsr_bit g4829 (.Q(w5012), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5307), .A1(w5011), .A2(w6620) );
	vdp_lfsr_bit g4830 (.Q(w5015), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5308), .A1(w5012), .A2(w6619) );
	vdp_lfsr_bit g4831 (.Q(w5016), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5309), .A1(w5015), .A2(w6618) );
	vdp_lfsr_bit g4832 (.Q(w5021), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5310), .A1(w5016), .A2(w6617) );
	vdp_lfsr_bit g4833 (.Q(w5020), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5311), .A1(w5021), .A2(w6616) );
	vdp_lfsr_bit g4834 (.Q(w5023), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5312), .A1(w5020), .A2(w6615) );
	vdp_lfsr_bit g4835 (.Q(w5025), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5313), .A1(w5023), .A2(w6614) );
	vdp_lfsr_bit g4836 (.Q(w5028), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5026), .A1(w5025), .A2(w6613) );
	vdp_lfsr_bit g4837 (.Q(w5030), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5316), .A1(w5028), .A2(w5317) );
	vdp_lfsr_bit g4838 (.Q(w5032), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5192), .A1(w5030), .A2(w5193) );
	vdp_lfsr_bit g4839 (.Q(w5034), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5189), .A1(w5032), .A2(w5190) );
	vdp_lfsr_bit g4840 (.Q(w5036), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5187), .A1(w5034), .A2(w5188) );
	vdp_lfsr_bit g4841 (.Q(w5039), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6612), .A1(w5036), .A2(w5186) );
	vdp_lfsr_bit g4842 (.Q(w5040), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5183), .A1(w5039), .A2(w5184) );
	vdp_lfsr_bit g4843 (.Q(w5041), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6610), .A1(w5040), .A2(w6611) );
	vdp_lfsr_bit g4844 (.Q(w5046), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6609), .A1(w5041), .A2(w6608) );
	vdp_lfsr_bit g4845 (.Q(w5045), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5180), .A1(w5046), .A2(w5181) );
	vdp_lfsr_bit g4846 (.Q(w5048), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5179), .A1(w5045), .A2(w5178) );
	vdp_lfsr_bit g4847 (.Q(w4990), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5176), .A1(w5048), .A2(w5177) );
	vdp_bufif0 g4848 (.A(w5025), .Z(w6411), .nE(w6607) );
	vdp_bufif0 g4849 (.A(w4987), .Z(w6411), .nE(w5200) );
	vdp_noif0 g4850 (.A(w4990), .nZ(DB[6]), .nE(w5318) );
	vdp_aon22 g4851 (.Z(w5049), .B2(w4978), .B1(w5050), .A1(w4989), .A2(w4988) );
	vdp_sr_bit g4852 (.Q(w5003), .D(w5001), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g4853 (.Q(w4997), .D(w4996), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_and g4854 (.Z(w4999), .B(w5001), .A(DCLK2) );
	vdp_and g4855 (.Z(w5005), .B(DCLK2), .A(w5003) );
	vdp_and g4856 (.Z(w5002), .B(w4997), .A(DCLK2) );
	vdp_sr_bit g4857 (.Q(w5063), .D(w6595), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4858 (.Q(w6595), .D(w6596), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4859 (.Q(w6596), .D(w5004), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4860 (.Z(w5008), .B2(w5063), .B1(w4944), .A1(w160), .A2(w4992) );
	vdp_noif0 g4861 (.A(w5061), .nZ(VRAMA[4]), .nE(w5166) );
	vdp_lfsr_bit g4862 (.Q(w5010), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6622), .A1(w5008), .A2(w6621) );
	vdp_lfsr_bit g4863 (.Q(w5013), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5307), .A1(w5010), .A2(w6620) );
	vdp_lfsr_bit g4864 (.Q(w5014), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5308), .A1(w5013), .A2(w6619) );
	vdp_lfsr_bit g4865 (.Q(w5017), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5309), .A1(w5014), .A2(w6618) );
	vdp_lfsr_bit g4866 (.Q(w5018), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5310), .A1(w5017), .A2(w6617) );
	vdp_lfsr_bit g4867 (.Q(w5019), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5311), .A1(w5018), .A2(w6616) );
	vdp_lfsr_bit g4868 (.Q(w5022), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5312), .A1(w5019), .A2(w6615) );
	vdp_lfsr_bit g4869 (.Q(w5024), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5313), .A1(w5022), .A2(w6614) );
	vdp_lfsr_bit g4870 (.Q(w5027), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5026), .A1(w5024), .A2(w6613) );
	vdp_lfsr_bit g4871 (.Q(w5029), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5316), .A1(w5027), .A2(w5317) );
	vdp_lfsr_bit g4872 (.Q(w5031), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5192), .A1(w5029), .A2(w5193) );
	vdp_lfsr_bit g4873 (.Q(w5033), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5189), .A1(w5031), .A2(w5190) );
	vdp_lfsr_bit g4874 (.Q(w5035), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5187), .A1(w5033), .A2(w5188) );
	vdp_lfsr_bit g4875 (.Q(w5038), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6612), .A1(w5035), .A2(w5186) );
	vdp_lfsr_bit g4876 (.Q(w5037), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5183), .A1(w5038), .A2(w5184) );
	vdp_lfsr_bit g4877 (.Q(w5042), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6610), .A1(w5037), .A2(w6611) );
	vdp_lfsr_bit g4878 (.Q(w5043), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6609), .A1(w5042), .A2(w6608) );
	vdp_lfsr_bit g4879 (.Q(w5044), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5180), .A1(w5043), .A2(w5181) );
	vdp_lfsr_bit g4880 (.Q(w5047), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5179), .A1(w5044), .A2(w5178) );
	vdp_lfsr_bit g4881 (.Q(w5065), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5176), .A1(w5047), .A2(w5177) );
	vdp_bufif0 g4882 (.A(w5024), .Z(VRAMA[4]), .nE(w6607) );
	vdp_bufif0 g4883 (.A(w5049), .Z(VRAMA[4]), .nE(w5200) );
	vdp_noif0 g4884 (.A(w5065), .nZ(w160), .nE(w5318) );
	vdp_aon22 g4885 (.Z(w5066), .B2(w5041), .B1(w5050), .A1(w4989), .A2(w4990) );
	vdp_aon22 g4886 (.Z(w5060), .B2(w5053), .B1(w132), .A1(w5006), .A2(w5059) );
	vdp_not g4887 (.nZ(w5006), .A(w132) );
	vdp_comp_str g4888 (.nZ(w5054), .A(w5002), .Z(w5055) );
	vdp_comp_str g4889 (.nZ(w5058), .A(w5005), .Z(w5057) );
	vdp_sr_bit g4890 (.Q(w5062), .D(w6598), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4891 (.Q(w6598), .D(w6597), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4892 (.Q(w6597), .D(w5056), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4893 (.Z(w5107), .B2(w5062), .B1(w4944), .A1(DB[8]), .A2(w4992) );
	vdp_noif0 g4894 (.A(w5060), .nZ(VRAMA[5]), .nE(w5166) );
	vdp_lfsr_bit g4895 (.Q(w5105), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6622), .A1(w5107), .A2(w6621) );
	vdp_lfsr_bit g4896 (.Q(w5102), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5307), .A1(w5105), .A2(w6620) );
	vdp_lfsr_bit g4897 (.Q(w5101), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5308), .A1(w5102), .A2(w6619) );
	vdp_lfsr_bit g4898 (.Q(w5098), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5309), .A1(w5101), .A2(w6618) );
	vdp_lfsr_bit g4899 (.Q(w5097), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5310), .A1(w5098), .A2(w6617) );
	vdp_lfsr_bit g4900 (.Q(w5094), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5311), .A1(w5097), .A2(w6616) );
	vdp_lfsr_bit g4901 (.Q(w5093), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5312), .A1(w5094), .A2(w6615) );
	vdp_lfsr_bit g4902 (.Q(w5071), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5313), .A1(w5093), .A2(w6614) );
	vdp_lfsr_bit g4903 (.Q(w5090), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5026), .A1(w5071), .A2(w6613) );
	vdp_lfsr_bit g4904 (.Q(w5064), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5316), .A1(w5090), .A2(w5317) );
	vdp_lfsr_bit g4905 (.Q(w5087), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5192), .A1(w5064), .A2(w5193) );
	vdp_lfsr_bit g4906 (.Q(w5086), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5189), .A1(w5087), .A2(w5190) );
	vdp_lfsr_bit g4907 (.Q(w5083), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5187), .A1(w5086), .A2(w5188) );
	vdp_lfsr_bit g4908 (.Q(w5081), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6612), .A1(w5083), .A2(w5186) );
	vdp_lfsr_bit g4909 (.Q(w5080), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5183), .A1(w5081), .A2(w5184) );
	vdp_lfsr_bit g4910 (.Q(w5069), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6610), .A1(w5080), .A2(w6611) );
	vdp_lfsr_bit g4911 (.Q(w5076), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6609), .A1(w5069), .A2(w6608) );
	vdp_lfsr_bit g4912 (.Q(w5074), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5180), .A1(w5076), .A2(w5181) );
	vdp_lfsr_bit g4913 (.Q(w5072), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5179), .A1(w5074), .A2(w5178) );
	vdp_lfsr_bit g4914 (.Q(w5089), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5176), .A1(w5072), .A2(w5177) );
	vdp_bufif0 g4915 (.A(w5071), .Z(VRAMA[5]), .nE(w6607) );
	vdp_bufif0 g4916 (.A(w5066), .Z(VRAMA[5]), .nE(w5200) );
	vdp_noif0 g4917 (.A(w5089), .nZ(DB[8]), .nE(w5318) );
	vdp_aon22 g4918 (.Z(w5068), .B2(w5042), .B1(w5050), .A1(w4989), .A2(w5065) );
	vdp_slatch g4919 (.D(S[0]), .nC(w5058), .C(w5057), .Q(w5112) );
	vdp_slatch g4920 (.D(S[0]), .nC(w5054), .C(w5055), .Q(w5052) );
	vdp_aoi22 g4921 (.Z(w5059), .B2(w5111), .B1(w5112), .A1(w5110), .A2(w5052) );
	vdp_sr_bit g4922 (.Q(w5120), .D(w6600), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4923 (.Q(w6600), .D(w6599), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4924 (.Q(w6599), .D(w5108), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4925 (.Z(w5106), .B2(w5120), .B1(w4944), .A1(DB[9]), .A2(w4992) );
	vdp_noif0 g4926 (.A(w5109), .nZ(VRAMA[6]), .nE(w5166) );
	vdp_lfsr_bit g4927 (.Q(w5104), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6622), .A1(w5106), .A2(w6621) );
	vdp_lfsr_bit g4928 (.Q(w5103), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w5307), .A1(w5104), .A2(w6620) );
	vdp_lfsr_bit g4929 (.Q(w5100), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w5308), .A1(w5103), .A2(w6619) );
	vdp_lfsr_bit g4930 (.Q(w5099), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w5309), .A1(w5100), .A2(w6618) );
	vdp_lfsr_bit g4931 (.Q(w5096), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w5310), .A1(w5099), .A2(w6617) );
	vdp_lfsr_bit g4932 (.Q(w5095), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w5311), .A1(w5096), .A2(w6616) );
	vdp_lfsr_bit g4933 (.Q(w5092), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w5312), .A1(w5095), .A2(w6615) );
	vdp_lfsr_bit g4934 (.Q(w5070), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w5313), .A1(w5092), .A2(w6614) );
	vdp_lfsr_bit g4935 (.Q(w5091), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5026), .A1(w5070), .A2(w6613) );
	vdp_lfsr_bit g4936 (.Q(w5118), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5316), .A1(w5091), .A2(w5317) );
	vdp_lfsr_bit g4937 (.Q(w5088), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5192), .A1(w5118), .A2(w5193) );
	vdp_lfsr_bit g4938 (.Q(w5085), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5189), .A1(w5088), .A2(w5190) );
	vdp_lfsr_bit g4939 (.Q(w5084), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5187), .A1(w5085), .A2(w5188) );
	vdp_lfsr_bit g4940 (.Q(w5082), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6612), .A1(w5084), .A2(w5186) );
	vdp_lfsr_bit g4941 (.Q(w5079), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5183), .A1(w5082), .A2(w5184) );
	vdp_lfsr_bit g4942 (.Q(w5078), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6610), .A1(w5079), .A2(w6611) );
	vdp_lfsr_bit g4943 (.Q(w5077), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6609), .A1(w5078), .A2(w6608) );
	vdp_lfsr_bit g4944 (.Q(w5075), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5180), .A1(w5077), .A2(w5181) );
	vdp_lfsr_bit g4945 (.Q(w5073), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5179), .A1(w5075), .A2(w5178) );
	vdp_lfsr_bit g4946 (.Q(w5115), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5176), .A1(w5073), .A2(w5177) );
	vdp_bufif0 g4947 (.A(w5070), .Z(VRAMA[6]), .nE(w6607) );
	vdp_bufif0 g4948 (.A(w5068), .Z(VRAMA[6]), .nE(w5200) );
	vdp_noif0 g4949 (.A(w5115), .nZ(DB[9]), .nE(w5318) );
	vdp_aon22 g4950 (.Z(w5117), .B2(w5069), .B1(w5050), .A1(w4989), .A2(w5089) );
	vdp_aoi22 g4951 (.Z(w5109), .B2(w5111), .B1(w5122), .A1(w5110), .A2(w5113) );
	vdp_slatch g4952 (.D(S[1]), .nC(w5058), .C(w5057), .Q(w5122) );
	vdp_slatch g4953 (.D(S[1]), .nC(w5054), .C(w5055), .Q(w5113) );
	vdp_sr_bit g4954 (.Q(w5119), .D(w6602), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4955 (.Q(w6602), .D(w6601), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4956 (.Q(w6601), .D(w5123), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4957 (.Z(w5165), .B2(w5119), .B1(w4944), .A1(DB[10]), .A2(w4992) );
	vdp_noif0 g4958 (.A(w5168), .nZ(VRAMA[7]), .nE(w5169) );
	vdp_lfsr_bit g4959 (.Q(w5164), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6622), .A1(w5165), .A2(w6621) );
	vdp_lfsr_bit g4960 (.Q(w5159), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5307), .A1(w5164), .A2(w6620) );
	vdp_lfsr_bit g4961 (.Q(w5160), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5308), .A1(w5159), .A2(w6619) );
	vdp_lfsr_bit g4962 (.Q(w5154), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5309), .A1(w5160), .A2(w6618) );
	vdp_lfsr_bit g4963 (.Q(w5155), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5310), .A1(w5154), .A2(w6617) );
	vdp_lfsr_bit g4964 (.Q(w5152), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5311), .A1(w5155), .A2(w6616) );
	vdp_lfsr_bit g4965 (.Q(w5150), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5312), .A1(w5152), .A2(w6615) );
	vdp_lfsr_bit g4966 (.Q(w5116), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5313), .A1(w5150), .A2(w6614) );
	vdp_lfsr_bit g4967 (.Q(w5147), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5026), .A1(w5116), .A2(w6613) );
	vdp_lfsr_bit g4968 (.Q(w5143), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5316), .A1(w5147), .A2(w5317) );
	vdp_lfsr_bit g4969 (.Q(w5145), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5192), .A1(w5143), .A2(w5193) );
	vdp_lfsr_bit g4970 (.Q(w5142), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5189), .A1(w5145), .A2(w5190) );
	vdp_lfsr_bit g4971 (.Q(w5141), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5187), .A1(w5142), .A2(w5188) );
	vdp_lfsr_bit g4972 (.Q(w5138), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6612), .A1(w5141), .A2(w5186) );
	vdp_lfsr_bit g4973 (.Q(w5136), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5183), .A1(w5138), .A2(w5184) );
	vdp_lfsr_bit g4974 (.Q(w5134), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6610), .A1(w5136), .A2(w6611) );
	vdp_lfsr_bit g4975 (.Q(w5132), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6609), .A1(w5134), .A2(w6608) );
	vdp_lfsr_bit g4976 (.Q(w5130), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5180), .A1(w5132), .A2(w5181) );
	vdp_lfsr_bit g4977 (.Q(w5128), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5179), .A1(w5130), .A2(w5178) );
	vdp_lfsr_bit g4978 (.Q(w5126), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5176), .A1(w5128), .A2(w5177) );
	vdp_bufif0 g4979 (.A(w5116), .Z(VRAMA[7]), .nE(w6607) );
	vdp_bufif0 g4980 (.A(w5117), .Z(VRAMA[7]), .nE(w5200) );
	vdp_noif0 g4981 (.A(w5126), .nZ(DB[10]), .nE(w5318) );
	vdp_aon22 g4982 (.Z(w5125), .B2(w5078), .B1(w5050), .A1(w4989), .A2(w5115) );
	vdp_aoi22 g4983 (.Z(w5168), .B2(w5111), .B1(w5170), .A1(w5110), .A2(w5121) );
	vdp_slatch g4984 (.D(S[2]), .nC(w5058), .C(w5057), .Q(w5170) );
	vdp_slatch g4985 (.D(S[2]), .nC(w5054), .C(w5055), .Q(w5121) );
	vdp_sr_bit g4986 (.Q(w5195), .D(w29), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4987 (.Q(w5194), .D(w22), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4988 (.Z(w5162), .B2(w4582), .B1(w4944), .A1(w170), .A2(w4992) );
	vdp_noif0 g4989 (.A(w5167), .nZ(VRAMA[8]), .nE(w5169) );
	vdp_lfsr_bit g4990 (.Q(w5163), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6622), .A1(w5162), .A2(w6621) );
	vdp_lfsr_bit g4991 (.Q(w5158), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5307), .A1(w5163), .A2(w6620) );
	vdp_lfsr_bit g4992 (.Q(w5161), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5308), .A1(w5158), .A2(w6619) );
	vdp_lfsr_bit g4993 (.Q(w5157), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5309), .A1(w5161), .A2(w6618) );
	vdp_lfsr_bit g4994 (.Q(w5156), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5310), .A1(w5157), .A2(w6617) );
	vdp_lfsr_bit g4995 (.Q(w5153), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5311), .A1(w5156), .A2(w6616) );
	vdp_lfsr_bit g4996 (.Q(w5151), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5312), .A1(w5153), .A2(w6615) );
	vdp_lfsr_bit g4997 (.Q(w5149), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5313), .A1(w5151), .A2(w6614) );
	vdp_lfsr_bit g4998 (.Q(w5148), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5026), .A1(w5149), .A2(w6613) );
	vdp_lfsr_bit g4999 (.Q(w5146), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5316), .A1(w5148), .A2(w5317) );
	vdp_lfsr_bit g5000 (.Q(w5144), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5192), .A1(w5146), .A2(w5193) );
	vdp_lfsr_bit g5001 (.Q(w5140), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5189), .A1(w5144), .A2(w5190) );
	vdp_lfsr_bit g5002 (.Q(w5139), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5187), .A1(w5140), .A2(w5188) );
	vdp_lfsr_bit g5003 (.Q(w5137), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6612), .A1(w5139), .A2(w5186) );
	vdp_lfsr_bit g5004 (.Q(w5135), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5183), .A1(w5137), .A2(w5184) );
	vdp_lfsr_bit g5005 (.Q(w5133), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6610), .A1(w5135), .A2(w6611) );
	vdp_lfsr_bit g5006 (.Q(w5131), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6609), .A1(w5133), .A2(w6608) );
	vdp_lfsr_bit g5007 (.Q(w5129), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5180), .A1(w5131), .A2(w5181) );
	vdp_lfsr_bit g5008 (.Q(w5127), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5179), .A1(w5129), .A2(w5178) );
	vdp_lfsr_bit g5009 (.Q(w5191), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5176), .A1(w5127), .A2(w5177) );
	vdp_bufif0 g5010 (.A(1'b0), .Z(VRAMA[0]), .nE(w6607) );
	vdp_bufif0 g5011 (.A(w5125), .Z(VRAMA[8]), .nE(w5200) );
	vdp_noif0 g5012 (.A(w5191), .nZ(w170), .nE(w5318) );
	vdp_aon22 g5013 (.Z(w5201), .B2(w5174), .B1(w5050), .A1(w4989), .A2(w5126) );
	vdp_aoi22 g5014 (.Z(w5167), .B2(w5111), .B1(w5171), .A1(w5110), .A2(w5172) );
	vdp_slatch g5015 (.D(S[3]), .nC(w5058), .C(w5057), .Q(w5171) );
	vdp_slatch g5016 (.D(S[3]), .nC(w5054), .C(w5055), .Q(w5172) );
	vdp_bufif0 g5017 (.A(1'b0), .Z(VRAMA[0]), .nE(w5200) );
	vdp_bufif0 g5018 (.A(w5204), .Z(VRAMA[8]), .nE(w5208) );
	vdp_aon22 g5019 (.Z(w5231), .B2(w4592), .B1(w4944), .A1(w156), .A2(w4992) );
	vdp_lfsr_bit g5020 (.Q(w5229), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6622), .A1(w5231), .A2(w6621) );
	vdp_lfsr_bit g5021 (.Q(w5227), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5307), .A1(w5229), .A2(w6620) );
	vdp_lfsr_bit g5022 (.Q(w5225), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5308), .A1(w5227), .A2(w6619) );
	vdp_lfsr_bit g5023 (.Q(w5223), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5309), .A1(w5225), .A2(w6618) );
	vdp_lfsr_bit g5024 (.Q(w5220), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5310), .A1(w5223), .A2(w6617) );
	vdp_lfsr_bit g5025 (.Q(w5219), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5311), .A1(w5220), .A2(w6616) );
	vdp_lfsr_bit g5026 (.Q(w5217), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5312), .A1(w5219), .A2(w6615) );
	vdp_lfsr_bit g5027 (.Q(w5215), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5313), .A1(w5217), .A2(w6614) );
	vdp_lfsr_bit g5028 (.Q(w5199), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5026), .A1(w5215), .A2(w6613) );
	vdp_lfsr_bit g5029 (.Q(w5197), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5316), .A1(w5199), .A2(w5317) );
	vdp_noif0 g5030 (.A(w5197), .nZ(w156), .nE(w5318) );
	vdp_not g5031 (.nZ(w5185), .A(M5) );
	vdp_not g5032 (.nZ(w5196), .A(H40) );
	vdp_noif0 g5033 (.A(1'b1), .nZ(VRAMA[0]), .nE(w5166) );
	vdp_aoi22 g5034 (.Z(w5053), .B2(w5236), .B1(w5199), .A1(w5110), .A2(w5197) );
	vdp_not g5035 (.nZ(w5233), .A(M5) );
	vdp_or g5036 (.Z(w5234), .B(w5195), .A(w5194) );
	vdp_sr_bit g5037 (.Q(w5205), .D(w9), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5038 (.Q(w5211), .D(w30), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_comp_we g5039 (.nZ(w5176), .A(w5203), .Z(w5177) );
	vdp_comp_we g5040 (.nZ(w5179), .A(w5203), .Z(w5178) );
	vdp_comp_we g5041 (.nZ(w5180), .A(w5203), .Z(w5181) );
	vdp_comp_we g5042 (.nZ(w6609), .A(w5203), .Z(w6608) );
	vdp_comp_we g5043 (.nZ(w6610), .A(w5203), .Z(w6611) );
	vdp_comp_we g5044 (.nZ(w5050), .A(H40), .Z(w4989) );
	vdp_comp_we g5045 (.nZ(w5183), .A(w5203), .Z(w5184) );
	vdp_comp_we g5046 (.nZ(w6612), .A(w5203), .Z(w5186) );
	vdp_comp_we g5047 (.nZ(w5187), .A(w5203), .Z(w5188) );
	vdp_comp_we g5048 (.nZ(w5189), .A(w5203), .Z(w5190) );
	vdp_comp_we g5049 (.nZ(w5192), .A(w5203), .Z(w5193) );
	vdp_comp_we g5050 (.nZ(w5111), .A(w5194), .Z(w5110) );
	vdp_not g5051 (.nZ(w5169), .A(w5198) );
	vdp_not g5052 (.nZ(w5166), .A(w5198) );
	vdp_not g5053 (.nZ(w5200), .A(w5207) );
	vdp_not g5054 (.nZ(w6607), .A(w5182) );
	vdp_and g5055 (.Z(w5182), .B(w5205), .A(w5185) );
	vdp_oai21 g5056 (.Z(w5210), .B(w5185), .A1(w5211), .A2(w5205) );
	vdp_aon333 g5057 (.Z(w4543), .B1(M5), .A1(1'b1), .C1(M5), .A2(w5185), .A3(w5149), .B2(w5133), .B3(w5196), .C2(H40), .C3(w5191) );
	vdp_aon22 g5058 (.Z(w5230), .B2(w4598), .B1(w4944), .A1(DB[2]), .A2(w4992) );
	vdp_lfsr_bit g5059 (.Q(w5228), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6622), .A1(w5230), .A2(w6621) );
	vdp_lfsr_bit g5060 (.Q(w5226), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5307), .A1(w5228), .A2(w6620) );
	vdp_lfsr_bit g5061 (.Q(w5224), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5308), .A1(w5226), .A2(w6619) );
	vdp_lfsr_bit g5062 (.Q(w5222), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5309), .A1(w5224), .A2(w6618) );
	vdp_lfsr_bit g5063 (.Q(w5221), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5310), .A1(w5222), .A2(w6617) );
	vdp_lfsr_bit g5064 (.Q(w5218), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5311), .A1(w5221), .A2(w6616) );
	vdp_lfsr_bit g5065 (.Q(w5216), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5312), .A1(w5218), .A2(w6615) );
	vdp_lfsr_bit g5066 (.Q(w5214), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5313), .A1(w5216), .A2(w6614) );
	vdp_lfsr_bit g5067 (.Q(w5213), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5026), .A1(w5214), .A2(w6613) );
	vdp_lfsr_bit g5068 (.Q(w5212), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5316), .A1(w5213), .A2(w5317) );
	vdp_noif0 g5069 (.A(w5212), .nZ(DB[2]), .nE(w5318) );
	vdp_aoi22 g5070 (.Z(w5061), .B2(w5236), .B1(w5213), .A1(w5110), .A2(w5212) );
	vdp_aoi22 g5071 (.Z(w5249), .B2(w5236), .B1(w5250), .A1(w5110), .A2(w4545) );
	vdp_noif0 g5072 (.A(w5249), .nZ(VRAMA[9]), .nE(w5169) );
	vdp_slatch g5074 (.D(S[4]), .nC(w5055), .C(w5054), .Q(w4545) );
	vdp_and g5075 (.Z(w5198), .B(w5233), .A(w5234) );
	vdp_slatch g5076 (.D(w612), .nC(w5315), .C(w5314), .Q(w5174) );
	vdp_slatch g5077 (.D(w617), .nC(w5315), .C(w5314), .Q(w5206) );
	vdp_bufif0 g5078 (.A(w5201), .Z(VRAMA[9]), .nE(w5239) );
	vdp_bufif0 g5079 (.A(w5206), .Z(VRAMA[16]), .nE(w5239) );
	vdp_and g5080 (.Z(w5207), .B(w5205), .A(M5) );
	vdp_not g5081 (.nZ(w5239), .A(w5207) );
	vdp_not g5082 (.nZ(w5208), .A(w5209) );
	vdp_not g5083 (.nZ(w5209), .A(w5210) );
	vdp_xor g5084 (.Z(w5238), .B(w5206), .A(VRAMA[16]) );
	vdp_xor g5085 (.Z(w5242), .B(w5244), .A(w5243) );
	vdp_and3 g5086 (.Z(w5235), .B(w5248), .A(w5245), .C(M5) );
	vdp_nor g5087 (.Z(w5244), .B(H40), .A(w5174) );
	vdp_nor g5088 (.Z(w5243), .B(H40), .A(VRAMA[9]) );
	vdp_aon22 g5089 (.Z(w5269), .B2(w4589), .B1(w4944), .A1(DB[1]), .A2(w4992) );
	vdp_lfsr_bit g5090 (.Q(w5268), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6622), .A1(w5269), .A2(w6621) );
	vdp_lfsr_bit g5091 (.Q(w5267), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5307), .A1(w5268), .A2(w6620) );
	vdp_lfsr_bit g5092 (.Q(w5266), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5308), .A1(w5267), .A2(w6619) );
	vdp_lfsr_bit g5093 (.Q(w5265), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5309), .A1(w5266), .A2(w6618) );
	vdp_lfsr_bit g5094 (.Q(w5264), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5310), .A1(w5265), .A2(w6617) );
	vdp_lfsr_bit g5095 (.Q(w5263), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5311), .A1(w5264), .A2(w6616) );
	vdp_lfsr_bit g5096 (.Q(w5262), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5312), .A1(w5263), .A2(w6615) );
	vdp_lfsr_bit g5097 (.Q(w5261), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5313), .A1(w5262), .A2(w6614) );
	vdp_lfsr_bit g5098 (.Q(w5247), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5026), .A1(w5261), .A2(w6613) );
	vdp_lfsr_bit g5099 (.Q(w5259), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5316), .A1(w5247), .A2(w5317) );
	vdp_noif0 g5100 (.A(w5259), .nZ(DB[1]), .nE(w5318) );
	vdp_slatch g5101 (.D(w685), .nC(w5315), .C(w5314), .Q(w5204) );
	vdp_slatch g5102 (.D(w661), .nC(w5315), .C(w5314), .Q(w5258) );
	vdp_xor g5103 (.Z(w5241), .B(w5258), .A(VRAMA[15]) );
	vdp_xor g5104 (.Z(w5240), .B(w5204), .A(VRAMA[10]) );
	vdp_aon22 g5105 (.Z(w5278), .B2(w4588), .B1(w4944), .A1(DB[0]), .A2(w4992) );
	vdp_lfsr_bit g5106 (.Q(w5279), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6622), .A1(w5278), .A2(w6621) );
	vdp_lfsr_bit g5107 (.Q(w5280), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5307), .A1(w5279), .A2(w6620) );
	vdp_lfsr_bit g5108 (.Q(w5281), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5308), .A1(w5280), .A2(w6619) );
	vdp_lfsr_bit g5109 (.Q(w5283), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5309), .A1(w5281), .A2(w6618) );
	vdp_lfsr_bit g5110 (.Q(w5282), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5310), .A1(w5283), .A2(w6617) );
	vdp_lfsr_bit g5111 (.Q(w5285), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5311), .A1(w5282), .A2(w6616) );
	vdp_lfsr_bit g5112 (.Q(w5284), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5312), .A1(w5285), .A2(w6615) );
	vdp_lfsr_bit g5113 (.Q(w5286), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5313), .A1(w5284), .A2(w6614) );
	vdp_lfsr_bit g5114 (.Q(w5260), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5026), .A1(w5286), .A2(w6613) );
	vdp_lfsr_bit g5115 (.Q(w6606), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5316), .A1(w5260), .A2(w5317) );
	vdp_noif0 g5116 (.A(w6606), .nZ(DB[0]), .nE(w5318) );
	vdp_slatch g5117 (.D(w698), .nC(w5315), .C(w5314), .Q(w5257) );
	vdp_slatch g5118 (.D(w681), .nC(w5315), .C(w5314), .Q(w5301) );
	vdp_xor g5119 (.Z(w5254), .B(w5301), .A(VRAMA[14]) );
	vdp_xor g5120 (.Z(w5253), .B(w5257), .A(VRAMA[11]) );
	vdp_slatch g5121 (.D(S[5]), .nC(w5057), .C(w5058), .Q(w5272) );
	vdp_slatch g5122 (.D(S[5]), .nC(w5055), .C(w5054), .Q(w5251) );
	vdp_slatch g5123 (.D(S[6]), .nC(w5057), .C(w5058), .Q(w5273) );
	vdp_slatch g5124 (.D(S[6]), .nC(w5055), .C(w5054), .Q(w5271) );
	vdp_slatch g5125 (.D(S[7]), .nC(w5057), .C(w5058), .Q(w5306) );
	vdp_slatch g5126 (.D(S[7]), .nC(w5055), .C(w5054), .Q(w5236) );
	vdp_slatch g5127 (.D(w698), .nC(w5276), .C(w5277), .Q(w5274) );
	vdp_slatch g5128 (.D(w681), .nC(w5276), .C(w5277), .Q(w5270) );
	vdp_bufif0 g5129 (.A(w5257), .Z(VRAMA[9]), .nE(w5208) );
	vdp_bufif0 g5130 (.A(w5204), .Z(VRAMA[10]), .nE(w5239) );
	vdp_bufif0 g5131 (.A(w5295), .Z(VRAMA[10]), .nE(w5208) );
	vdp_bufif0 g5132 (.A(w5258), .Z(VRAMA[13]), .nE(w5208) );
	vdp_bufif0 g5133 (.A(w5301), .Z(VRAMA[14]), .nE(w5239) );
	vdp_bufif0 g5134 (.A(w5257), .Z(VRAMA[11]), .nE(w5239) );
	vdp_bufif0 g5135 (.A(w5294), .Z(VRAMA[13]), .nE(w5239) );
	vdp_bufif0 g5136 (.A(w5295), .Z(VRAMA[12]), .nE(w5239) );
	vdp_bufif0 g5137 (.A(w5294), .Z(VRAMA[11]), .nE(w5208) );
	vdp_bufif0 g5138 (.A(w5301), .Z(VRAMA[12]), .nE(w5208) );
	vdp_bufif0 g5139 (.A(w5258), .Z(VRAMA[15]), .nE(w5239) );
	vdp_slatch g5140 (.D(w719), .nC(w5315), .C(w5314), .Q(w5295) );
	vdp_slatch g5141 (.D(w725), .nC(w5315), .C(w5314), .Q(w5294) );
	vdp_xor g5142 (.Z(w5256), .B(w5294), .A(VRAMA[13]) );
	vdp_xor g5143 (.Z(w5255), .B(w5295), .A(VRAMA[12]) );
	vdp_dlatch_inv g5144 (.nQ(w5293), .D(w5298), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5145 (.nQ(w5292), .D(w5299), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5146 (.nQ(w5291), .D(w6728), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5147 (.nQ(w5290), .D(w6730), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5148 (.nQ(w5289), .D(w5300), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5149 (.nQ(w5288), .D(w5297), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5150 (.nQ(w5287), .D(w6729), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5151 (.nQ(w6404), .D(w5296), .nC(nDCLK1), .C(DCLK1) );
	vdp_comp_we g5152 (.nZ(w5316), .A(w5203), .Z(w5317) );
	vdp_comp_we g5153 (.nZ(w5026), .A(w5203), .Z(w6613) );
	vdp_comp_we g5154 (.nZ(w5313), .A(w5203), .Z(w6614) );
	vdp_comp_we g5155 (.nZ(w5312), .A(w5203), .Z(w6615) );
	vdp_comp_we g5156 (.nZ(w5311), .A(w5203), .Z(w6616) );
	vdp_comp_we g5157 (.nZ(w5310), .A(w5203), .Z(w6617) );
	vdp_comp_we g5158 (.nZ(w5309), .A(w5203), .Z(w6618) );
	vdp_comp_we g5159 (.nZ(w5308), .A(w5203), .Z(w6619) );
	vdp_comp_we g5160 (.nZ(w5307), .A(w5203), .Z(w6620) );
	vdp_comp_we g5161 (.nZ(w6622), .A(w5203), .Z(w6621) );
	vdp_comp_we g5162 (.nZ(w4944), .A(w119), .Z(w4992) );
	vdp_noif0 g5163 (.A(w5246), .nZ(VRAMA[10]), .nE(w5169) );
	vdp_noif0 g5164 (.A(w5275), .nZ(VRAMA[13]), .nE(w5169) );
	vdp_noif0 g5165 (.A(w5305), .nZ(VRAMA[11]), .nE(w5169) );
	vdp_noif0 g5166 (.A(w5304), .nZ(VRAMA[12]), .nE(w5169) );
	vdp_not g5167 (.nZ(w5248), .A(VRAMA[2]) );
	vdp_not g5168 (.nZ(w5275), .A(w5274) );
	vdp_not g5169 (.nZ(w5303), .A(w124) );
	vdp_aoi22 g5170 (.Z(w5007), .B2(w5236), .B1(w5247), .A1(w5110), .A2(w5259) );
	vdp_aoi22 g5171 (.Z(w5246), .B2(w5236), .B1(w5272), .A1(w5110), .A2(w5251) );
	vdp_aoi22 g5172 (.Z(w5000), .B2(w5236), .B1(w5260), .A1(w5110), .A2(w6606) );
	vdp_aoi22 g5173 (.Z(w5305), .B2(w5236), .B1(w5273), .A1(w5110), .A2(w5271) );
	vdp_aoi22 g5174 (.Z(w5304), .B2(w5236), .B1(w5306), .A1(w5110), .A2(w5236) );
	vdp_and g5175 (.Z(w5302), .B(w5303), .A(w4580) );
	vdp_nor8 g5176 (.Z(w5245), .B(w5255), .A(w5256), .C(w5254), .D(w5253), .F(w5242), .E(w5238), .G(w5240), .H(w5241) );
	vdp_not g5177 (.nZ(w5318), .A(w123) );
	vdp_comp_str g5178 (.nZ(w5315), .A(w142), .Z(w5314) );
	vdp_comp_str g5179 (.nZ(w5277), .A(w143), .Z(w5276) );
	vdp_or3 g5180 (.Z(w5203), .B(w119), .A(w123), .C(w5302) );
	vdp_not g5181 (.nZ(S[7]), .A(w5293) );
	vdp_not g5182 (.nZ(S[6]), .A(w5292) );
	vdp_not g5183 (.nZ(S[5]), .A(w5291) );
	vdp_not g5184 (.nZ(S[4]), .A(w5290) );
	vdp_not g5185 (.nZ(S[3]), .A(w5289) );
	vdp_not g5186 (.nZ(S[2]), .A(w5288) );
	vdp_not g5187 (.nZ(S[1]), .A(w5287) );
	vdp_not g5188 (.nZ(S[0]), .A(w6404) );
	vdp_aon21_sr g5189 (.Q(w5394), .A1(w5393), .A2(w6507), .B(w6514), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5190 (.Q(w6514), .A1(w5361), .A2(w6507), .B(w6513), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5191 (.Q(w6513), .A1(w5360), .A2(w6507), .B(w6512), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5192 (.Q(w6512), .A1(w5359), .A2(w6507), .B(w6511), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5193 (.Q(w6511), .A1(w5358), .A2(w6507), .B(w6510), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5194 (.Q(w6510), .A1(w5357), .A2(w6507), .B(w6509), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5195 (.Q(w6509), .A1(w5356), .A2(w6507), .B(w6508), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5196 (.Q(w6508), .A1(w5355), .A2(w6507), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5197 (.Q(w6516), .A1(w5350), .A2(w6515), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5198 (.Q(w6517), .A1(w5349), .A2(w6515), .B(w6516), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5199 (.Q(w6518), .A1(w5348), .A2(w6515), .B(w6517), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5200 (.Q(w6519), .A1(w5347), .A2(w6515), .B(w6518), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5201 (.Q(w6520), .A1(w5346), .A2(w6515), .B(w6519), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5202 (.Q(w6521), .A1(w5345), .A2(w6515), .B(w6520), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5203 (.Q(w6522), .A1(w5344), .A2(w6515), .B(w6521), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5204 (.Q(w5375), .A1(w5364), .A2(w6515), .B(w6522), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5205 (.Q(w5503), .A1(w5339), .A2(w6499), .B(w6500), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5206 (.Q(w6500), .A1(w5338), .A2(w6499), .B(w6501), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5207 (.Q(w6501), .A1(w5337), .A2(w6499), .B(w6502), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5208 (.Q(w6502), .A1(w5336), .A2(w6499), .B(w6503), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5209 (.Q(w6503), .A1(w5335), .A2(w6499), .B(w6504), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5210 (.Q(w6504), .A1(w5334), .A2(w6499), .B(w6505), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5211 (.Q(w6505), .A1(w5333), .A2(w6499), .B(w6506), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5212 (.Q(w6506), .A1(w5332), .A2(w6499), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5213 (.Q(w6492), .A1(w5327), .A2(w6491), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5214 (.Q(w6493), .A1(w5326), .A2(w6491), .B(w6492), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5215 (.Q(w6494), .A1(w5325), .A2(w6491), .B(w6493), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5216 (.Q(w6495), .A1(w5324), .A2(w6491), .B(w6494), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5217 (.Q(w6497), .A1(w5402), .A2(w6491), .B(w6495), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5218 (.Q(w6496), .A1(w5407), .A2(w6491), .B(w6497), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5219 (.Q(w6498), .A1(w5401), .A2(w6491), .B(w6496), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5220 (.Q(w5323), .A1(w5322), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .A2(w6491), .B(w6498) );
	vdp_not g5221 (.nZ(w6499), .A(w5387) );
	vdp_not g5222 (.nZ(w6491), .A(w5387) );
	vdp_not g5223 (.nZ(w6515), .A(w5387) );
	vdp_not g5224 (.nZ(w6507), .A(w5387) );
	vdp_or4 g5225 (.Z(w5392), .B(w5353), .A(w5410), .D(w5388), .C(w5354) );
	vdp_or4 g5226 (.Z(w5379), .B(w5351), .A(w5382), .D(w5386), .C(w5352) );
	vdp_or4 g5227 (.Z(w5395), .B(w5363), .A(w5322), .D(w5745), .C(w5362) );
	vdp_or4 g5228 (.Z(w5378), .B(w5343), .A(w5741), .D(w5401), .C(w5342) );
	vdp_or4 g5229 (.Z(w5374), .B(w5341), .A(w5740), .D(w5407), .C(w5340) );
	vdp_or4 g5230 (.Z(w5398), .B(w5329), .A(w5328), .D(w6405), .C(w5330) );
	vdp_or4 g5231 (.Z(w5369), .B(w5367), .A(w5368), .D(w5331), .C(w5366) );
	vdp_slatch g5232 (.Q(w5388), .D(w5448), .nC(w5383), .C(w5384) );
	vdp_comp_str g5233 (.nZ(w5383), .A(w5418), .Z(w5384) );
	vdp_slatch g5234 (.Q(w5354), .D(w5446), .nC(w5383), .C(w5384) );
	vdp_slatch g5235 (.Q(w5353), .D(w5445), .nC(w5383), .C(w5384) );
	vdp_slatch g5236 (.Q(w5410), .D(w5444), .nC(w5383), .C(w5384) );
	vdp_slatch g5237 (.Q(w5386), .D(w5443), .nC(w5383), .C(w5384) );
	vdp_slatch g5238 (.Q(w5352), .D(w5442), .nC(w5383), .C(w5384) );
	vdp_slatch g5239 (.Q(w5351), .D(w5440), .nC(w5383), .C(w5384) );
	vdp_slatch g5240 (.Q(w5382), .D(w5436), .nC(w5383), .C(w5384) );
	vdp_slatch g5241 (.Q(w5331), .D(w6488), .nC(w5365), .C(w5400) );
	vdp_slatch g5242 (.Q(w5366), .D(w6489), .nC(w5365), .C(w5400) );
	vdp_slatch g5243 (.Q(w5367), .D(w6490), .nC(w5365), .C(w5400) );
	vdp_slatch g5244 (.Q(w5368), .D(w5424), .nC(w5365), .C(w5400) );
	vdp_slatch g5245 (.Q(w6405), .D(w5422), .nC(w5365), .C(w5400) );
	vdp_slatch g5246 (.Q(w5330), .D(w5421), .nC(w5365), .C(w5400) );
	vdp_slatch g5247 (.Q(w5329), .D(w5420), .nC(w5365), .C(w5400) );
	vdp_slatch g5248 (.Q(w5328), .D(w5417), .nC(w5365), .C(w5400) );
	vdp_aon22 g5249 (.Z(w5456), .B2(w5371), .B1(w5405), .A1(w5398), .A2(w5377) );
	vdp_comp_we g5250 (.nZ(w5371), .A(w5404), .Z(w5377) );
	vdp_notif0 g5251 (.A(w5399), .nZ(w170), .nE(w5416) );
	vdp_notif0 g5252 (.A(w5403), .nZ(w156), .nE(w5416) );
	vdp_notif0 g5253 (.A(w5372), .nZ(DB[10]), .nE(w5427) );
	vdp_notif0 g5254 (.A(w5373), .nZ(DB[2]), .nE(w5427) );
	vdp_notif0 g5255 (.A(w5381), .nZ(DB[1]), .nE(w5427) );
	vdp_notif0 g5256 (.A(w5408), .nZ(DB[9]), .nE(w5427) );
	vdp_notif0 g5257 (.A(w5390), .nZ(DB[8]), .nE(w5427) );
	vdp_notif0 g5258 (.A(w5391), .nZ(DB[0]), .nE(w5427) );
	vdp_not g5259 (.nZ(w5396), .A(w5395) );
	vdp_aon22 g5260 (.Z(w5429), .B2(w5371), .B1(w5376), .A1(w5369), .A2(w5377) );
	vdp_aon22 g5261 (.Z(w5434), .B2(w5371), .B1(w5380), .A1(w5379), .A2(w5377) );
	vdp_aon22 g5262 (.Z(w5451), .B2(w5371), .B1(w5396), .A1(w5392), .A2(w5377) );
	vdp_comp_str g5263 (.nZ(w5365), .A(w5418), .Z(w5400) );
	vdp_not g5264 (.nZ(w5405), .A(w5406) );
	vdp_not g5265 (.nZ(w5376), .A(w5374) );
	vdp_not g5266 (.nZ(w5380), .A(w5378) );
	vdp_and3 g5267 (.Z(w5841), .B(w5432), .A(w5379), .C(w5378) );
	vdp_and3 g5268 (.Z(w5438), .B(w5452), .A(w5392), .C(w5395) );
	vdp_and3 g5269 (.Z(w5454), .B(w5430), .A(w5369), .C(w5374) );
	vdp_and3 g5270 (.Z(w5798), .B(w5398), .A(w5411), .C(w5406) );
	vdp_aon2222 g5271 (.Z(w5403), .B2(w5324), .B1(w5414), .A1(w5415), .A2(w5326), .D2(w5322), .D1(w5412), .C1(w5413), .C2(w5407) );
	vdp_aon2222 g5272 (.Z(w5399), .B2(w5325), .B1(w5414), .A1(w5415), .A2(w5327), .D2(w5401), .D1(w5412), .C1(w5413), .C2(w5402) );
	vdp_aon2222 g5273 (.Z(w5372), .B2(w5334), .B1(w5414), .A1(w5415), .A2(w5332), .D2(w5338), .D1(w5412), .C1(w5413), .C2(w5336) );
	vdp_aon2222 g5274 (.Z(w5373), .B2(w5335), .B1(w5414), .A1(w5415), .A2(w5333), .D2(w5339), .D1(w5412), .C1(w5413), .C2(w5337) );
	vdp_aon2222 g5275 (.Z(w5381), .B2(w5347), .B1(w5414), .A1(w5415), .A2(w5349), .D2(w5364), .D1(w5412), .C1(w5413), .C2(w5345) );
	vdp_aon2222 g5276 (.Z(w5408), .B2(w5348), .B1(w5414), .A1(w5415), .A2(w5350), .D2(w5344), .D1(w5412), .C1(w5413), .C2(w5346) );
	vdp_aon2222 g5277 (.Z(w5390), .B2(w5357), .B1(w5414), .A1(w5415), .A2(w5355), .D2(w5361), .D1(w5412), .C1(w5413), .C2(w5359) );
	vdp_aon2222 g5278 (.Z(w5391), .B2(w5358), .B1(w5414), .A1(w5415), .A2(w5356), .D2(w5393), .D1(w5412), .C1(w5413), .C2(w5360) );
	vdp_slatch g5279 (.Q(w5448), .D(w5469), .nC(w5468), .C(w5447) );
	vdp_comp_str g5280 (.nZ(w5468), .A(w5467), .Z(w5447) );
	vdp_slatch g5281 (.Q(w5446), .D(w5473), .nC(w5468), .C(w5447) );
	vdp_slatch g5282 (.Q(w5445), .D(w5474), .nC(w5468), .C(w5447) );
	vdp_slatch g5283 (.Q(w5444), .D(w5477), .nC(w5468), .C(w5447) );
	vdp_slatch g5284 (.Q(w5443), .D(w5482), .nC(w5483), .C(w5441) );
	vdp_comp_str g5285 (.nZ(w5483), .A(w5478), .Z(w5441) );
	vdp_slatch g5286 (.Q(w5442), .D(w5485), .nC(w5483), .C(w5441) );
	vdp_slatch g5287 (.Q(w5440), .D(w5486), .nC(w5483), .C(w5441) );
	vdp_slatch g5288 (.Q(w5436), .D(w5488), .nC(w5483), .C(w5441) );
	vdp_sr_bit g5289 (.Q(w5490), .D(w5375), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5290 (.nQ(w5435), .D(w5493), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5291 (.nQ(w5495), .D(w5433), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5292 (.nQ(w5431), .D(w5502), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5293 (.nQ(w5508), .D(w5428), .nC(nDCLK2), .C(DCLK2) );
	vdp_slatch g5294 (.Q(w5424), .D(w5469), .nC(w5510), .C(w5426) );
	vdp_slatch g5295 (.Q(w6488), .D(w5473), .nC(w5510), .C(w5426) );
	vdp_slatch g5296 (.Q(w6489), .D(w5474), .nC(w5510), .C(w5426) );
	vdp_slatch g5297 (.Q(w6490), .D(w5477), .nC(w5510), .C(w5426) );
	vdp_comp_str g5298 (.nZ(w5510), .A(w5509), .Z(w5426) );
	vdp_slatch g5299 (.Q(w5422), .D(w5482), .nC(w5521), .C(w5419) );
	vdp_slatch g5300 (.Q(w5421), .D(w5485), .nC(w5521), .C(w5419) );
	vdp_slatch g5301 (.Q(w5420), .D(w5486), .nC(w5521), .C(w5419) );
	vdp_slatch g5302 (.Q(w5417), .D(w5488), .nC(w5521), .C(w5419) );
	vdp_comp_str g5303 (.nZ(w5521), .A(w5526), .Z(w5419) );
	vdp_dlatch_inv g5304 (.nQ(w5519), .D(w5518), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5305 (.nQ(w5522), .D(w6446), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5306 (.nQ(w5455), .D(w5525), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5307 (.Z(w5524), .B(w5455), .A(w5460) );
	vdp_xor g5308 (.Z(w6484), .B(w5431), .A(w5460) );
	vdp_xor g5309 (.Z(w5491), .B(w5435), .A(w5460) );
	vdp_xor g5310 (.Z(w6414), .B(w6413), .A(w5460) );
	vdp_sr_bit g5311 (.Q(w6487), .D(w5394), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5312 (.nQ(w6413), .D(w5458), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5313 (.nQ(w6415), .D(w5450), .nC(nDCLK2), .C(DCLK2) );
	vdp_and g5314 (.Z(w5452), .B(w6414), .A(w5461) );
	vdp_and g5315 (.Z(w5453), .B(w6415), .A(DCLK1) );
	vdp_and g5316 (.Z(w5437), .B(w5495), .A(DCLK1) );
	vdp_and g5317 (.Z(w5432), .B(w5491), .A(w5461) );
	vdp_and g5318 (.Z(w5412), .B(w5497), .A(w5496) );
	vdp_and g5319 (.Z(w5413), .B(w82), .A(w5497) );
	vdp_and g5320 (.Z(w5414), .B(w83), .A(w5496) );
	vdp_and g5321 (.Z(w5415), .B(w82), .A(w83) );
	vdp_and g5322 (.Z(w5430), .B(w6484), .A(w83) );
	vdp_and g5323 (.Z(w5449), .B(w5508), .A(DCLK1) );
	vdp_and g5324 (.Z(w5439), .B(w5522), .A(DCLK1) );
	vdp_and g5325 (.Z(w5411), .B(w5524), .A(w5461) );
	vdp_sr_bit g5326 (.Q(w5500), .D(w5503), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5327 (.Q(w5511), .D(w5480), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_not g5328 (.nZ(w5418), .A(w5425) );
	vdp_not g5329 (.nZ(w5423), .A(w4528) );
	vdp_not g5330 (.nZ(w5496), .A(w82) );
	vdp_not g5331 (.nZ(w5497), .A(w83) );
	vdp_aoi21 g5332 (.Z(w5450), .B(w5464), .A1(w5451), .A2(w5452) );
	vdp_aoi21 g5333 (.Z(w5433), .B(w5492), .A1(w5434), .A2(w5432) );
	vdp_aoi21 g5334 (.Z(w5428), .B(w5507), .A1(w5429), .A2(w5430) );
	vdp_oai21 g5335 (.Z(w5425), .B(DCLK2), .A1(w5512), .A2(w5511) );
	vdp_aoi21 g5336 (.Z(w6446), .B(w5507), .A1(w5411), .A2(w5456) );
	vdp_not g5337 (.nZ(w5416), .A(w121) );
	vdp_nand g5338 (.Z(w5480), .B(w5519), .A(w5423) );
	vdp_sr_bit g5339 (.Q(w5471), .D(w5528), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5340 (.Q(w5476), .D(w6416), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5341 (.Q(w5487), .D(w6486), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5342 (.Q(w5472), .D(w5489), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5343 (.Q(w5494), .D(w2725), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5344 (.Q(w5498), .D(w5499), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5345 (.Q(w6456), .D(w5515), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5346 (.Q(w5515), .D(w5527), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5347 (.Q(w5530), .D(w5323), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g5348 (.Z(w5527), .B2(w5323), .B1(w5534), .A1(w5533), .A2(w5530) );
	vdp_aon22 g5349 (.Z(w5499), .B2(w5503), .B1(w5534), .A1(w5533), .A2(w5500) );
	vdp_aon22 g5350 (.Z(w5489), .B2(w5375), .B1(w5534), .A1(w5533), .A2(w5490) );
	vdp_aon22 g5351 (.Z(w5528), .B2(w5394), .B1(w5534), .A1(w5533), .A2(w6487) );
	vdp_not g5352 (.nZ(w5470), .A(w5525) );
	vdp_not g5353 (.nZ(w5462), .A(w83) );
	vdp_not g5354 (.nZ(w5467), .A(w5546) );
	vdp_not g5355 (.nZ(w5475), .A(M5) );
	vdp_not g5356 (.nZ(w5478), .A(w5479) );
	vdp_not g5357 (.nZ(w5465), .A(w5539) );
	vdp_not g5358 (.nZ(w5459), .A(w5537) );
	vdp_not g5359 (.nZ(w5509), .A(w5506) );
	vdp_not g5360 (.nZ(w5526), .A(w5514) );
	vdp_not g5361 (.nZ(w5520), .A(w5515) );
	vdp_comp_we g5362 (.nZ(w5534), .A(M5), .Z(w5533) );
	vdp_and g5363 (.Z(w2844), .B(w5472), .A(w5471) );
	vdp_or g5364 (.Z(w6416), .B(w5471), .A(w5475) );
	vdp_or g5365 (.Z(w5481), .B(w5484), .A(w5480) );
	vdp_and g5366 (.Z(w6486), .B(w5472), .A(M5) );
	vdp_and g5367 (.Z(w2725), .B(w5498), .A(M5) );
	vdp_or g5368 (.Z(w5523), .B(w5480), .A(w5513) );
	vdp_not g5369 (.nZ(w5545), .A(SPR_PRIO) );
	vdp_bufif0 g5370 (.A(w6456), .Z(COL[0]), .nE(w5545) );
	vdp_oai21 g5371 (.Z(w5506), .B(DCLK2), .A1(w5481), .A2(w5505) );
	vdp_bufif0 g5372 (.A(w5494), .Z(COL[6]), .nE(w5545) );
	vdp_bufif0 g5373 (.A(w5487), .Z(COL[5]), .nE(w5545) );
	vdp_bufif0 g5374 (.A(w5476), .Z(COL[4]), .nE(w5545) );
	vdp_oai21 g5375 (.Z(w5479), .B(DCLK2), .A1(w5481), .A2(w5466) );
	vdp_oai21 g5376 (.Z(w5546), .B(DCLK2), .A1(w5540), .A2(w5466) );
	vdp_and3 g5377 (.Z(w5466), .B(w5544), .A(w5465), .C(w5543) );
	vdp_and3 g5378 (.Z(w5484), .B(w5544), .A(w5465), .C(w5531) );
	vdp_and3 g5379 (.Z(w5505), .B(w5543), .A(w5532), .C(w5465) );
	vdp_and3 g5380 (.Z(w5513), .B(w5531), .A(w5532), .C(w5465) );
	vdp_or4 g5381 (.Z(w2724), .B(w5536), .A(w5517), .D(w5515), .C(w5516) );
	vdp_and4 g5382 (.Z(w2785), .B(w5516), .A(w5536), .D(w5520), .C(w5517) );
	vdp_and4 g5383 (.Z(w2784), .B(w5516), .A(w5536), .D(w5515), .C(w5517) );
	vdp_oai21 g5384 (.Z(w5514), .B(DCLK2), .A1(w5505), .A2(w5523) );
	vdp_nand3 g5385 (.Z(w5458), .B(w5459), .A(w5470), .C(w5542) );
	vdp_nand3 g5386 (.Z(w5463), .B(w5541), .A(w120), .C(w5462) );
	vdp_nand3 g5387 (.Z(w5504), .B(w82), .A(w120), .C(w5462) );
	vdp_nand g5388 (.Z(w5507), .B(w5504), .A(w5535) );
	vdp_nand g5389 (.Z(w5501), .B(w5538), .A(w5537) );
	vdp_nand g5390 (.Z(w5502), .B(w5470), .A(w5501) );
	vdp_nand g5391 (.Z(w5493), .B(w5459), .A(w5470) );
	vdp_nand g5392 (.Z(w5464), .B(w5463), .A(w5535) );
	vdp_sr_bit g5393 (.Q(w6419), .D(w6418), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5394 (.Q(w6420), .D(w6419), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5395 (.Q(w5614), .D(w6420), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5396 (.Q(w5621), .D(w5614), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5397 (.Q(w5612), .D(w6421), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5398 (.Q(w6485), .D(w5622), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5399 (.Q(w5624), .D(w6523), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5400 (.Q(w5604), .D(w6417), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_dlatch_inv g5401 (.nQ(w5571), .D(w5562), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5402 (.nQ(w5576), .D(w5561), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5403 (.nQ(w5582), .D(w5560), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5404 (.nQ(w5587), .D(w5559), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5405 (.nQ(w5588), .D(w5558), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5406 (.nQ(w5591), .D(w5557), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5407 (.nQ(w5592), .D(w5556), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5408 (.nQ(w5595), .D(w5554), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5409 (.nQ(w5618), .D(w5619), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5410 (.nQ(w5616), .D(w5600), .nC(nDCLK1), .C(DCLK1) );
	vdp_cnt_bit_load g5411 (.Q(w5619), .D(w5620), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1), .R(1'b0), .CI(w6525), .L(w5551), .nL(w5597) );
	vdp_cnt_bit_load g5412 (.Q(w5600), .D(w5599), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1), .R(1'b0), .CI(w5552), .L(w5551), .nL(w5597), .CO(w6525) );
	vdp_aon22 g5413 (.Z(w5482), .B2(w5553), .B1(w170), .A1(w5595), .A2(w5572) );
	vdp_aon22 g5414 (.Z(w5554), .B2(w5555), .B1(w5584), .A1(w5583), .A2(w5575) );
	vdp_aon22 g5415 (.Z(w5485), .B2(w5553), .B1(DB[12]), .A1(w5592), .A2(w5572) );
	vdp_aon22 g5416 (.Z(w5556), .B2(w5555), .B1(w5580), .A1(w5581), .A2(w5575) );
	vdp_aon22 g5417 (.Z(w5563), .B2(w5553), .B1(DB[13]), .A1(w5591), .A2(w5572) );
	vdp_aon22 g5418 (.Z(w5557), .B2(w5555), .B1(w5573), .A1(w5574), .A2(w5575) );
	vdp_aon22 g5419 (.Z(w5488), .B2(w5553), .B1(DB[14]), .A1(w5588), .A2(w5572) );
	vdp_aon22 g5420 (.Z(w5558), .B2(w5555), .B1(w5564), .A1(w5565), .A2(w5575) );
	vdp_aon22 g5421 (.Z(w5469), .B2(w5553), .B1(w156), .A1(w5587), .A2(w5572) );
	vdp_aon22 g5422 (.Z(w5559), .B2(w5555), .B1(w5583), .A1(w5584), .A2(w5575) );
	vdp_aon22 g5423 (.Z(w5473), .B2(w5553), .B1(DB[4]), .A1(w5582), .A2(w5572) );
	vdp_aon22 g5424 (.Z(w5560), .B2(w5555), .B1(w5581), .A1(w5580), .A2(w5575) );
	vdp_aon22 g5425 (.Z(w5474), .B2(w5553), .B1(DB[5]), .A1(w5576), .A2(w5572) );
	vdp_aon22 g5426 (.Z(w5561), .B2(w5555), .B1(w5574), .A1(w5573), .A2(w5575) );
	vdp_aon22 g5427 (.Z(w5548), .B2(w5553), .B1(DB[6]), .A1(w5571), .A2(w5572) );
	vdp_aon22 g5428 (.Z(w5562), .B2(w5555), .B1(w5565), .A1(w5564), .A2(w5575) );
	vdp_slatch g5429 (.Q(w6417), .D(w5607), .nC(w5550), .C(w5608) );
	vdp_dlatch_inv g5430 (.nQ(w5605), .D(w5604), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5431 (.nQ(w5622), .D(w26), .nC(nHCLK1), .C(HCLK1) );
	vdp_xnor g5432 (.Z(w5532), .B(1'b0), .A(w5616) );
	vdp_xor g5433 (.Z(w5596), .B(w5604), .A(w5606) );
	vdp_aon22 g5434 (.Z(w6523), .B2(w5614), .B1(M5), .A1(w5621), .A2(w6524) );
	vdp_not g5435 (.nZ(w5623), .A(w5622) );
	vdp_not g5436 (.nZ(w6524), .A(M5) );
	vdp_not g5437 (.nZ(w5550), .A(w5608) );
	vdp_not g5438 (.nZ(w6418), .A(w5611) );
	vdp_not g5439 (.nZ(w5531), .A(w5605) );
	vdp_not g5440 (.nZ(w5539), .A(w5618) );
	vdp_not g5441 (.nZ(w5552), .A(w5608) );
	vdp_comp_we g5442 (.nZ(w5572), .A(w4528), .Z(w5553) );
	vdp_comp_we g5443 (.nZ(w5575), .A(w5596), .Z(w5555) );
	vdp_comp_we g5444 (.nZ(w5597), .A(w5608), .Z(w5551) );
	vdp_and g5445 (.Z(w6421), .B(w6485), .A(w5623) );
	vdp_aoi21 g5446 (.Z(w5611), .B(w25), .A1(M5), .A2(w22) );
	vdp_sr_bit g5447 (.Q(w5606), .D(w5670), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_aon22 g5448 (.Z(w5678), .B2(w5672), .B1(w5671), .A1(w5668), .A2(w5615) );
	vdp_aon22 g5449 (.Z(w5677), .B2(w5672), .B1(w5675), .A1(w5673), .A2(w5615) );
	vdp_aon22 g5450 (.Z(w5674), .B2(w5672), .B1(w5673), .A1(w5675), .A2(w5615) );
	vdp_aon22 g5451 (.Z(w5679), .B2(w5672), .B1(w5668), .A1(w5671), .A2(w5615) );
	vdp_not g5452 (.nZ(w5634), .A(w5671) );
	vdp_not g5453 (.nZ(w5635), .A(w5675) );
	vdp_not g5454 (.nZ(w5640), .A(w5673) );
	vdp_not g5455 (.nZ(w5639), .A(w5668) );
	vdp_not g5456 (.nZ(w5567), .A(w5677) );
	vdp_not g5457 (.nZ(w5568), .A(w5678) );
	vdp_not g5458 (.nZ(w5569), .A(w5679) );
	vdp_not g5459 (.nZ(w5570), .A(w5674) );
	vdp_not g5460 (.nZ(w5613), .A(M5) );
	vdp_comp_we g5461 (.nZ(w5672), .A(w5606), .Z(w5615) );
	vdp_not g5462 (.nZ(w5608), .A(w5669) );
	vdp_not g5463 (.nZ(w5667), .A(w5666) );
	vdp_dlatch_inv g5464 (.nQ(w5666), .D(w5665), .nC(nHCLK1), .C(HCLK1) );
	vdp_aon2222 g5465 (.Z(w5566), .B2(w5568), .B1(w5628), .A1(w5627), .A2(w5567), .D2(w5570), .D1(w5646), .C1(w5644), .C2(w5569) );
	vdp_aon2222 g5466 (.Z(w5617), .B2(w5640), .B1(w5632), .A1(w5639), .A2(w5627), .D2(w5634), .D1(w5636), .C1(w5635), .C2(w5680) );
	vdp_aon2222 g5467 (.Z(w5586), .B2(w5568), .B1(w5633), .A1(w5632), .A2(w5567), .D2(w5570), .D1(w5637), .C1(w5645), .C2(w5569) );
	vdp_aon2222 g5468 (.Z(w5577), .B2(w5640), .B1(w5633), .A1(w5639), .A2(w5628), .D2(w5634), .D1(w5648), .C1(w5635), .C2(w5641) );
	vdp_aon2222 g5469 (.Z(w5594), .B2(w5568), .B1(w5641), .A1(w5680), .A2(w5567), .D2(w5570), .D1(w5643), .C1(w5642), .C2(w5569) );
	vdp_aon2222 g5470 (.Z(w5585), .B2(w5640), .B1(w5645), .A1(w5639), .A2(w5644), .D2(w5634), .D1(w5647), .C1(w5635), .C2(w5642) );
	vdp_aon2222 g5471 (.Z(w5603), .B2(w5568), .B1(w5648), .A1(w5636), .A2(w5567), .D2(w5570), .D1(w5649), .C1(w5647), .C2(w5569) );
	vdp_aon2222 g5472 (.Z(w5589), .B2(w5640), .B1(w5637), .A1(w5639), .A2(w5646), .D2(w5634), .D1(w5649), .C1(w5635), .C2(w5643) );
	vdp_aon2222 g5473 (.Z(w5578), .B2(w5568), .B1(w5651), .A1(w5650), .A2(w5567), .D2(w5570), .D1(w5663), .C1(w5652), .C2(w5569) );
	vdp_aon2222 g5474 (.Z(w5593), .B2(w5640), .B1(w5653), .A1(w5639), .A2(w5650), .D2(w5634), .D1(w5654), .C1(w5635), .C2(w5655) );
	vdp_aon2222 g5475 (.Z(w5590), .B2(w5568), .B1(w5657), .A1(w5653), .A2(w5567), .D2(w5570), .D1(w5656), .C1(w5658), .C2(w5569) );
	vdp_aon2222 g5476 (.Z(w5601), .B2(w5640), .B1(w5657), .A1(w5639), .A2(w5651), .D2(w5634), .D1(w5659), .C1(w5635), .C2(w5660) );
	vdp_aon2222 g5477 (.Z(w5590), .B2(w5568), .B1(w5660), .A1(w5655), .A2(w5567), .D2(w5570), .D1(w5661), .C1(w5662), .C2(w5569) );
	vdp_aon2222 g5478 (.Z(w5602), .B2(w5640), .B1(w5658), .A1(w5639), .A2(w5652), .D2(w5634), .D1(w5664), .C1(w5635), .C2(w5662) );
	vdp_aon2222 g5479 (.Z(w5610), .B2(w5568), .B1(w5659), .A1(w5654), .A2(w5567), .D2(w5570), .D1(w5676), .C1(w5664), .C2(w5569) );
	vdp_aon2222 g5480 (.Z(w5609), .B2(w5640), .B1(w5656), .A1(w5639), .A2(w5663), .D2(w5634), .D1(w5676), .C1(w5635), .C2(w5661) );
	vdp_aoi22 g5481 (.Z(w5564), .B2(w5626), .B1(w5566), .A1(w5579), .A2(w5617) );
	vdp_aoi22 g5482 (.Z(w5573), .B2(w5626), .B1(w5578), .A1(w5579), .A2(w5577) );
	vdp_aoi22 g5483 (.Z(w5580), .B2(w5626), .B1(w5586), .A1(w5579), .A2(w5585) );
	vdp_aoi22 g5484 (.Z(w5584), .B2(w5626), .B1(w5590), .A1(w5579), .A2(w5589) );
	vdp_aoi22 g5485 (.Z(w5565), .B2(w5626), .B1(w5594), .A1(w5579), .A2(w5593) );
	vdp_aoi22 g5486 (.Z(w5574), .B2(w5626), .B1(w5590), .A1(w5579), .A2(w5601) );
	vdp_aoi22 g5487 (.Z(w5581), .B2(w5626), .B1(w5603), .A1(w5579), .A2(w5602) );
	vdp_aoi22 g5488 (.Z(w5583), .B2(w5626), .B1(w5610), .A1(w5579), .A2(w5609) );
	vdp_nand g5489 (.Z(w5669), .B(w5667), .A(HCLK2) );
	vdp_nor g5490 (.Z(w5626), .B(w5613), .A(w5612) );
	vdp_nor g5491 (.Z(w5579), .B(M5), .A(w5612) );
	vdp_sr_bit g5492 (.Q(w5671), .D(w5675), .nC2(w5682), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5493 (.Q(w5675), .D(w5673), .nC2(w5682), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5494 (.Q(w5673), .D(w5668), .nC2(w5682), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5495 (.Q(w5668), .D(w5669), .nC2(w5682), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_dlatch_inv g5496 (.nQ(w5512), .D(w5671), .nC(nDCLK1), .C(DCLK1) );
	vdp_comp_str g5497 (.nZ(w5631), .A(w5683), .Z(w5685) );
	vdp_comp_str g5498 (.nZ(w5630), .A(w5683), .Z(w5688) );
	vdp_comp_str g5499 (.nZ(w5638), .A(w5683), .Z(w5689) );
	vdp_comp_str g5500 (.nZ(w5629), .A(w5683), .Z(w5684) );
	vdp_slatch g5501 (.D(w5698), .Q(w5627), .nC(w5629), .C(w5684) );
	vdp_slatch g5502 (.D(w6549), .Q(w5628), .nC(w5638), .C(w5689) );
	vdp_slatch g5503 (.D(w6548), .Q(w5644), .nC(w5630), .C(w5688) );
	vdp_slatch g5504 (.D(w6547), .Q(w5646), .nC(w5631), .C(w5685) );
	vdp_slatch g5505 (.D(w5697), .Q(w5632), .nC(w5629), .C(w5684) );
	vdp_slatch g5506 (.D(w6546), .Q(w5633), .nC(w5638), .C(w5689) );
	vdp_slatch g5507 (.D(w6545), .Q(w5645), .nC(w5630), .C(w5688) );
	vdp_slatch g5508 (.D(w6544), .Q(w5637), .nC(w5631), .C(w5685) );
	vdp_slatch g5509 (.D(w5696), .Q(w5680), .nC(w5629), .C(w5684) );
	vdp_slatch g5510 (.D(w6543), .Q(w5641), .nC(w5638), .C(w5689) );
	vdp_slatch g5511 (.D(w6542), .Q(w5642), .nC(w5630), .C(w5688) );
	vdp_slatch g5512 (.D(w6541), .Q(w5643), .nC(w5631), .C(w5685) );
	vdp_slatch g5513 (.D(w5695), .Q(w5636), .nC(w5629), .C(w5684) );
	vdp_slatch g5514 (.D(w6540), .Q(w5648), .nC(w5638), .C(w5689) );
	vdp_slatch g5515 (.D(w6539), .Q(w5647), .nC(w5630), .C(w5688) );
	vdp_slatch g5516 (.D(w6538), .Q(w5649), .nC(w5631), .C(w5685) );
	vdp_slatch g5517 (.D(w5694), .Q(w5650), .nC(w5629), .C(w5684) );
	vdp_slatch g5518 (.D(w6537), .Q(w5651), .nC(w5638), .C(w5689) );
	vdp_slatch g5519 (.D(w6536), .Q(w5652), .nC(w5630), .C(w5688) );
	vdp_slatch g5520 (.D(w6535), .Q(w5663), .nC(w5631), .C(w5685) );
	vdp_slatch g5521 (.D(w5693), .Q(w5653), .nC(w5629), .C(w5684) );
	vdp_slatch g5522 (.D(w6534), .Q(w5657), .nC(w5638), .C(w5689) );
	vdp_slatch g5523 (.D(w6533), .Q(w5658), .nC(w5630), .C(w5688) );
	vdp_slatch g5524 (.D(w6532), .Q(w5656), .nC(w5631), .C(w5685) );
	vdp_slatch g5525 (.D(w5692), .Q(w5655), .nC(w5629), .C(w5684) );
	vdp_slatch g5526 (.D(w6531), .Q(w5660), .nC(w5638), .C(w5689) );
	vdp_slatch g5527 (.D(w6530), .Q(w5662), .nC(w5630), .C(w5688) );
	vdp_slatch g5528 (.D(w6529), .Q(w5661), .nC(w5631), .C(w5685) );
	vdp_slatch g5529 (.D(w5691), .Q(w5654), .nC(w5629), .C(w5684) );
	vdp_slatch g5530 (.D(w6528), .Q(w5659), .nC(w5638), .C(w5689) );
	vdp_slatch g5531 (.D(w6527), .Q(w5664), .nC(w5630), .C(w5688) );
	vdp_slatch g5532 (.D(w6526), .nC(w5631), .C(w5685), .Q(w5676) );
	vdp_sr_bit g5533 (.Q(w5700), .D(w5701), .nC2(nDCLK1), .nC1(w5682), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g5534 (.Q(w6422), .D(w5700), .nC2(nDCLK1), .nC1(w5682), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g5535 (.Q(w5714), .D(w6422), .nC2(nDCLK1), .nC1(w5682), .C2(DCLK1), .C1(DCLK2) );
	vdp_comp_str g5536 (.nZ(w5704), .A(w5715), .Z(w5690) );
	vdp_comp_str g5537 (.nZ(w5707), .A(w5715), .Z(w5687) );
	vdp_comp_str g5538 (.nZ(w5709), .A(w5715), .Z(w5686) );
	vdp_dlatch_inv g5539 (.nQ(w5701), .D(w5710), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g5540 (.Z(w5683), .B(DCLK2), .A(w5714) );
	vdp_and g5541 (.Z(w5715), .B(DCLK2), .A(w5700) );
	vdp_and g5542 (.Z(w5716), .B(DCLK2), .A(w5701) );
	vdp_slatch g5543 (.Q(w6528), .D(w6552), .nC(w5704), .C(w5690) );
	vdp_slatch g5544 (.Q(w6527), .D(w6551), .nC(w5707), .C(w5687) );
	vdp_slatch g5545 (.Q(w6526), .D(w6550), .nC(w5709), .C(w5686) );
	vdp_slatch g5546 (.Q(w6531), .D(w6555), .nC(w5704), .C(w5690) );
	vdp_slatch g5547 (.Q(w6530), .D(w6554), .nC(w5707), .C(w5687) );
	vdp_slatch g5548 (.Q(w6529), .D(w6553), .nC(w5709), .C(w5686) );
	vdp_slatch g5549 (.Q(w6534), .D(w6558), .nC(w5704), .C(w5690) );
	vdp_slatch g5550 (.Q(w6533), .D(w6557), .nC(w5707), .C(w5687) );
	vdp_slatch g5551 (.Q(w6532), .D(w6556), .nC(w5709), .C(w5686) );
	vdp_slatch g5552 (.Q(w6537), .D(w6561), .nC(w5704), .C(w5690) );
	vdp_slatch g5553 (.Q(w6536), .D(w6560), .nC(w5707), .C(w5687) );
	vdp_slatch g5554 (.Q(w6535), .D(w6559), .nC(w5709), .C(w5686) );
	vdp_slatch g5555 (.Q(w6540), .D(w6564), .nC(w5704), .C(w5690) );
	vdp_slatch g5556 (.Q(w6539), .D(w6563), .nC(w5707), .C(w5687) );
	vdp_slatch g5557 (.Q(w6538), .D(w6562), .nC(w5709), .C(w5686) );
	vdp_slatch g5558 (.Q(w6543), .D(w6567), .nC(w5704), .C(w5690) );
	vdp_slatch g5559 (.Q(w6542), .D(w6566), .nC(w5707), .C(w5687) );
	vdp_slatch g5560 (.Q(w6541), .D(w6565), .nC(w5709), .C(w5686) );
	vdp_slatch g5561 (.Q(w6546), .D(w6570), .nC(w5704), .C(w5690) );
	vdp_slatch g5562 (.Q(w6545), .D(w6569), .nC(w5707), .C(w5687) );
	vdp_slatch g5563 (.Q(w6544), .D(w6568), .nC(w5709), .C(w5686) );
	vdp_slatch g5564 (.Q(w6549), .D(w6573), .nC(w5704), .C(w5690) );
	vdp_slatch g5565 (.Q(w6548), .D(w6572), .nC(w5707), .C(w5687) );
	vdp_slatch g5566 (.Q(w6547), .D(w6571), .nC(w5709), .C(w5686) );
	vdp_sr_bit g5567 (.Q(w5713), .D(w5712), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_dlatch_inv g5568 (.nQ(w5712), .D(w5711), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g5569 (.Z(w5723), .B(w5712), .A(DCLK2) );
	vdp_nand g5570 (.Z(w5711), .B(w5614), .A(HCLK1) );
	vdp_nand g5571 (.Z(w5710), .B(w5624), .A(HCLK1) );
	vdp_and g5572 (.Z(w5722), .B(w5713), .A(DCLK2) );
	vdp_comp_str g5573 (.nZ(w5708), .A(w5723), .Z(w5721) );
	vdp_comp_str g5574 (.nZ(w5706), .A(w5722), .Z(w5720) );
	vdp_comp_str g5575 (.nZ(w5705), .A(w5716), .Z(w5719) );
	vdp_comp_str g5576 (.nZ(w5703), .A(w5715), .Z(w5718) );
	vdp_slatch g5577 (.D(S[7]), .Q(w5698), .nC(w5703), .C(w5718) );
	vdp_slatch g5578 (.D(S[7]), .Q(w6573), .nC(w5705), .C(w5719) );
	vdp_slatch g5579 (.D(S[7]), .Q(w6572), .nC(w5706), .C(w5720) );
	vdp_slatch g5580 (.D(S[7]), .Q(w6571), .nC(w5708), .C(w5721) );
	vdp_slatch g5581 (.D(S[5]), .Q(w5697), .nC(w5703), .C(w5718) );
	vdp_slatch g5582 (.D(S[5]), .Q(w6570), .nC(w5705), .C(w5719) );
	vdp_slatch g5583 (.D(S[5]), .Q(w6569), .nC(w5706), .C(w5720) );
	vdp_slatch g5584 (.D(S[5]), .Q(w6568), .nC(w5708), .C(w5721) );
	vdp_slatch g5585 (.D(S[3]), .Q(w5696), .nC(w5703), .C(w5718) );
	vdp_slatch g5586 (.D(S[3]), .Q(w6567), .nC(w5705), .C(w5719) );
	vdp_slatch g5587 (.D(S[3]), .Q(w6566), .nC(w5706), .C(w5720) );
	vdp_slatch g5588 (.D(S[3]), .Q(w6565), .nC(w5708), .C(w5721) );
	vdp_slatch g5589 (.D(S[1]), .Q(w5695), .nC(w5703), .C(w5718) );
	vdp_slatch g5590 (.D(S[1]), .Q(w6564), .nC(w5705), .C(w5719) );
	vdp_slatch g5591 (.D(S[1]), .Q(w6563), .nC(w5706), .C(w5720) );
	vdp_slatch g5592 (.D(S[1]), .Q(w6562), .nC(w5708), .C(w5721) );
	vdp_slatch g5593 (.D(S[6]), .Q(w5694), .nC(w5703), .C(w5718) );
	vdp_slatch g5594 (.D(S[6]), .Q(w6561), .nC(w5705), .C(w5719) );
	vdp_slatch g5595 (.D(S[6]), .Q(w6560), .nC(w5706), .C(w5720) );
	vdp_slatch g5596 (.D(S[6]), .Q(w6559), .nC(w5708), .C(w5721) );
	vdp_slatch g5597 (.D(S[4]), .Q(w5693), .nC(w5703), .C(w5718) );
	vdp_slatch g5598 (.D(S[4]), .Q(w6558), .nC(w5705), .C(w5719) );
	vdp_slatch g5599 (.D(S[4]), .Q(w6557), .nC(w5706), .C(w5720) );
	vdp_slatch g5600 (.D(S[4]), .Q(w6556), .nC(w5708), .C(w5721) );
	vdp_slatch g5601 (.D(S[2]), .Q(w5692), .nC(w5703), .C(w5718) );
	vdp_slatch g5602 (.D(S[2]), .Q(w6555), .nC(w5705), .C(w5719) );
	vdp_slatch g5603 (.D(S[2]), .Q(w6554), .nC(w5706), .C(w5720) );
	vdp_slatch g5604 (.D(S[2]), .Q(w6553), .nC(w5708), .C(w5721) );
	vdp_slatch g5605 (.D(S[0]), .Q(w5691), .nC(w5703), .C(w5718) );
	vdp_slatch g5606 (.D(S[0]), .Q(w6552), .nC(w5705), .C(w5719) );
	vdp_slatch g5607 (.D(S[0]), .Q(w6551), .nC(w5706), .C(w5720) );
	vdp_slatch g5608 (.D(S[0]), .nC(w5708), .C(w5721), .Q(w6550) );
	vdp_aon21_sr g5609 (.Q(w5779), .A1(w5738), .A2(w6749), .B(w6460), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5610 (.Q(w6460), .A1(w5342), .A2(w6749), .B(w6461), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5611 (.Q(w6461), .A1(w5340), .A2(w6749), .B(w6462), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5612 (.Q(w6462), .A1(w5739), .A2(w6749), .B(w6463), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5613 (.Q(w6463), .A1(w5768), .A2(w6749), .B(w6464), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5614 (.Q(w6464), .A1(w5730), .A2(w6749), .B(w6459), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5615 (.Q(w6459), .A1(w5731), .A2(w6749), .B(w6458), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5616 (.Q(w6458), .A1(w5732), .A2(w6749), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5617 (.Q(w6471), .A1(w5734), .A2(w6750), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5618 (.Q(w6470), .A1(w5735), .A2(w6750), .B(w6471), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5619 (.Q(w6469), .A1(w5749), .A2(w6750), .B(w6470), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5620 (.Q(w6468), .A1(w5736), .A2(w6750), .B(w6469), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5621 (.Q(w6467), .A1(w5737), .A2(w6750), .B(w6468), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5622 (.Q(w6466), .A1(w5341), .A2(w6750), .B(w6467), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5623 (.Q(w6465), .A1(w5343), .A2(w6750), .B(w6466), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5624 (.Q(w5783), .A1(w5362), .A2(w6750), .B(w6465), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5625 (.Q(w5788), .A1(w5745), .A2(w6751), .B(w6478), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5626 (.Q(w6478), .A1(w5741), .A2(w6751), .B(w6477), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5627 (.Q(w6477), .A1(w5740), .A2(w6751), .B(w6476), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5628 (.Q(w6476), .A1(w5747), .A2(w6751), .B(w6475), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5629 (.Q(w6475), .A1(w5748), .A2(w6751), .B(w6474), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5630 (.Q(w6474), .A1(w5750), .A2(w6751), .B(w6473), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5631 (.Q(w6473), .A1(w5762), .A2(w6751), .B(w6472), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5632 (.Q(w6472), .A1(w5763), .A2(w6751), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_or4 g5633 (.Z(w5771), .B(w5768), .A(w5324), .C(w5736), .D(w5748) );
	vdp_or4 g5634 (.Z(w5406), .B(w5739), .A(w5402), .C(w5737), .D(w5747) );
	vdp_aon22 g5635 (.Z(w5758), .B2(w4529), .B1(w5765), .A1(w5793), .A2(DB[0]) );
	vdp_aon22 g5636 (.Z(w5757), .B2(w4530), .B1(w5765), .A1(w5793), .A2(DB[1]) );
	vdp_aon22 g5637 (.Z(w5756), .B2(w4538), .B1(w5765), .A1(w5793), .A2(DB[2]) );
	vdp_aon22 g5638 (.Z(w5755), .B2(w4529), .B1(w5765), .A1(w5793), .A2(DB[8]) );
	vdp_aon22 g5639 (.Z(w5754), .B2(w4530), .B1(w5765), .A1(w5793), .A2(DB[9]) );
	vdp_aon22 g5640 (.Z(w5753), .B2(w4538), .B1(w5765), .A1(w5793), .A2(DB[10]) );
	vdp_or4 g5641 (.Z(w5780), .B(w5728), .A(w5729), .C(w5733), .D(w5767) );
	vdp_or4 g5642 (.Z(w5772), .B(w5742), .A(w5770), .C(w5743), .D(w5769) );
	vdp_or4 g5643 (.Z(w5787), .B(w5731), .A(w5326), .C(w5735), .D(w5762) );
	vdp_or4 g5644 (.Z(w5784), .B(w5749), .A(w5750), .C(w5730), .D(w5325) );
	vdp_or4 g5645 (.Z(w5794), .B(w5744), .A(w5746), .C(w5752), .D(w5751) );
	vdp_or4 g5646 (.Z(w5785), .B(w5760), .A(w5761), .C(w5764), .D(w5759) );
	vdp_or4 g5647 (.Z(w5796), .B(w5732), .A(w5327), .C(w5734), .D(w5763) );
	vdp_comp_we g5648 (.nZ(w5765), .A(w4528), .Z(w5793) );
	vdp_not g5649 (.nZ(w6749), .A(w5387) );
	vdp_not g5650 (.nZ(w6750), .A(w5387) );
	vdp_not g5651 (.nZ(w6751), .A(w5387) );
	vdp_slatch g5652 (.Q(w5769), .D(w5811), .nC(w5777), .C(w5810) );
	vdp_comp_str g5653 (.nZ(w5777), .A(w5418), .Z(w5810) );
	vdp_slatch g5654 (.Q(w5743), .D(w5813), .nC(w5777), .C(w5810) );
	vdp_slatch g5655 (.Q(w5742), .D(w5814), .nC(w5777), .C(w5810) );
	vdp_slatch g5656 (.Q(w5770), .D(w5815), .nC(w5777), .C(w5810) );
	vdp_slatch g5657 (.Q(w5729), .D(w5816), .nC(w5777), .C(w5810) );
	vdp_slatch g5658 (.Q(w5728), .D(w5818), .nC(w5777), .C(w5810) );
	vdp_slatch g5659 (.Q(w5733), .D(w5819), .nC(w5777), .C(w5810) );
	vdp_slatch g5660 (.Q(w5767), .D(w5820), .nC(w5777), .C(w5810) );
	vdp_slatch g5661 (.Q(w5759), .D(w5829), .nC(w5791), .C(w5828) );
	vdp_comp_str g5662 (.nZ(w5791), .A(w5418), .Z(w5828) );
	vdp_slatch g5663 (.Q(w5764), .D(w5831), .nC(w5791), .C(w5828) );
	vdp_slatch g5664 (.Q(w5760), .D(w5832), .nC(w5791), .C(w5828) );
	vdp_slatch g5665 (.Q(w5761), .D(w5833), .nC(w5791), .C(w5828) );
	vdp_slatch g5666 (.Q(w5746), .D(w5834), .nC(w5791), .C(w5828) );
	vdp_slatch g5667 (.Q(w5744), .D(w5836), .nC(w5791), .C(w5828) );
	vdp_slatch g5668 (.Q(w5752), .D(w5837), .nC(w5791), .C(w5828) );
	vdp_slatch g5669 (.Q(w5751), .D(w5838), .nC(w5791), .C(w5828) );
	vdp_comp_we g5670 (.nZ(w5774), .A(1'b0), .Z(w5404) );
	vdp_aon22 g5671 (.Z(w5840), .B2(w5774), .B1(w5795), .A1(w5794), .A2(w5404) );
	vdp_not g5672 (.nZ(w5387), .A(w4540) );
	vdp_not g5673 (.nZ(w5795), .A(w5796) );
	vdp_not g5674 (.nZ(w5786), .A(w5787) );
	vdp_not g5675 (.nZ(w5782), .A(w5784) );
	vdp_not g5676 (.nZ(w5773), .A(w5771) );
	vdp_and3 g5677 (.Z(w5800), .B(w5799), .A(w5772), .C(w5771) );
	vdp_aon22 g5678 (.Z(w5808), .B2(w5774), .B1(w5773), .A1(w5772), .A2(w5404) );
	vdp_notif0 g5679 (.A(w5775), .nZ(DB[4]), .nE(w5776) );
	vdp_aon2222 g5680 (.Z(w5775), .B2(w5768), .B1(w5806), .A1(w5807), .A2(w5731), .D2(w5738), .D1(w5804), .C1(w5805), .C2(w5340) );
	vdp_notif0 g5681 (.A(w5778), .nZ(DB[12]), .nE(w5776) );
	vdp_aon2222 g5682 (.Z(w5778), .B2(w5730), .B1(w5806), .A1(w5807), .A2(w5732), .D2(w5342), .D1(w5804), .C1(w5805), .C2(w5739) );
	vdp_notif0 g5683 (.A(w6455), .nZ(DB[13]), .nE(w5776) );
	vdp_aon2222 g5684 (.Z(w6455), .B2(w5749), .B1(w5806), .A1(w5807), .A2(w5734), .D2(w5343), .D1(w5804), .C1(w5805), .C2(w5737) );
	vdp_notif0 g5685 (.A(w5781), .nZ(DB[5]), .nE(w5776) );
	vdp_aon2222 g5686 (.Z(w5781), .B2(w5736), .B1(w5806), .A1(w5807), .A2(w5735), .D2(w5362), .D1(w5804), .C1(w5805), .C2(w5341) );
	vdp_notif0 g5687 (.A(w5790), .nZ(DB[14]), .nE(w5776) );
	vdp_aon2222 g5688 (.Z(w5790), .B2(w5750), .B1(w5806), .A1(w5807), .A2(w5763), .D2(w5741), .D1(w5804), .C1(w5805), .C2(w5747) );
	vdp_notif0 g5689 (.A(w5789), .nZ(DB[6]), .nE(w5776) );
	vdp_aon2222 g5690 (.Z(w5789), .B2(w5748), .B1(w5806), .A1(w5807), .A2(w5762), .D2(w5745), .D1(w5804), .C1(w5805), .C2(w5740) );
	vdp_aon22 g5691 (.Z(w5821), .B2(w5774), .B1(w5782), .A1(w5780), .A2(w5404) );
	vdp_aon22 g5692 (.Z(w5824), .B2(w5774), .B1(w5786), .A1(w5785), .A2(w5404) );
	vdp_and3 g5693 (.Z(w5802), .B(w5823), .A(w5780), .C(w5784) );
	vdp_and3 g5694 (.Z(w5803), .B(w5825), .A(w5785), .C(w5787) );
	vdp_and3 g5695 (.Z(w5801), .B(w5839), .A(w5794), .C(w5796) );
	vdp_not g5696 (.nZ(w5776), .A(w121) );
	vdp_slatch g5697 (.Q(w5834), .D(w5482), .nC(w5869), .C(w5835) );
	vdp_slatch g5698 (.Q(w5836), .D(w5485), .nC(w5869), .C(w5835) );
	vdp_slatch g5699 (.Q(w5837), .D(w5486), .nC(w5869), .C(w5835) );
	vdp_slatch g5700 (.Q(w5838), .D(w5488), .nC(w5869), .C(w5835) );
	vdp_comp_str g5701 (.nZ(w5869), .A(w5870), .Z(w5835) );
	vdp_slatch g5702 (.Q(w5829), .D(w5469), .nC(w5865), .C(w5830) );
	vdp_slatch g5703 (.Q(w5831), .D(w5473), .nC(w5865), .C(w5830) );
	vdp_slatch g5704 (.Q(w5832), .D(w5474), .nC(w5865), .C(w5830) );
	vdp_slatch g5705 (.Q(w5833), .D(w5548), .nC(w5865), .C(w5830) );
	vdp_comp_str g5706 (.nZ(w5865), .A(w5868), .Z(w5830) );
	vdp_slatch g5707 (.Q(w5816), .D(w5482), .nC(w5852), .C(w5817) );
	vdp_slatch g5708 (.Q(w5818), .D(w5485), .nC(w5852), .C(w5817) );
	vdp_slatch g5709 (.Q(w5819), .D(w5486), .nC(w5852), .C(w5817) );
	vdp_slatch g5710 (.Q(w5820), .D(w5488), .nC(w5852), .C(w5817) );
	vdp_comp_str g5711 (.nZ(w5852), .A(w6746), .Z(w5817) );
	vdp_slatch g5712 (.Q(w5811), .D(w5469), .nC(w5851), .C(w5812) );
	vdp_slatch g5713 (.Q(w5813), .D(w5473), .nC(w5851), .C(w5812) );
	vdp_slatch g5714 (.Q(w5814), .D(w5474), .nC(w5851), .C(w5812) );
	vdp_slatch g5715 (.Q(w5815), .D(w5548), .nC(w5851), .C(w5812) );
	vdp_comp_str g5716 (.nZ(w5851), .A(w5849), .Z(w5812) );
	vdp_dlatch_inv g5717 (.nQ(w6454), .D(w5844), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5718 (.Z(w5846), .B(w5460), .A(w6454) );
	vdp_sr_bit g5719 (.Q(w126), .D(w6452), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g5720 (.Q(w5843), .D(w5779), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5721 (.nQ(w5848), .D(w5809), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5722 (.nQ(w6447), .D(w5822), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5723 (.nQ(w6449), .D(w5858), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5724 (.Z(w6448), .B(w6449), .A(w5460) );
	vdp_sr_bit g5725 (.Q(w6457), .D(w5783), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5726 (.nQ(w5826), .D(w6744), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5727 (.Z(w6450), .B(w5826), .A(w5460) );
	vdp_sr_bit g5728 (.Q(w5862), .D(w5788), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5729 (.nQ(w5859), .D(w6453), .nC(nDCLK2), .C(DCLK2) );
	vdp_not g5730 (.nZ(w5874), .A(w5460) );
	vdp_not g5731 (.nZ(w5827), .A(w83) );
	vdp_not g5732 (.nZ(w5863), .A(w82) );
	vdp_dlatch_inv g5733 (.nQ(w5872), .D(w6451), .nC(nDCLK2), .C(DCLK2) );
	vdp_and g5734 (.Z(w5839), .B(w5874), .A(w5461) );
	vdp_aoi21 g5735 (.Z(w6451), .B(w5860), .A1(w5840), .A2(w5839) );
	vdp_and g5736 (.Z(w5725), .B(w5872), .A(DCLK1) );
	vdp_and g5737 (.Z(w5726), .B(w5859), .A(DCLK1) );
	vdp_and g5738 (.Z(w5825), .B(w6450), .A(w5461) );
	vdp_aoi21 g5739 (.Z(w6453), .B(w5860), .A1(w5824), .A2(w5825) );
	vdp_and g5740 (.Z(w5823), .B(w6448), .A(w5461) );
	vdp_aoi21 g5741 (.Z(w5822), .B(w5847), .A1(w5821), .A2(w5823) );
	vdp_and g5742 (.Z(w5799), .B(w5461), .A(w5846) );
	vdp_aoi21 g5743 (.Z(w5809), .B(w5847), .A1(w5808), .A2(w5799) );
	vdp_and g5744 (.Z(w5766), .B(DCLK1), .A(w5848) );
	vdp_and g5745 (.Z(w5727), .B(w6447), .A(DCLK1) );
	vdp_and g5746 (.Z(w5804), .B(w5827), .A(w5863) );
	vdp_and g5747 (.Z(w5806), .B(w83), .A(w5863) );
	vdp_and g5748 (.Z(w5805), .B(w5827), .A(w82) );
	vdp_and g5749 (.Z(w5807), .B(w83), .A(w82) );
	vdp_or8 g5750 (.Z(w6452), .B(w5800), .A(w5454), .C(w5801), .D(w5841), .F(w5803), .E(w5798), .G(w5438), .H(w5802) );
	vdp_sr_bit g5751 (.Q(w5517), .D(w5881), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5752 (.Q(w5845), .D(w5517), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5753 (.Q(w5516), .D(w5857), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5754 (.Q(w5875), .D(w5516), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5755 (.Q(w5536), .D(w6438), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5756 (.Q(w5864), .D(w5536), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_comp_we g5757 (.nZ(w5879), .A(M5), .Z(w5878) );
	vdp_not g5758 (.nZ(w5870), .A(w5871) );
	vdp_or g5759 (.Z(w5540), .B(w5873), .A(w5480) );
	vdp_and3 g5760 (.Z(w5873), .B(w5532), .A(w5539), .C(w5531) );
	vdp_and3 g5761 (.Z(w5867), .B(w5532), .A(w5539), .C(w5543) );
	vdp_and3 g5762 (.Z(w6744), .B(w5537), .A(w5525), .C(w5538) );
	vdp_and3 g5763 (.Z(w5854), .B(w5544), .A(w5539), .C(w5531) );
	vdp_and3 g5764 (.Z(w5876), .B(w5544), .A(w5539), .C(w5543) );
	vdp_aoi21 g5765 (.Z(w5844), .B(w5470), .A1(w5459), .A2(w5542) );
	vdp_aon22 g5766 (.Z(w5881), .B2(w5779), .B1(w5879), .A1(w5878), .A2(w5843) );
	vdp_aon22 g5767 (.Z(w5857), .B2(w5783), .B1(w5879), .A1(w5878), .A2(w6457) );
	vdp_aon22 g5768 (.Z(w6438), .B2(w5788), .B1(w5879), .A1(w5878), .A2(w5862) );
	vdp_bufif0 g5769 (.A(w5875), .Z(COL[2]), .nE(w5880) );
	vdp_oai21 g5770 (.Z(w5855), .B(DCLK2), .A1(w5876), .A2(w5856) );
	vdp_and g5771 (.Z(w5858), .B(w5537), .A(w5525) );
	vdp_or g5772 (.Z(w5876), .B(w5854), .A(w5480) );
	vdp_bufif0 g5773 (.A(w5864), .Z(COL[3]), .nE(w5880) );
	vdp_oai21 g5774 (.Z(w5866), .B(DCLK2), .A1(w5856), .A2(w5867) );
	vdp_oai21 g5775 (.Z(w5871), .B(DCLK2), .A1(w5867), .A2(w5540) );
	vdp_not g5776 (.nZ(w5543), .A(w5531) );
	vdp_not g5777 (.nZ(w5868), .A(w5866) );
	vdp_not g5778 (.nZ(w5541), .A(w82) );
	vdp_not g5779 (.nZ(w5544), .A(w5532) );
	vdp_not g5780 (.nZ(w6746), .A(w5855) );
	vdp_not g5781 (.nZ(w5542), .A(w5538) );
	vdp_not g5782 (.nZ(w5849), .A(w5850) );
	vdp_bufif0 g5783 (.A(w5845), .Z(COL[1]), .nE(w5880) );
	vdp_oai21 g5784 (.Z(w5850), .B(DCLK2), .A1(w5523), .A2(w5876) );
	vdp_not g5785 (.nZ(w5880), .A(SPR_PRIO) );
	vdp_nand3 g5786 (.Z(w5853), .B(w120), .A(w83), .C(w5541) );
	vdp_nand g5787 (.Z(w5847), .B(w5535), .A(w5853) );
	vdp_nand3 g5788 (.Z(w5861), .B(w120), .A(w83), .C(w82) );
	vdp_nand g5789 (.Z(w5860), .B(w5535), .A(w5861) );
	vdp_sr_bit g5790 (.Q(w5908), .D(w5949), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5791 (.Q(w5909), .D(w5947), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5792 (.Q(w5906), .D(w5954), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5793 (.Q(w5907), .D(w5946), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5794 (.Z(w4535), .B2(w5908), .B1(w5943), .A1(w5942), .A2(w81), .C1(w5897), .C2(w5909) );
	vdp_aon222 g5795 (.Z(w4534), .B2(w5906), .B1(w5943), .A1(w5942), .A2(w80), .C1(w5897), .C2(w5907) );
	vdp_sr_bit g5796 (.Q(w5904), .D(w5953), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5797 (.Q(w5905), .D(w5945), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5798 (.Z(w4533), .B2(w5904), .B1(w5943), .A1(w5942), .A2(w79), .C1(w5897), .C2(w5905) );
	vdp_sr_bit g5799 (.Q(w5902), .D(w5952), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5800 (.Q(w5903), .D(w5944), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5801 (.Z(w4532), .B2(w5902), .B1(w5943), .A1(w5942), .A2(w78), .C1(w5897), .C2(w5903) );
	vdp_sr_bit g5802 (.Q(w5898), .D(w5951), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5803 (.Q(w5901), .D(w5955), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5804 (.Z(w4531), .B2(w5898), .B1(w5943), .A1(w5942), .A2(w77), .C1(w5897), .C2(w5901) );
	vdp_sr_bit g5805 (.Q(w5899), .D(w5950), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5806 (.Q(w5900), .D(w5941), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5807 (.Z(w4536), .B2(w5899), .B1(w5943), .A1(w5942), .A2(w76), .C1(w5897), .C2(w5900) );
	vdp_sr_bit g5808 (.Q(w5525), .D(w6723), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_slatch g5809 (.Q(w6723), .D(w5620), .nC(w5933), .C(w5894) );
	vdp_sr_bit g5810 (.Q(w5537), .D(w6721), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_slatch g5811 (.Q(w6721), .D(w5599), .nC(w5933), .C(w5894) );
	vdp_sr_bit g5812 (.Q(w5538), .D(w6722), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_slatch g5813 (.Q(w6722), .D(w5607), .nC(w5933), .C(w5894) );
	vdp_sr_bit g5814 (.Q(w5910), .D(w26), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5815 (.Q(w5893), .D(w5910), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5816 (.Q(w5892), .D(w5938), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5817 (.Q(w5926), .D(w5936), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5818 (.Q(w5925), .D(w5935), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5819 (.Q(w5889), .D(w4540), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5820 (.Q(w5888), .D(w5921), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5821 (.Q(w5916), .D(w6481), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5822 (.Q(w6481), .D(w5957), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_xor g5823 (.Z(w5918), .B(w5916), .A(w5917) );
	vdp_dlatch_inv g5824 (.nQ(w5887), .D(w5921), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5825 (.nQ(w5919), .D(w5918), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5826 (.nQ(w5890), .D(w5891), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5827 (.nQ(w5924), .D(w5923), .nC(nHCLK1), .C(HCLK1) );
	vdp_comp_str g5828 (.nZ(w5933), .A(w5930), .Z(w5894) );
	vdp_oai21 g5829 (.Z(w6480), .B(w5920), .A1(w5957), .A2(w5916) );
	vdp_and g5830 (.Z(w4529), .B(w5914), .A(w5886) );
	vdp_not g5831 (.nZ(w5460), .A(w5919) );
	vdp_not g5832 (.nZ(w5921), .A(w6480) );
	vdp_and g5833 (.Z(w4530), .B(w5913), .A(w5886) );
	vdp_and g5834 (.Z(w4538), .B(w5912), .A(w5886) );
	vdp_or g5835 (.Z(w5922), .B(w5888), .A(w5921) );
	vdp_not g5836 (.nZ(w5940), .A(w4528) );
	vdp_not g5837 (.nZ(w4540), .A(w5923) );
	vdp_not g5838 (.nZ(w5956), .A(M5) );
	vdp_not g5839 (.nZ(w5943), .A(w6714) );
	vdp_not g5840 (.nZ(w5895), .A(w5894) );
	vdp_not g5841 (.nZ(w5942), .A(w5940) );
	vdp_not g5842 (.nZ(w5897), .A(w5896) );
	vdp_or4 g5843 (.Z(w4537), .B(w4540), .A(w4528), .C(w5889), .D(w5922) );
	vdp_or4 g5844 (.Z(w5923), .B(w5926), .A(w5886), .C(w5892), .D(w5925) );
	vdp_nand g5845 (.Z(w5891), .B(w5924), .A(HCLK2) );
	vdp_nand g5846 (.Z(w5535), .B(w5940), .A(w5890) );
	vdp_nor g5847 (.Z(w5461), .B(w5887), .A(w4528) );
	vdp_nand g5848 (.Z(w5896), .B(w5940), .A(w5895) );
	vdp_nand g5849 (.Z(w6714), .B(w5940), .A(w5886) );
	vdp_aoi22 g5850 (.Z(w5886), .B2(w5956), .B1(w26), .A1(M5), .A2(w5893) );
	vdp_cnt_bit_load g5851 (.Q(w5985), .D(w5934), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w7), .CI(w6047), .L(w5932), .nL(w5978) );
	vdp_cnt_bit_load g5852 (.Q(w5931), .D(w5982), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w7), .CI(w5927), .L(w5932), .nL(w5978), .CO(w6047) );
	vdp_sr_bit g5853 (.Q(w5920), .D(w6445), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5854 (.SUM(w5938), .CO(w6702), .CI(1'b1), .A(HPOS[0]), .B(M5) );
	vdp_fa g5855 (.SUM(w5936), .CO(w6703), .CI(w6702), .A(HPOS[1]), .B(1'b0) );
	vdp_fa g5856 (.SUM(w5935), .CO(w6704), .CI(w6703), .A(HPOS[2]), .B(1'b1) );
	vdp_fa g5857 (.SUM(w5941), .CO(w6705), .CI(w6704), .A(w5990), .B(M5) );
	vdp_fa g5858 (.SUM(w5955), .CO(w6706), .CI(w6705), .A(HPOS[4]), .B(w5994) );
	vdp_fa g5859 (.SUM(w5944), .CO(w6707), .CI(w6706), .A(HPOS[5]), .B(1'b1) );
	vdp_fa g5860 (.SUM(w5945), .CO(w6708), .CI(w6707), .A(HPOS[6]), .B(1'b1) );
	vdp_fa g5861 (.SUM(w5946), .CO(w6709), .CI(w6708), .A(HPOS[7]), .B(1'b1) );
	vdp_fa g5862 (.SUM(w5947), .CI(w6709), .A(HPOS[8]), .B(1'b1) );
	vdp_not g5863 (.nZ(w5994), .A(M5) );
	vdp_aoi33 g5864 (.Z(w6445), .B2(w6720), .B1(w5949), .A1(H40), .A2(w5949), .A3(w5948), .B3(w6720) );
	vdp_not g5865 (.nZ(w6720), .A(H40) );
	vdp_or g5866 (.Z(w5948), .B(w5953), .A(w5954) );
	vdp_and g5867 (.Z(w5929), .B(w5927), .A(w5928) );
	vdp_sr_bit g5868 (.Q(w5927), .D(w6479), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5869 (.Q(w6479), .D(w5665), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5870 (.nQ(w5975), .D(w5512), .nC(nDCLK2), .C(DCLK2) );
	vdp_slatch g5871 (.Q(w5974), .D(w5961), .nC(w5915), .C(w5965) );
	vdp_slatch g5872 (.Q(w5914), .D(w5974), .nC(w5911), .C(w5967) );
	vdp_slatch g5873 (.Q(w5968), .D(w5960), .nC(w5915), .C(w5965) );
	vdp_slatch g5874 (.Q(w5912), .D(w5968), .nC(w5911), .C(w5967) );
	vdp_slatch g5875 (.Q(w5969), .D(w5961), .nC(w5915), .C(w5965) );
	vdp_slatch g5876 (.Q(w5913), .D(w5969), .nC(w5911), .C(w5967) );
	vdp_slatch g5877 (.Q(w6482), .D(w5670), .nC(w5915), .C(w5965) );
	vdp_sr_bit g5878 (.Q(w5917), .D(w6482), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_and g5879 (.Z(w5959), .B(DCLK2), .A(w5512) );
	vdp_comp_str g5880 (.nZ(w5911), .A(w5959), .Z(w5967) );
	vdp_comp_str g5881 (.nZ(w5915), .A(w5930), .Z(w5965) );
	vdp_not g5882 (.nZ(w5957), .A(w5975) );
	vdp_comp_we g5883 (.nZ(w5978), .A(w5929), .Z(w5932) );
	vdp_and3 g5884 (.Z(w5930), .B(HCLK1), .A(w5928), .C(w5927) );
	vdp_nand g5885 (.Z(w5982), .B(w5963), .A(M5) );
	vdp_nand g5886 (.Z(w5934), .B(w5962), .A(M5) );
	vdp_nor g5887 (.Z(w5928), .B(w5985), .A(w5931) );
	vdp_fa g5888 (.SUM(w5949), .CI(w6004), .A(w6003), .B(w6016) );
	vdp_aon22 g5889 (.Z(w6003), .B2(w6008), .B1(w6002), .A1(w6040), .A2(w5971) );
	vdp_sr_bit g5890 (.Q(w6002), .D(w5949), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5891 (.Q(w6040), .D(w6041), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5892 (.SUM(w6041), .CI(w6000), .A(w6001), .B(w6036) );
	vdp_aon22 g5893 (.Z(w6001), .B2(w6013), .B1(w6039), .A1(1'b0), .A2(w5964) );
	vdp_fa g5894 (.SUM(w5954), .CO(w6004), .CI(w5999), .A(w5998), .B(w6016) );
	vdp_aon22 g5895 (.Z(w5998), .B2(w6008), .B1(w5997), .A1(w6037), .A2(w5971) );
	vdp_sr_bit g5896 (.Q(w5997), .D(w5954), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5897 (.Q(w6037), .D(w6043), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5898 (.SUM(w6043), .CO(w6000), .CI(w5996), .A(w5995), .B(w6036) );
	vdp_aon22 g5899 (.Z(w5995), .B2(w6013), .B1(w6034), .A1(w6035), .A2(w5964) );
	vdp_fa g5900 (.SUM(w5953), .CO(w5999), .CI(w5993), .A(w5992), .B(w6016) );
	vdp_aon22 g5901 (.Z(w5992), .B2(w6008), .B1(w5991), .A1(w6033), .A2(w5971) );
	vdp_fa g5902 (.SUM(w6044), .CO(w5996), .CI(w5989), .A(w5988), .B(w6019) );
	vdp_aon22 g5903 (.Z(w5988), .B2(w6013), .B1(w6031), .A1(w6032), .A2(w5964) );
	vdp_sr_bit g5904 (.Q(w5991), .D(w5953), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5905 (.Q(w6033), .D(w6044), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5906 (.SUM(w6005), .CO(w5993), .CI(w6006), .A(w5987), .B(w6016) );
	vdp_aon22 g5907 (.Z(w5987), .B2(w6008), .B1(w5986), .A1(w6030), .A2(w5971) );
	vdp_sr_bit g5908 (.Q(w5986), .D(w6005), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5909 (.Q(w6030), .D(w6029), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5910 (.SUM(w6029), .CO(w5989), .CI(w5983), .A(w5984), .B(w6019) );
	vdp_aon22 g5911 (.Z(w5984), .B2(w6013), .B1(w6717), .A1(w6028), .A2(w5964) );
	vdp_fa g5912 (.SUM(w5951), .CO(w6006), .CI(w5980), .A(w5981), .B(w6016) );
	vdp_aon22 g5913 (.Z(w5981), .B2(w6008), .B1(w5979), .A1(w6027), .A2(w5971) );
	vdp_sr_bit g5914 (.Q(w5979), .D(w5951), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5915 (.Q(w6027), .D(w6710), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5916 (.SUM(w6710), .CO(w5983), .CI(w5977), .A(w5976), .B(w6026) );
	vdp_aon22 g5917 (.Z(w5976), .B2(w6013), .B1(w6045), .A1(w6025), .A2(w5964) );
	vdp_fa g5918 (.SUM(w5950), .CO(w5980), .CI(w5973), .A(w5972), .B(w6016) );
	vdp_aon22 g5919 (.Z(w5972), .B2(w6008), .B1(w5970), .A1(w6024), .A2(w5971) );
	vdp_sr_bit g5920 (.Q(w5970), .D(w5950), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5921 (.Q(w6024), .D(w6023), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5922 (.SUM(w6023), .CO(w5977), .CI(w6021), .A(w5966), .B(w6018) );
	vdp_aon22 g5923 (.Z(w5966), .B2(w6013), .B1(w6020), .A1(w6022), .A2(w5964) );
	vdp_aon22 g5924 (.Z(w5620), .B2(w6013), .B1(w6017), .A1(w6042), .A2(w5964) );
	vdp_aon22 g5925 (.Z(w5599), .B2(w6013), .B1(w6012), .A1(w6015), .A2(w5964) );
	vdp_aon22 g5926 (.Z(w5607), .B2(w6013), .B1(w6011), .A1(w6014), .A2(w5964) );
	vdp_and g5927 (.Z(w5973), .B(w6010), .A(w6716) );
	vdp_comp_we g5928 (.nZ(w5964), .A(M5), .Z(w6013) );
	vdp_comp_we g5929 (.nZ(w6008), .A(w6715), .Z(w5971) );
	vdp_sr_bit g5930 (.Q(w6715), .D(w5930), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5931 (.Q(w6009), .D(w5975), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5932 (.Q(w6057), .D(w6060), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5933 (.Q(w6060), .D(w6061), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5934 (.Q(w6061), .D(w6065), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5935 (.Q(w6065), .D(w6066), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5936 (.Q(w6066), .D(w6067), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5937 (.nQ(w6067), .D(w6070), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5938 (.nZ(w6017), .A(w6057) );
	vdp_sr_bit g5939 (.Q(w6071), .D(w6072), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5940 (.Q(w6072), .D(w6076), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5941 (.Q(w6076), .D(w6077), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5942 (.Q(w6077), .D(w6079), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5943 (.Q(w6079), .D(w6082), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5944 (.nQ(w6082), .D(w6081), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5945 (.nZ(w6020), .A(w6071) );
	vdp_sr_bit g5946 (.Q(w6083), .D(w6483), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5947 (.Q(w6483), .D(w6086), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5948 (.Q(w6086), .D(w6088), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5949 (.Q(w6088), .D(w6089), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5950 (.Q(w6089), .D(w6090), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5951 (.nQ(w6090), .D(w6094), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5952 (.nZ(w6045), .A(w6083) );
	vdp_sr_bit g5953 (.Q(w6095), .D(w6098), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5954 (.Q(w6098), .D(w6102), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5955 (.Q(w6102), .D(w6101), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5956 (.Q(w6101), .D(w6103), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5957 (.Q(w6103), .D(w6106), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5958 (.nQ(w6106), .D(w6107), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5959 (.nZ(w6717), .A(w6095) );
	vdp_sr_bit g5960 (.Q(w6110), .D(w6113), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5961 (.Q(w6113), .D(w6114), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5962 (.Q(w6114), .D(w6115), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5963 (.Q(w6115), .D(w6139), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5964 (.Q(w6139), .D(w6140), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5965 (.nQ(w6140), .D(w6120), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5966 (.nZ(w6031), .A(w6110) );
	vdp_sr_bit g5967 (.Q(w6141), .D(w6135), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5968 (.Q(w6135), .D(w6134), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5969 (.Q(w6134), .D(w6132), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5970 (.Q(w6132), .D(w6131), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5971 (.Q(w6131), .D(w6129), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5972 (.nQ(w6129), .D(w6119), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5973 (.nZ(w6034), .A(w6141) );
	vdp_sr_bit g5974 (.Q(w6718), .D(w6125), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5975 (.Q(w6125), .D(w6126), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5976 (.Q(w6126), .D(w6122), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5977 (.Q(w6122), .D(w6121), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5978 (.Q(w6121), .D(w6117), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5979 (.nQ(w6117), .D(w6118), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5980 (.nZ(w6039), .A(w6718) );
	vdp_and g5981 (.Z(w6016), .B(w6010), .A(w5917) );
	vdp_and g5982 (.Z(w6053), .B(w5670), .A(w5963) );
	vdp_and g5983 (.Z(w6054), .B(w6021), .A(w5962) );
	vdp_or g5984 (.Z(w6018), .B(w6053), .A(w6019) );
	vdp_and g5985 (.B(w6056), .A(M5) );
	vdp_or g5986 (.Z(w6026), .B(w6054), .A(w6019) );
	vdp_and g5987 (.Z(w6019), .B(w23), .A(w6727) );
	vdp_or g5988 (.Z(w6036), .B(w6019), .A(M5) );
	vdp_not g5989 (.nZ(w6727), .A(M5) );
	vdp_not g5990 (.nZ(w6716), .A(w5917) );
	vdp_nor g5991 (.Z(w6010), .B(w6715), .A(w6009) );
	vdp_sr_bit g5992 (.Q(w6069), .D(w6073), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5993 (.Q(w6073), .D(w6074), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5994 (.Q(w6074), .D(w6075), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5995 (.Q(w6075), .D(w6078), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5996 (.Q(w6078), .D(w6719), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5997 (.nQ(w6719), .D(w6148), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5998 (.nZ(w5961), .A(w6069) );
	vdp_sr_bit g5999 (.Q(w6058), .D(w6059), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6000 (.Q(w6059), .D(w6062), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6001 (.Q(w6062), .D(w6063), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6002 (.Q(w6063), .D(w6064), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6003 (.Q(w6064), .D(w6068), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6004 (.nQ(w6068), .D(w6147), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6005 (.nZ(w5961), .A(w6058) );
	vdp_sr_bit g6006 (.Q(w6048), .D(w6049), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6007 (.Q(w6049), .D(w6050), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6008 (.Q(w6050), .D(w6052), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6009 (.Q(w6052), .D(w6051), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6010 (.Q(w6051), .D(w6055), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6011 (.nQ(w6055), .D(w6146), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6012 (.nZ(w6056), .A(w6048) );
	vdp_sr_bit g6013 (.Q(w6080), .D(w6084), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6014 (.Q(w6084), .D(w6085), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6015 (.Q(w6085), .D(w6087), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6016 (.Q(w6087), .D(w6091), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6017 (.Q(w6091), .D(w6092), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6018 (.nQ(w6092), .D(w6153), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6019 (.nZ(w5960), .A(w6080) );
	vdp_sr_bit g6020 (.Q(w6093), .D(w6096), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6021 (.Q(w6096), .D(w6097), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6022 (.Q(w6097), .D(w6099), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6023 (.Q(w6099), .D(w6100), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6024 (.Q(w6100), .D(w6104), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6025 (.nQ(w6104), .D(w6149), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6026 (.nZ(w5963), .A(w6093) );
	vdp_sr_bit g6027 (.Q(w6105), .D(w6108), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6028 (.Q(w6108), .D(w6109), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6029 (.Q(w6109), .D(w6111), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6030 (.Q(w6111), .D(w6112), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6031 (.Q(w6112), .D(w6116), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6032 (.nQ(w6116), .D(w6150), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6033 (.nZ(w5962), .A(w6105) );
	vdp_sr_bit g6034 (.Q(w6137), .D(w6138), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6035 (.Q(w6138), .D(w6142), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6036 (.Q(w6142), .D(w6143), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6037 (.Q(w6143), .D(w6136), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6038 (.Q(w6136), .D(w6133), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6039 (.nQ(w6133), .D(w6151), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6040 (.nZ(w6011), .A(w6137) );
	vdp_sr_bit g6041 (.Q(w6128), .D(w6130), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6042 (.Q(w6130), .D(w6127), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6043 (.Q(w6127), .D(w6124), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6044 (.Q(w6124), .D(w6123), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6045 (.Q(w6123), .D(w6144), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6046 (.nQ(w6144), .D(w6152), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6047 (.nZ(w6012), .A(w6128) );
	vdp_slatch g6048 (.D(w6178), .nC(w6216), .C(w6156), .nQ(w6014) );
	vdp_slatch g6049 (.D(S[1]), .nC(w6217), .C(w6160), .Q(w6177) );
	vdp_slatch g6050 (.D(S[1]), .nC(w6218), .C(w6159), .Q(w6176) );
	vdp_aoi22 g6051 (.Z(w6175), .B2(w6222), .B1(w6177), .A1(w6176), .A2(w6157) );
	vdp_slatch g6052 (.D(S[0]), .nC(w6217), .C(w6160), .Q(w6180) );
	vdp_slatch g6053 (.D(S[0]), .nC(w6218), .C(w6159), .Q(w6179) );
	vdp_aoi22 g6054 (.Z(w6178), .B2(w6222), .B1(w6180), .A1(w6179), .A2(w6157) );
	vdp_slatch g6055 (.D(w6175), .nC(w6216), .C(w6156), .nQ(w6015) );
	vdp_slatch g6056 (.D(S[2]), .nC(w6217), .C(w6160), .Q(w6174) );
	vdp_slatch g6057 (.D(S[2]), .nC(w6218), .C(w6159), .Q(w6173) );
	vdp_aoi22 g6058 (.Z(w6259), .B2(w6222), .B1(w6174), .A1(w6173), .A2(w6157) );
	vdp_slatch g6059 (.D(w6259), .nC(w6216), .C(w6156), .nQ(w6042) );
	vdp_slatch g6060 (.D(S[3]), .nC(w6217), .C(w6160), .Q(w6172) );
	vdp_slatch g6061 (.D(S[3]), .nC(w6218), .C(w6159), .Q(w6171) );
	vdp_aoi22 g6062 (.Z(w6170), .B2(w6222), .B1(w6172), .A1(w6171), .A2(w6157) );
	vdp_slatch g6063 (.D(w6170), .nC(w6216), .C(w6156), .nQ(w6022) );
	vdp_slatch g6064 (.D(S[4]), .nC(w6217), .C(w6160), .Q(w6169) );
	vdp_slatch g6065 (.D(S[4]), .nC(w6218), .C(w6159), .Q(w6168) );
	vdp_aoi22 g6066 (.Z(w6167), .B2(w6222), .B1(w6169), .A1(w6168), .A2(w6157) );
	vdp_slatch g6067 (.D(w6167), .nC(w6216), .C(w6156), .nQ(w6025) );
	vdp_slatch g6068 (.D(S[5]), .nC(w6217), .C(w6160), .Q(w6166) );
	vdp_slatch g6069 (.D(S[5]), .nC(w6218), .C(w6159), .Q(w6165) );
	vdp_aoi22 g6070 (.Z(w6164), .B2(w6222), .B1(w6166), .A1(w6165), .A2(w6157) );
	vdp_slatch g6071 (.D(w6164), .nC(w6216), .C(w6156), .nQ(w6028) );
	vdp_slatch g6072 (.D(S[6]), .nC(w6217), .C(w6160), .Q(w6163) );
	vdp_slatch g6073 (.D(S[6]), .nC(w6218), .C(w6159), .Q(w6161) );
	vdp_aoi22 g6074 (.Z(w6162), .B2(w6222), .B1(w6163), .A1(w6161), .A2(w6157) );
	vdp_slatch g6075 (.D(w6162), .nC(w6216), .C(w6156), .nQ(w6032) );
	vdp_slatch g6076 (.D(S[7]), .nC(w6217), .C(w6160), .Q(w6158) );
	vdp_slatch g6077 (.D(S[7]), .nC(w6218), .C(w6159), .Q(w6154) );
	vdp_aoi22 g6078 (.Z(w6155), .B2(w6222), .B1(w6158), .A1(w6154), .A2(w6157) );
	vdp_slatch g6079 (.D(w6155), .nC(w6216), .C(w6156), .nQ(w6035) );
	vdp_comp_str g6080 (.nZ(w6216), .A(w5665), .Z(w6156) );
	vdp_comp_str g6081 (.nZ(w6217), .A(w4995), .Z(w6160) );
	vdp_comp_str g6082 (.nZ(w6218), .A(w4999), .Z(w6159) );
	vdp_comp_we g6083 (.nZ(w6222), .A(w6215), .Z(w6157) );
	vdp_sr_bit g6084 (.Q(w6213), .D(w6209), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6085 (.Z(w6209), .B(w6214), .A(w6181) );
	vdp_fa g6086 (.SUM(w6214), .CI(w6183), .A(w6213), .B(1'b0) );
	vdp_sr_bit g6087 (.Q(w6248), .D(w6204), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6088 (.Z(w6204), .B(w6210), .A(w6181) );
	vdp_fa g6089 (.SUM(w6210), .CO(w6183), .CI(w6184), .A(w6248), .B(1'b0) );
	vdp_sr_bit g6090 (.Q(w6205), .D(w6228), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6091 (.Z(w6228), .B(w6206), .A(w6181) );
	vdp_fa g6092 (.SUM(w6206), .CO(w6184), .CI(w6186), .A(w6205), .B(w6185) );
	vdp_sr_bit g6093 (.Q(w6201), .D(w6200), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6094 (.Z(w6200), .B(w6202), .A(w6181) );
	vdp_fa g6095 (.SUM(w6202), .CO(w6186), .CI(w6188), .A(w6201), .B(w6187) );
	vdp_sr_bit g6096 (.Q(w6191), .D(w6724), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6097 (.Q(w6724), .D(w22), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6098 (.nQ(w6189), .D(w6191), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g6099 (.nQ(w6181), .D(w6190), .nC(nHCLK1), .C(HCLK1) );
	vdp_and g6100 (.Z(w6185), .B(w6188), .A(w6197) );
	vdp_and g6101 (.Z(w6187), .B(w6188), .A(w6196) );
	vdp_and g6102 (.Z(w4618), .B(w6724), .A(w6273) );
	vdp_or g6103 (.Z(w6190), .B(w6194), .A(w6260) );
	vdp_not g6104 (.nZ(w6193), .A(M5) );
	vdp_not g6105 (.nZ(w6188), .A(w6189) );
	vdp_fa g6106 (.SUM(w6233), .CO(w6236), .CI(w6234), .A(w6287), .B(w6207) );
	vdp_aoi22 g6107 (.Z(w6299), .B2(w6219), .B1(w6235), .A1(w6233), .A2(w6283) );
	vdp_notif0 g6108 (.A(w6299), .nZ(VRAMA[9]), .nE(w6276) );
	vdp_fa g6109 (.SUM(w6224), .CO(w6234), .CI(w6230), .A(w6286), .B(w6211) );
	vdp_aoi22 g6110 (.Z(w6232), .B2(w6219), .B1(w6233), .A1(w6224), .A2(w6283) );
	vdp_notif0 g6111 (.A(w6232), .nZ(VRAMA[8]), .nE(w6276) );
	vdp_fa g6112 (.SUM(w6220), .CO(w6230), .CI(w6223), .A(w6285), .B(w6203) );
	vdp_aoi22 g6113 (.Z(w6231), .B2(w6219), .B1(w6224), .A1(w6220), .A2(w6283) );
	vdp_notif0 g6114 (.A(w6231), .nZ(VRAMA[7]), .nE(w6276) );
	vdp_fa g6115 (.SUM(w6226), .CO(w6223), .CI(1'b0), .A(w6284), .B(w6199) );
	vdp_aoi22 g6116 (.Z(w6221), .B2(w6219), .B1(w6220), .A1(w6226), .A2(w6283) );
	vdp_notif0 g6117 (.A(w6221), .nZ(VRAMA[6]), .nE(w6276) );
	vdp_not g6118 (.nZ(w6276), .A(w6290) );
	vdp_ha g6119 (.SUM(w6235), .B(w6288), .A(w6236), .CO(w6237) );
	vdp_aoi22 g6120 (.Z(w6239), .B2(w6219), .B1(w6238), .A1(w6235), .A2(w6283) );
	vdp_notif0 g6121 (.A(w6239), .nZ(VRAMA[10]), .nE(w6293) );
	vdp_ha g6122 (.SUM(w6238), .B(w6289), .A(w6237), .CO(w6240) );
	vdp_aoi22 g6123 (.Z(w6241), .B2(w6219), .B1(w6249), .A1(w6238), .A2(w6283) );
	vdp_notif0 g6124 (.A(w6241), .nZ(VRAMA[11]), .nE(w6293) );
	vdp_ha g6125 (.SUM(w6249), .B(w6292), .A(w6240), .CO(w6242) );
	vdp_aoi22 g6126 (.Z(w6244), .B2(w6219), .B1(w6243), .A1(w6249), .A2(w6283) );
	vdp_notif0 g6127 (.A(w6244), .nZ(VRAMA[12]), .nE(w6293) );
	vdp_ha g6128 (.SUM(w6243), .B(w6291), .A(w6242), .CO(w6246) );
	vdp_aoi22 g6129 (.Z(w6247), .B2(w6219), .B1(w6245), .A1(w6243), .A2(w6283) );
	vdp_notif0 g6130 (.A(w6247), .nZ(VRAMA[13]), .nE(w6293) );
	vdp_ha g6131 (.SUM(w6245), .B(w6295), .A(w6246), .CO(w6252) );
	vdp_aoi22 g6132 (.Z(w6250), .B2(w6219), .B1(w6251), .A1(w6245), .A2(w6283) );
	vdp_notif0 g6133 (.A(w6250), .nZ(VRAMA[14]), .nE(w6293) );
	vdp_ha g6134 (.SUM(w6251), .B(w6294), .A(w6252), .CO(w6253) );
	vdp_aoi22 g6135 (.Z(w6256), .B2(w6219), .B1(w6257), .A1(w6251), .A2(w6283) );
	vdp_notif0 g6136 (.A(w6256), .nZ(VRAMA[15]), .nE(w6293) );
	vdp_ha g6137 (.SUM(w6257), .B(w6297), .A(w6253) );
	vdp_aoi22 g6138 (.Z(w6255), .B2(w6219), .B1(w5270), .A1(w6257), .A2(w6283) );
	vdp_notif0 g6139 (.A(w6255), .nZ(VRAMA[16]), .nE(w6293) );
	vdp_not g6140 (.nZ(w6293), .A(w6290) );
	vdp_sr_bit g6141 (.Q(w6290), .D(w6444), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6142 (.nQ(w4539), .D(w6254), .nC(nHCLK2), .C(HCLK2) );
	vdp_and g6143 (.Z(w6444), .B(M5), .A(w22) );
	vdp_or9 g6144 (.Z(w6254), .B(w6152), .A(w6151), .C(w6070), .D(w6081), .F(w6107), .E(w6094), .G(w6120), .H(w6119), .I(w6118) );
	vdp_sr_bit g6145 (.Q(w4612), .D(w6588), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_sr_bit g6146 (.D(w6725), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_fa g6147 (.SUM(w6199), .CO(w6711), .CI(1'b0), .A(w6271), .B(w6200) );
	vdp_fa g6148 (.SUM(w6203), .CO(w6712), .CI(w6711), .A(w6272), .B(w6228) );
	vdp_fa g6149 (.SUM(w6211), .CO(w6713), .CI(w6712), .A(1'b0), .B(w6204) );
	vdp_fa g6150 (.SUM(w6207), .CI(w6713), .A(1'b0), .B(w6209) );
	vdp_notif0 g6151 (.A(1'b1), .nZ(VRAMA[0]), .nE(w6276) );
	vdp_notif0 g6152 (.A(1'b1), .nZ(VRAMA[1]), .nE(w6276) );
	vdp_not g6153 (.nZ(w6208), .A(w6277) );
	vdp_notif0 g6154 (.A(w6208), .nZ(VRAMA[2]), .nE(w6276) );
	vdp_not g6155 (.nZ(w6212), .A(w6279) );
	vdp_notif0 g6156 (.A(w6212), .nZ(VRAMA[3]), .nE(w6276) );
	vdp_not g6157 (.nZ(w6225), .A(w6278) );
	vdp_notif0 g6158 (.A(w6225), .nZ(VRAMA[4]), .nE(w6276) );
	vdp_notif0 g6159 (.A(w6227), .nZ(VRAMA[5]), .nE(w6276) );
	vdp_aoi22 g6160 (.Z(w6227), .B2(w6219), .B1(w6226), .A1(w6269), .A2(w6283) );
	vdp_comp_we g6161 (.nZ(w6219), .A(w1), .Z(w6283) );
	vdp_aon22 g6162 (.Z(w6271), .B2(w6195), .B1(w6269), .A1(w6267), .A2(w6270) );
	vdp_aon22 g6163 (.Z(w6272), .B2(w6195), .B1(w6267), .A1(w6266), .A2(w6270) );
	vdp_comp_we g6164 (.nZ(w6195), .A(w1), .Z(w6270) );
	vdp_or g6165 (.Z(w6725), .B(w6260), .A(w4618) );
	vdp_nor g6166 (.Z(w6588), .B(w6194), .A(w6193) );
	vdp_comp_str g6167 (.nZ(w6323), .A(w6280), .Z(w6296) );
	vdp_slatch g6168 (.D(w6326), .nC(w6323), .C(w6296), .Q(w6151) );
	vdp_aon22 g6169 (.Z(w6327), .B2(w6300), .B1(w6179), .A1(DB[0]), .A2(w6281) );
	vdp_slatch g6170 (.D(w6328), .nC(w6323), .C(w6296), .Q(w6152) );
	vdp_aon22 g6171 (.Z(w6329), .B2(w6300), .B1(w6176), .A1(DB[1]), .A2(w6281) );
	vdp_slatch g6172 (.D(w6330), .nC(w6323), .C(w6296), .Q(w6070) );
	vdp_aon22 g6173 (.Z(w6331), .B2(w6300), .B1(w6173), .A1(DB[2]), .A2(w6281) );
	vdp_slatch g6174 (.D(w6332), .nC(w6323), .C(w6296), .Q(w6081) );
	vdp_aon22 g6175 (.Z(w6333), .B2(w6300), .B1(w6171), .A1(w156), .A2(w6281) );
	vdp_slatch g6176 (.D(w6334), .nC(w6323), .C(w6296), .Q(w6094) );
	vdp_aon22 g6177 (.Z(w6335), .B2(w6300), .B1(w6168), .A1(DB[4]), .A2(w6281) );
	vdp_slatch g6178 (.D(w6336), .nC(w6323), .C(w6296), .Q(w6107) );
	vdp_aon22 g6179 (.Z(w6337), .B2(w6300), .B1(w6165), .A1(DB[5]), .A2(w6281) );
	vdp_slatch g6180 (.D(w6338), .nC(w6323), .C(w6296), .Q(w6120) );
	vdp_aon22 g6181 (.Z(w6339), .B2(w6300), .B1(w6161), .A1(DB[6]), .A2(w6281) );
	vdp_slatch g6182 (.D(w6341), .nC(w6323), .C(w6296), .Q(w6119) );
	vdp_aon22 g6183 (.Z(w6342), .B2(w6300), .B1(w6154), .A1(w160), .A2(w6281) );
	vdp_slatch g6184 (.D(w6340), .nC(w6323), .C(w6296), .Q(w6118) );
	vdp_aon22 g6185 (.Z(w6343), .B2(w6300), .B1(w5112), .A1(DB[8]), .A2(w6281) );
	vdp_slatch g6186 (.D(w6314), .nC(w6311), .C(w6282), .Q(w6286) );
	vdp_aon22 g6187 (.Z(w6350), .B2(w6300), .B1(w6174), .A1(DB[2]), .A2(w6281) );
	vdp_slatch g6188 (.D(w6313), .nC(w6311), .C(w6282), .Q(w6287) );
	vdp_aon22 g6189 (.Z(w6345), .B2(w6300), .B1(w6172), .A1(w156), .A2(w6281) );
	vdp_slatch g6190 (.D(w6320), .nC(w6311), .C(w6282), .Q(w6288) );
	vdp_aon22 g6191 (.Z(w6346), .B2(w6300), .B1(w6169), .A1(DB[4]), .A2(w6281) );
	vdp_slatch g6192 (.D(w6319), .nC(w6311), .C(w6282), .Q(w6289) );
	vdp_aon22 g6193 (.Z(w6349), .B2(w6300), .B1(w6166), .A1(DB[5]), .A2(w6281) );
	vdp_slatch g6194 (.D(w6317), .nC(w6311), .C(w6282), .Q(w6292) );
	vdp_aon22 g6195 (.Z(w6351), .B2(w6300), .B1(w6163), .A1(DB[6]), .A2(w6281) );
	vdp_slatch g6196 (.D(w6318), .nC(w6311), .C(w6282), .Q(w6291) );
	vdp_aon22 g6197 (.Z(w6352), .B2(w6300), .B1(w6158), .A1(w160), .A2(w6281) );
	vdp_slatch g6198 (.D(w6316), .nC(w6311), .C(w6282), .Q(w6295) );
	vdp_aon22 g6199 (.Z(w6353), .B2(w6300), .B1(w5052), .A1(DB[8]), .A2(w6281) );
	vdp_slatch g6200 (.D(w6309), .nC(w6311), .C(w6282), .Q(w6294) );
	vdp_aon22 g6201 (.Z(w6308), .B2(w6300), .B1(w5113), .A1(DB[9]), .A2(w6281) );
	vdp_slatch g6202 (.D(w6324), .nC(w6311), .C(w6282), .Q(w6297) );
	vdp_aon22 g6203 (.Z(w6325), .B2(w6300), .B1(w5121), .A1(DB[10]), .A2(w6281) );
	vdp_slatch g6204 (.D(w6312), .nC(w6311), .C(w6282), .Q(w6284) );
	vdp_aon22 g6205 (.Z(w6347), .B2(w6300), .B1(w6180), .A1(DB[0]), .A2(w6281) );
	vdp_slatch g6206 (.D(w6355), .nC(w6311), .C(w6282), .Q(w6285) );
	vdp_aon22 g6207 (.Z(w6348), .B2(w6300), .B1(w6177), .A1(DB[1]), .A2(w6281) );
	vdp_comp_str g6208 (.nZ(w6311), .A(w6280), .Z(w6282) );
	vdp_not g6209 (.nZ(w6280), .A(w6439) );
	vdp_oai21 g6210 (.Z(w6439), .B(HCLK1), .A1(w6194), .A2(w122) );
	vdp_sr_bit g6211 (.Q(w6440), .D(w6442), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6212 (.Q(w5665), .D(w6441), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6213 (.Q(w6215), .D(w6443), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6214 (.Q(w6344), .D(w5624), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g6215 (.Q(w6263), .D(w6268), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w6260), .CI(w22), .L(w6265), .nL(w6303), .CO(w6304) );
	vdp_cnt_bit_load g6216 (.Q(w6302), .D(w6264), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w6260), .CI(w6304), .L(w6265), .nL(w6303) );
	vdp_comp_we g6217 (.nZ(w6303), .A(w6194), .Z(w6265) );
	vdp_not g6218 (.nZ(w6268), .A(w6305) );
	vdp_not g6219 (.nZ(w6264), .A(w6301) );
	vdp_not g6220 (.nZ(w6261), .A(w125) );
	vdp_nand g6221 (.Z(w6356), .B(w125), .A(w4612) );
	vdp_nand g6222 (.Z(w6262), .B(w6261), .A(w4612) );
	vdp_not g6223 (.nZ(w6300), .A(w6262) );
	vdp_nor g6224 (.Z(w6273), .B(w6302), .A(w6263) );
	vdp_and g6225 (.Z(w6194), .B(w6273), .A(w22) );
	vdp_rs_FF g6226 (.Q(w6442), .R(w6274), .S(w6260) );
	vdp_and3 g6227 (.Z(w6441), .B(w5624), .A(w4619), .C(w6440) );
	vdp_cnt_bit g6228 (.Q(w6443), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w7), .CI(w6344) );
	vdp_not g6229 (.nZ(w6281), .A(w6356) );
	vdp_not g6230 (.nZ(w6307), .A(w4574) );
	vdp_not g6231 (.nZ(w6310), .A(w4575) );
	vdp_comp_str g6232 (.nZ(w6306), .A(w6280), .Z(w6358) );
	vdp_not g6233 (.nZ(w6366), .A(w122) );
	vdp_aon22 g6234 (.Z(w6368), .B2(w6300), .B1(w5172), .A1(DB[0]), .A2(w6281) );
	vdp_slatch g6235 (.D(w6357), .nC(w6306), .C(w6358), .Q(w6146) );
	vdp_bufif0 g6236 (.A(w6365), .Z(DB[0]), .nE(w6366) );
	vdp_aon222 g6237 (.Z(w6365), .B2(w4576), .B1(w6151), .A1(w6146), .A2(w6307), .C1(w6284), .C2(w6310) );
	vdp_aon22 g6238 (.Z(w6371), .B2(w6300), .B1(w5251), .A1(DB[1]), .A2(w6281) );
	vdp_slatch g6239 (.D(w6367), .nC(w6306), .C(w6358), .Q(w6147) );
	vdp_bufif0 g6240 (.A(w6369), .Z(DB[1]), .nE(w6366) );
	vdp_aon222 g6241 (.Z(w6369), .B2(w4576), .B1(w6152), .A1(w6147), .A2(w6307), .C1(w6285), .C2(w6310) );
	vdp_aon22 g6242 (.Z(w6373), .B2(w6300), .B1(w5271), .A1(DB[2]), .A2(w6281) );
	vdp_slatch g6243 (.D(w6370), .nC(w6306), .C(w6358), .Q(w6148) );
	vdp_bufif0 g6244 (.A(w6372), .Z(DB[2]), .nE(w6366) );
	vdp_aon222 g6245 (.Z(w6372), .B2(w4576), .B1(w6070), .A1(w6148), .A2(w6307), .C1(w6286), .C2(w6310) );
	vdp_aon22 g6246 (.Z(w6382), .B2(w6300), .B1(w5236), .A1(w156), .A2(w6281) );
	vdp_slatch g6247 (.D(w6374), .nC(w6306), .C(w6358), .Q(w6153) );
	vdp_bufif0 g6248 (.A(w6381), .Z(w156), .nE(w6366) );
	vdp_aon222 g6249 (.Z(w6381), .B2(w4576), .B1(w6081), .A1(w6153), .A2(w6307), .C1(w6287), .C2(w6310) );
	vdp_aon22 g6250 (.Z(w6379), .B2(w6300), .B1(w4556), .A1(DB[4]), .A2(w6281) );
	vdp_slatch g6251 (.D(w6305), .nC(w6306), .C(w6358), .Q(w6149) );
	vdp_bufif0 g6252 (.A(w6380), .Z(DB[4]), .nE(w6366) );
	vdp_aon222 g6253 (.Z(w6380), .B2(w4576), .B1(w6094), .A1(w6149), .A2(w6307), .C1(w6288), .C2(w6310) );
	vdp_aon22 g6254 (.Z(w6377), .B2(w6300), .B1(w4602), .A1(DB[5]), .A2(w6281) );
	vdp_slatch g6255 (.D(w6301), .nC(w6306), .C(w6358), .Q(w6150) );
	vdp_bufif0 g6256 (.A(w6378), .Z(DB[5]), .nE(w6366) );
	vdp_aon222 g6257 (.Z(w6378), .B2(w4576), .B1(w6107), .A1(w6150), .A2(w6307), .C1(w6289), .C2(w6310) );
	vdp_aon22 g6258 (.Z(w6375), .B2(w6300), .B1(w4557), .A1(DB[6]), .A2(w6281) );
	vdp_slatch g6259 (.D(w6376), .nC(w6306), .C(w6358), .Q(w6196) );
	vdp_bufif0 g6260 (.A(w6398), .Z(DB[6]), .nE(w6366) );
	vdp_aon222 g6261 (.Z(w6398), .B2(w4576), .B1(w6120), .A1(w6196), .A2(w6307), .C1(w6292), .C2(w6310) );
	vdp_aon22 g6262 (.Z(w6394), .B2(w6300), .B1(w4552), .A1(w160), .A2(w6281) );
	vdp_slatch g6263 (.D(w6395), .nC(w6315), .C(w6396), .Q(w6197) );
	vdp_bufif0 g6264 (.A(w6397), .Z(w160), .nE(w6366) );
	vdp_aon222 g6265 (.Z(w6397), .B2(w4576), .B1(w6119), .A1(w6197), .A2(w6307), .C1(w6291), .C2(w6310) );
	vdp_aon22 g6266 (.Z(w6392), .B2(w6300), .B1(w6359), .A1(DB[8]), .A2(w6281) );
	vdp_slatch g6267 (.D(w6393), .nC(w6315), .C(w6396), .Q(w6277) );
	vdp_bufif0 g6268 (.A(w6726), .Z(DB[8]), .nE(w6366) );
	vdp_aon222 g6269 (.Z(w6726), .B2(w4576), .B1(w6118), .A1(w6277), .A2(w6307), .C1(w6295), .C2(w6310) );
	vdp_aon22 g6270 (.Z(w6390), .B2(w6300), .B1(w6364), .A1(DB[9]), .A2(w6281) );
	vdp_slatch g6271 (.D(w6391), .nC(w6315), .C(w6396), .Q(w6279) );
	vdp_bufif0 g6272 (.A(w6399), .Z(DB[9]), .nE(w6366) );
	vdp_aon222 g6273 (.Z(w6399), .B2(w4576), .B1(1'b0), .A1(w6279), .A2(w6307), .C1(w6294), .C2(w6310) );
	vdp_aon22 g6274 (.Z(w6388), .B2(w6300), .B1(w6363), .A1(DB[10]), .A2(w6281) );
	vdp_slatch g6275 (.D(w6389), .nC(w6315), .C(w6396), .Q(w6278) );
	vdp_bufif0 g6276 (.A(w6400), .Z(DB[10]), .nE(w6366) );
	vdp_aon222 g6277 (.Z(w6400), .B2(w4576), .B1(1'b0), .A1(w6278), .A2(w6307), .C1(w6297), .C2(w6310) );
	vdp_aon22 g6278 (.Z(w6386), .B2(w6300), .B1(w6362), .A1(w170), .A2(w6281) );
	vdp_slatch g6279 (.D(w6387), .nC(w6315), .C(w6396), .Q(w6269) );
	vdp_bufif0 g6280 (.A(w6269), .Z(w170), .nE(w6366) );
	vdp_aon22 g6281 (.Z(w6385), .B2(w6300), .B1(w6361), .A1(DB[12]), .A2(w6281) );
	vdp_slatch g6282 (.D(w6401), .nC(w6315), .C(w6396), .Q(w6267) );
	vdp_bufif0 g6283 (.A(w6267), .Z(DB[12]), .nE(w6366) );
	vdp_aon22 g6284 (.Z(w6383), .B2(w6300), .B1(w6360), .A1(DB[13]), .A2(w6281) );
	vdp_slatch g6285 (.D(w6384), .nC(w6315), .C(w6396), .Q(w6266) );
	vdp_bufif0 g6286 (.A(w6266), .Z(DB[13]), .nE(w6366) );
	vdp_comp_str g6287 (.nZ(w6315), .A(w6280), .Z(w6396) );
	vdp_sr_bit g6288 (.Q(w4721), .D(w131), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6289 (.Q(w4722), .D(VRAMA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6290 (.Q(w6409), .D(w6403), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6291 (.Q(w4714), .D(VRAMA[3]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6292 (.Q(w4716), .D(VRAMA[4]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6293 (.Q(w4717), .D(VRAMA[5]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6294 (.Q(w4718), .D(VRAMA[6]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6295 (.Q(w4719), .D(VRAMA[7]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6296 (.Q(w4720), .D(VRAMA[8]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6297 (.Q(w4661), .D(w6407), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6298 (.Q(w4660), .D(w6408), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_and g6299 (.Z(w6407), .B(w134), .A(w5235) );
	vdp_and g6300 (.Z(w6408), .B(w133), .A(w5235) );
	vdp_sr_bit g6301 (.Q(w6423), .D(RD_DATA[0]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6302 (.Q(w6424), .D(RD_DATA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6303 (.Q(w6426), .D(w324), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6304 (.Q(w6425), .D(RD_DATA[2]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_V_PLA g6305 (.o[0](w1892), .o[1](w1893), .o[2](w1894), .o[3](w1895), .o[4](w1896), .o[5](w1897), .o[6](w1898), .o[7](w1899), .o[8](w1900), .o[9](w1901), .o[10](w1902), .o[11](w1903), .o[12](w1904), .o[13](w1905), .o[14](w1906), .o[15](w1907), .o[16](w1908), .o[17](w1909), .o[18](w1910), .o[19](w1911), .o[20](w1913), .o[21](w1912), .o[22](w2025), .o[23](w1915), .o[24](w1992), .o[25](w1916), .o[26](w1917), .o[27](w1993), .o[28](w2007), .o[29](w2006), .o[30](w1914), .o[31](w1919), .o[32](w1891), .o[33](w1890), .o[34](w1889), .o[35](w1920), .o[36](w1935), .o[37](w1936), .o[38](w1888), .o[39](w1887), .o[40](w1938), .o[41](w1887), .o[42](w1937), .o[43](w1885), .o[44](w1884), .o[45](w1883), .o[46](w1882), .o[47](w6733), .Vcnt[0](w1707), .Vcnt[1](w1850), .Vcnt[2](w1948), .Vcnt[3](w1835), .Vcnt[4](w1947), .Vcnt[5](w1791), .Vcnt[6](w1754), .Vcnt[7](w1824), .Vcnt[8](w1851), .ODD_EVEN(ODD/EVEN), .LS0(w1062), .PAL(w1205), .nPAL(w1843), .2(w1842), .3(w1831), .M5(M5) );
	vdp_not g6306 (.A(w594), .nZ(w6731) );
	vdp_not g6307 (.A(w969), .nZ(w6732) );
	vdp_not g6308 (.nZ(w2463), .A(w6731) );
	vdp_not g6309 (.nZ(w2464), .A(w6732) );
	vdp_cram g6310 (.q[8](w2770), .D[8](w2771), .q[7](w2872), .D[7](w2772), .q[6](w2769), .D[6](w2773), .q[5](w2775), .D[5](w2774), .q[4](w2768), .D[4](w2776), .q[3](w2777), .D[3](w3001), .q[2](w2767), .D[2](w2778), .q[1](w2766), .D[1](w2779), .q[0](w2764), .D[0](w2780), .A[0](w2800), .A[1](w2804), .CLK(HCLK1), .A[2](w2810), .A[3](w2819), .A[4](w2840), .A[5](w2839), .B(w2846), .A(w2845) );
	vdp_linebuf_ram g6311 (.q[0](w5358), .D[0](w5758), .q[1](w5347), .D[1](w5757), .q[2](w5335), .D[2](w5756), .q[3](w5324), .D[3](w5769), .q[4](w5768), .D[4](w5743), .q[5](w5736), .D[5](w5742), .q[6](w5748), .D[6](w5770), .q[7](w5357), .D[7](w5755), .q[8](w5348), .D[8](w5754), .q[9](w5334), .D[9](w5753), .q[10](w5325), .D[10](w5729), .q[11](w5730), .D[11](w5728), .q[12](w5749), .D[12](w5733), .q[13](w5750), .D[13](w5767), .q[14](w5356), .D[14](w5758), .q[15](w5349), .D[15](w5757), .q[16](w5333), .D[16](w5756), .q[17](w5326), .D[17](w5759), .q[18](w5731), .D[18](w5764), .q[19](w5735), .D[19](w5760), .q[20](w5762), .D[20](w5761), .q[21](w5355), .D[21](w5755), .q[22](w5350), .D[22](w5754), .q[23](w5332), .D[23](w5753), .q[24](w5327), .D[24](w5746), .q[25](w5732), .D[25](w5744), .q[26](w5734), .D[26](w5752), .q[27](w5763), .D[27](w5751), .CLK(w4537), .A[5](w4531), .A[4](w4532), .A[3](w4533), .A[2](w4534), .A[1](w4535), .A[0](w4536), .A(w5766), .B(w5727), .C(w5726), .D(w5725) );
	vdp_linebuf_ram g6312 (.q[0](w5393), .D[0](w5758), .q[1](w5364), .D[1](w5757), .q[2](w5339), .D[2](w5756), .q[3](w5322), .D[3](w5388), .q[4](w5363), .D[4](w5354), .q[5](w5362), .D[5](w5353), .q[6](w5745), .D[6](w5410), .q[7](w5361), .D[7](w5755), .q[8](w5344), .D[8](w5754), .q[9](w5338), .D[9](w5753), .q[10](w5401), .D[10](w5386), .q[11](w5342), .D[11](w5352), .q[12](w5343), .D[12](w5351), .q[13](w5741), .D[13](w5382), .q[14](w5360), .D[14](w5758), .q[15](w5345), .D[15](w5757), .q[16](w5337), .D[16](w5756), .q[17](w5407), .D[17](w5368), .q[18](w5340), .D[18](w5331), .q[19](w5341), .D[19](w5366), .q[20](w5740), .D[20](w5367), .q[21](w5359), .D[21](w5755), .q[22](w5346), .D[22](w5754), .q[23](w5336), .D[23](w5753), .q[24](w5402), .D[24](w6405), .q[25](w5739), .D[25](w5330), .q[26](w5737), .D[26](w5329), .q[27](w5747), .D[27](w5328), .A[0](w4536), .CLK(w4537), .A[5](w4531), .A[3](w4533), .A[4](w4532), .A[2](w4534), .A[1](w4535), .A(w5453), .B(w5437), .C(w5449), .D(w5439) );
	vdp_att_cashe_ram2 g6313 (.q[0](w4738), .D[0](FIFOo[0]), .q[1](w4737), .D[1](FIFOo[1]), .q[2](w4736), .D[2](FIFOo[2]), .q[3](w4735), .D[3](FIFOo[3]), .q[4](w4711), .D[4](FIFOo[4]), .q[5](w4710), .D[5](w172), .q[6](w4705), .D[6](FIFOo[6]), .q[7](w4879), .D[7](w6423), .q[8](w4917), .D[8](w6424), .q[9](w4902), .D[9](w6425), .q[10](w4899), .D[10](w6426), .CLK(HCLK1), .A[6](w6431), .A[5](w6432), .A[1](w6437), .A[0](w6436), .A[4](w6433), .A[3](w6434), .A[2](w6435), .A(w6428), .B(w4724) );
	vdp_att_cashe_ram1 g6314 (.q[0](w4770), .D[0](FIFOo[0]), .q[1](w4773), .D[1](FIFOo[1]), .q[2](w4766), .D[2](FIFOo[2]), .q[3](w4767), .D[3](FIFOo[3]), .q[4](w4749), .D[4](FIFOo[4]), .q[5](w4741), .D[5](w172), .q[6](w4742), .D[6](FIFOo[6]), .q[7](w4740), .D[7](FIFOo[7]), .q[8](w4739), .D[8](w6423), .q[9](w4734), .D[9](w6424), .CLK(HCLK1), .A[0](w6436), .A[1](w6437), .A[2](w6435), .A[3](w6434), .A[4](w6433), .A[5](w6432), .A[6](w6431), .A(w6430), .B(w6429) );
	vdp_att_temp_ram g6315 (.A[4](w4636), .A[0](w4640), .A[1](w4639), .A[2](w4638), .A[3](w4637), .q[0](w6312), .D[0](w6347), .q[1](w6355), .D[1](w6348), .q[2](w6314), .D[2](w6350), .q[3](w6313), .D[3](w6345), .q[4](w6320), .D[4](w6346), .q[5](w6319), .D[5](w6349), .q[6](w6317), .D[6](w6351), .q[7](w6318), .D[7](w6352), .q[8](w6316), .D[8](w6353), .q[9](w6309), .D[9](w6308), .q[10](w6324), .D[10](w6325), .q[11](w6326), .D[11](w6327), .q[12](w6328), .D[12](w6329), .q[13](w6330), .D[13](w6331), .q[14](w6332), .D[14](w6333), .q[15](w6334), .D[15](w6335), .q[16](w6336), .D[16](w6337), .q[17](w6338), .D[17](w6339), .q[18](w6341), .D[18](w6342), .q[19](w6340), .D[19](w6343), .q[20](w6357), .D[20](w6368), .q[21](w6367), .D[21](w6371), .q[22](w6370), .D[22](w6373), .q[23](w6374), .D[23](w6382), .q[24](w6305), .D[24](w6379), .q[25](w6301), .D[25](w6377), .q[26](w6376), .D[26](w6375), .q[26](w6395), .D[26](w6394), .q[27](w6393), .D[27](w6392), .q[28](w6391), .D[28](w6390), .q[29](w6389), .D[29](w6388), .q[30](w6387), .D[30](w6386), .q[31](w6401), .D[31](w6385), .q[32](w6384), .D[32](w6383), .CLK(HCLK1), .A(w4603), .B(w4604), .C(w4608) );
	vdp_vsram g6316 (.CLK(HCLK1), .D[10](w4024), .q[10](w3982), .D[9](w4028), .q[9](w3975), .D[8](w4026), .q[8](w4001), .D[7](w4025), .q[7](w3967), .D[6](w4013), .q[6](w3963), .D[5](w4011), .q[5](w3955), .D[4](w4018), .q[4](w3951), .D[3](w4020), .q[3](w3948), .D[2](w4023), .q[2](w4006), .D[1](w3981), .q[1](w3943), .D[0](w3999), .q[0](w3938), .A[1](w3756), .A[2](w3728), .A[3](w3727), .A[4](w3726), .A[5](w3725), .A[0](w3757), .A(w3724), .B(w3723) );
	vdp_not g6317 (.nZ(w1825), .A(w6733) );
	vdp_not g6318 (.nZ(w1205), .A(w6734) );
	vdp_H_PLA g6319 (.HPLA[0](w1950), .HPLA[1](w1932), .HPLA[2](w1924), .HPLA[3](w1755), .HPLA[4](w1922), .HPLA[5](w1925), .HPLA[7](w1756), .HPLA[8](w1757), .HPLA[9](w1875), .HPLA[6](w1758), .HPLA[10](w1878), .HPLA[11](w1928), .HPLA[16](w1879), .HPLA[15](w1930), .HPLA[14](w1929), .HPLA[13](w1933), .HPLA[12](w1934), .i0(w59), .HPLA[17](w1778), .HPLA[18](w1777), .HPLA[19](w1877), .HPLA[20](w1876), .HPLA[21](w1926), .HPLA[22](w1921), .Hcnt[0](w1951), .Hcnt[1](w1690), .Hcnt[2](w1695), .Hcnt[3](w1694), .Hcnt[4](w1742), .Hcnt[5](w1775), .Hcnt[6](w1927), .Hcnt[7](w1752), .Hcnt[8](w1780), .H40(H40), .M5(M5), .B(w1779), .C(w1674), .A(w1747), .HPLA[23](w1693), .HPLA[24](w1691), .HPLA[25](w1692), .HPLA[26](w1689), .HPLA[27](w1880), .HPLA[28](w1873), .HPLA[29](w1675), .HPLA[30](w1731), .HPLA[31](w1676), .HPLA[32](w1923), .HPLA[33](w1772), .3(w1931), .HPLA[35](w1808), .HPLA[36](w1770), .HPLA[34](w1952) );
	vdp_slatch g5073 (.D(S[4]), .nC(w5057), .C(w5058), .Q(w5250) );
endmodule // VDP

// Module Definitions [It is possible to wrap here on your primitives]

module vdp_slatch (  nQ, D, C, nC);

	output wire nQ;
	input wire D;
	input wire C;
	input wire nC;

endmodule // vdp_slatch

module vdp_sr_bit (  D, C2, C1, Q, nC2, nC1);

	input wire D;
	input wire C2;
	input wire C1;
	output wire Q;
	input wire nC2;
	input wire nC1;

endmodule // vdp_sr_bit

module vdp_notif0 (  A, nZ, nE);

	input wire A;
	output wire nZ;
	input wire nE;

endmodule // vdp_notif0

module vdp_aon22 (  Z, A1, A2, B1, B2);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire B1;
	input wire B2;

endmodule // vdp_aon22

module vdp_not (  A, nZ);

	input wire A;
	output wire nZ;

endmodule // vdp_not

module vdp_comp_str (  A, Z, nZ);

	input wire A;
	output wire Z;
	output wire nZ;

endmodule // vdp_comp_str

module vdp_comp_we (  A, Z, nZ);

	input wire A;
	output wire Z;
	output wire nZ;

endmodule // vdp_comp_we

module vdp_and (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_and

module vdp_nand (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_nand

module vdp_and3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_and3

module vdp_fa (  SUM, A, B, CO, CI);

	output wire SUM;
	input wire A;
	input wire B;
	output wire CO;
	input wire CI;

endmodule // vdp_fa

module vdp_comp_dff (  D, C2, C1, Q, nC2, nC1);

	input wire D;
	input wire C2;
	input wire C1;
	output wire Q;
	input wire nC2;
	input wire nC1;

endmodule // vdp_comp_dff

module vdp_or (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_or

module vdp_xor (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_xor

module vdp_aoi21 (  Z, B, A1, A2);

	output wire Z;
	input wire B;
	input wire A1;
	input wire A2;

endmodule // vdp_aoi21

module vdp_nor (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_nor

module vdp_and5 (  Z, A, B, C, D, E);

	output wire Z;
	input wire A;
	input wire B;
	input wire C;
	input wire D;
	input wire E;

endmodule // vdp_and5

module vdp_aon2222 (  C2, B2, A2, C1, B1, A1, Z, D2, D1);

	input wire C2;
	input wire B2;
	input wire A2;
	input wire C1;
	input wire B1;
	input wire A1;
	output wire Z;
	input wire D2;
	input wire D1;

endmodule // vdp_aon2222

module vdp_cnt_bit (  R, Q, C1, C2, nC1, nC2, CI);

	input wire R;
	output wire Q;
	input wire C1;
	input wire C2;
	input wire nC1;
	input wire nC2;
	input wire CI;

endmodule // vdp_cnt_bit

module vdp_oai21 (  A1, Z, A2, B);

	input wire A1;
	output wire Z;
	input wire A2;
	input wire B;

endmodule // vdp_oai21

module vdp_comb1 (  Z, A1, B, A2, C);

	output wire Z;
	input wire A1;
	input wire B;
	input wire A2;
	input wire C;

endmodule // vdp_comb1

module vdp_rs_ff (  Q, R, S);

	output wire Q;
	input wire R;
	input wire S;

endmodule // vdp_rs_ff

module vdp_and4 (  A, Z, B, C, D);

	input wire A;
	output wire Z;
	input wire B;
	input wire C;
	input wire D;

endmodule // vdp_and4

module vdp_or3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_or3

module vdp_bufif0 (  A, Z, nE);

	input wire A;
	output wire Z;
	input wire nE;

endmodule // vdp_bufif0

module vdp_aoi221 (  Z, A2, B1, B2, A1, C);

	output wire Z;
	input wire A2;
	input wire B1;
	input wire B2;
	input wire A1;
	input wire C;

endmodule // vdp_aoi221

module vdp_aon33 (  Z, A2, B1, B2, A1, A3, B3);

	output wire Z;
	input wire A2;
	input wire B1;
	input wire B2;
	input wire A1;
	input wire A3;
	input wire B3;

endmodule // vdp_aon33

module vdp_dlatch_inv (  D, C, Q, nC);

	input wire D;
	input wire C;
	output wire Q;
	input wire nC;

endmodule // vdp_dlatch_inv

module vdp_cnt_bit_load (  D, nL, L, R, Q, C1, C2, nC1, nC2, CI, CO);

	input wire D;
	input wire nL;
	input wire L;
	input wire R;
	output wire Q;
	input wire C1;
	input wire C2;
	input wire nC1;
	input wire nC2;
	input wire CI;
	output wire CO;

endmodule // vdp_cnt_bit_load

module vdp_nand3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_nand3

module vdp_nor3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_nor3

module vdp_dff (  Q, R, C, D);

	output wire Q;
	input wire R;
	input wire C;
	input wire D;

endmodule // vdp_dff

module vdp_ha (  SUM, A, B, CO);

	output wire SUM;
	input wire A;
	input wire B;
	output wire CO;

endmodule // vdp_ha

module vdp_slatch_r (  Q, D, R, C, nC);

	output wire Q;
	input wire D;
	input wire R;
	input wire C;
	input wire nC;

endmodule // vdp_slatch_r

module vdp_rs_FF (  nQ, R, S, Q);

	output wire nQ;
	input wire R;
	input wire S;
	output wire Q;

endmodule // vdp_rs_FF

module vdp_or5 (  C, A, B, Z, D, E);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;
	input wire E;

endmodule // vdp_or5

module vdp_2a3oi (  A1, B, Z, A2, C);

	input wire A1;
	input wire B;
	output wire Z;
	input wire A2;
	input wire C;

endmodule // vdp_2a3oi

module vdp_nor5 (  C, A, B, Z, D, E);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;
	input wire E;

endmodule // vdp_nor5

module vdp_or4 (  C, A, B, Z, D);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;

endmodule // vdp_or4

module vdp_aoi22 (  Z, A1, A2, B1, B2);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire B1;
	input wire B2;

endmodule // vdp_aoi22

module vdp_aon222 (  C2, B2, A2, C1, B1, A1, Z);

	input wire C2;
	input wire B2;
	input wire A2;
	input wire C1;
	input wire B1;
	input wire A1;
	output wire Z;

endmodule // vdp_aon222

module vdp_dslatch (  D, C, Q, nC);

	input wire D;
	input wire C;
	output wire Q;
	input wire nC;

endmodule // vdp_dslatch

module vdp_comp_DFF (  D, C2, C1, Q, nC2, nC1);

	input wire D;
	input wire C2;
	input wire C1;
	output wire Q;
	input wire nC2;
	input wire nC1;

endmodule // vdp_comp_DFF

module vdp_nor4 (  C, A, B, Z, D);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;

endmodule // vdp_nor4

module vdp_and6 (  C, A, B, Z, D, E, F);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;
	input wire E;
	input wire F;

endmodule // vdp_and6

module vdp_g1622 (  Z, A);

	output wire Z;
	input wire A;

endmodule // vdp_g1622

module vdp_g1623 (  Z, A);

	output wire Z;
	input wire A;

endmodule // vdp_g1623

module vdp_g1624 (  A, Z);

	input wire A;
	output wire Z;

endmodule // vdp_g1624

module vdp_g1625 (  A, Z);

	input wire A;
	output wire Z;

endmodule // vdp_g1625

module vdp_g1626 (  Z, A);

	output wire Z;
	input wire A;

endmodule // vdp_g1626

module vdp_g1627 (  Z, A);

	output wire Z;
	input wire A;

endmodule // vdp_g1627

module vdp_g1628 (  Z, A);

	output wire Z;
	input wire A;

endmodule // vdp_g1628

module vdp_g1629 (  Z, A);

	output wire Z;
	input wire A;

endmodule // vdp_g1629

module vdp_2?3?I (  Z, A1, A2, C, B);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire C;
	input wire B;

endmodule // vdp_2?3?I

module vdp_RS (  Q, S, R);

	output wire Q;
	input wire S;
	input wire R;

endmodule // vdp_RS

module vdp_TFF (  C2, C1, nC2, nC1, CI, R, A, Q);

	input wire C2;
	input wire C1;
	input wire nC2;
	input wire nC1;
	input wire CI;
	input wire R;
	input wire A;
	output wire Q;

endmodule // vdp_TFF

module vdp_comp_ (  Q, D, nC1, C1, nC2, C2);

	output wire Q;
	input wire D;
	input wire nC1;
	input wire C1;
	input wire nC2;
	input wire C2;

endmodule // vdp_comp_

module vdp_SDELAY8 (  Q, D, nC1, C1, nC2, C2, nC3, C3, nC4, C4, nC5, C5, nC6, C6, nC7, C7, nC8, C8, nC9, C9, nC10, C10, nC11, C11, nC12, C12, nC13, C13, nC14, C14, nC15, C15, nC16, C16);

	output wire Q;
	input wire D;
	input wire nC1;
	input wire C1;
	input wire nC2;
	input wire C2;
	input wire nC3;
	input wire C3;
	input wire nC4;
	input wire C4;
	input wire nC5;
	input wire C5;
	input wire nC6;
	input wire C6;
	input wire nC7;
	input wire C7;
	input wire nC8;
	input wire C8;
	input wire nC9;
	input wire C9;
	input wire nC10;
	input wire C10;
	input wire nC11;
	input wire C11;
	input wire nC12;
	input wire C12;
	input wire nC13;
	input wire C13;
	input wire nC14;
	input wire C14;
	input wire nC15;
	input wire C15;
	input wire nC16;
	input wire C16;

endmodule // vdp_SDELAY8

module vdp_SDELAY7 (  Q, D, C1, nC1, C2, nC2, nC3, C4, nC4, C5, nC5, C6, nC6, C7, nC7, C8, nC8, C9, nC9, C10, nC10, C11, nC11, C12, nC12, C13, nC13, C14, nC14, C3);

	output wire Q;
	input wire D;
	input wire C1;
	input wire nC1;
	input wire C2;
	input wire nC2;
	input wire nC3;
	input wire C4;
	input wire nC4;
	input wire C5;
	input wire nC5;
	input wire C6;
	input wire nC6;
	input wire C7;
	input wire nC7;
	input wire C8;
	input wire nC8;
	input wire C9;
	input wire nC9;
	input wire C10;
	input wire nC10;
	input wire C11;
	input wire nC11;
	input wire C12;
	input wire nC12;
	input wire C13;
	input wire nC13;
	input wire C14;
	input wire nC14;
	input wire C3;

endmodule // vdp_SDELAY7

module vdp_or8 (  Z, A, B, C, D, E, F, G, H);

	output wire Z;
	input wire A;
	input wire B;
	input wire C;
	input wire D;
	input wire E;
	input wire F;
	input wire G;
	input wire H;

endmodule // vdp_or8

module vdp_or7 (  Z, A, B, C, D, E, F, G);

	output wire Z;
	input wire A;
	input wire B;
	input wire C;
	input wire D;
	input wire E;
	input wire F;
	input wire G;

endmodule // vdp_or7

module vdp_dlatch (  Q, C, D, nC);

	output wire Q;
	input wire C;
	input wire D;
	input wire nC;

endmodule // vdp_dlatch

module vdp_clkgen (  PH, CLK1, nCLK1, CLK2, nCLK2);

	input wire PH;
	output wire CLK1;
	output wire nCLK1;
	output wire CLK2;
	output wire nCLK2;

endmodule // vdp_clkgen

module vdp_cgi2a (  Z, A, C, B);

	output wire Z;
	input wire A;
	input wire C;
	input wire B;

endmodule // vdp_cgi2a

module vdp_nand4 (  Z, A, B, D, C);

	output wire Z;
	input wire A;
	input wire B;
	input wire D;
	input wire C;

endmodule // vdp_nand4

module vdp_lfsr_bit (  Q, A, C2, C1, nC2, nC1, C, B);

	output wire Q;
	input wire A;
	input wire C2;
	input wire C1;
	input wire nC2;
	input wire nC1;
	input wire C;
	input wire B;

endmodule // vdp_lfsr_bit

module vdp_aoi222 (  Z, A1, B1, B2, A2, C1, C2);

	output wire Z;
	input wire A1;
	input wire B1;
	input wire B2;
	input wire A2;
	input wire C1;
	input wire C2;

endmodule // vdp_aoi222

module vdp_aon333 (  Z, A1, A2, A3, B1, B2, B3, C1, C2, C3);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire A3;
	input wire B1;
	input wire B2;
	input wire B3;
	input wire C1;
	input wire C2;
	input wire C3;

endmodule // vdp_aon333

module vdp_aoi33 (  Z, A1, A2, A3, B1, B2, B3);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire A3;
	input wire B1;
	input wire B2;
	input wire B3;

endmodule // vdp_aoi33

module vdp_comp_strong (  nZ, Z, A);

	output wire nZ;
	output wire Z;
	input wire A;

endmodule // vdp_comp_strong

module vdp_g2446 (  nZ, A);

	output wire nZ;
	input wire A;

endmodule // vdp_g2446

module vdp_g2447 (  nZ, A);

	output wire nZ;
	input wire A;

endmodule // vdp_g2447

module vdp_g2448 (  nZ, A);

	output wire nZ;
	input wire A;

endmodule // vdp_g2448

module vdp_neg_dff (  Q, C, D, R);

	output wire Q;
	input wire C;
	input wire D;
	input wire R;

endmodule // vdp_neg_dff

module vdp_buf (  Z, A);

	output wire Z;
	input wire A;

endmodule // vdp_buf

module vdp_g2925 (  Z, A, B, C, D);

	output wire Z;
	input wire A;
	input wire B;
	input wire C;
	input wire D;

endmodule // vdp_g2925

module vdp_g2938 (  A, Z);

	input wire A;
	output wire Z;

endmodule // vdp_g2938

module vdp_aon2*8 (  Z, A1, B1, C1, D2, A2, B2, C2, D1, E2, F1, E1, F2, G1, H2, G2, H1);

	output wire Z;
	input wire A1;
	input wire B1;
	input wire C1;
	input wire D2;
	input wire A2;
	input wire B2;
	input wire C2;
	input wire D1;
	input wire E2;
	input wire F1;
	input wire E1;
	input wire F2;
	input wire G1;
	input wire H2;
	input wire G2;
	input wire H1;

endmodule // vdp_aon2*8

module vdp_xnor (  Z, A, B);

	output wire Z;
	input wire A;
	input wire B;

endmodule // vdp_xnor

module vdp_oai211 (  Z, A1, A2, B, C);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire B;
	input wire C;

endmodule // vdp_oai211

module vdp_aoi31 (  Z, B3, B2, B1, A);

	output wire Z;
	input wire B3;
	input wire B2;
	input wire B1;
	input wire A;

endmodule // vdp_aoi31

module vdp_AOI222 (  Z, B1, A1, B2, A2, C1, C2);

	output wire Z;
	input wire B1;
	input wire A1;
	input wire B2;
	input wire A2;
	input wire C1;
	input wire C2;

endmodule // vdp_AOI222

module vdp_SR_bit (  Q, D, C1, C2, nC1, nC2);

	output wire Q;
	input wire D;
	input wire C1;
	input wire C2;
	input wire nC1;
	input wire nC2;

endmodule // vdp_SR_bit

module vdp_cnt_bit_rev (  nC2, nC1, C2, C1, Q, CI, B, A);

	input wire nC2;
	input wire nC1;
	input wire C2;
	input wire C1;
	output wire Q;
	input wire CI;
	input wire B;
	input wire A;

endmodule // vdp_cnt_bit_rev

module vdp_2x_sr_bit (  Q, D, nC2, nC1, C2, C1, nC4, nC3, C4, C3);

	output wire Q;
	input wire D;
	input wire nC2;
	input wire nC1;
	input wire C2;
	input wire C1;
	input wire nC4;
	input wire nC3;
	input wire C4;
	input wire C3;

endmodule // vdp_2x_sr_bit

module vdp_and9 (  Z, B, A, C, D, F, E, G, H, I);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;
	input wire I;

endmodule // vdp_and9

module vdp_nor12 (  Z, B, A, C, D, F, E, G, H, J, I, K, L);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;
	input wire J;
	input wire I;
	input wire K;
	input wire L;

endmodule // vdp_nor12

module vdp_noif0 (  A, nZ, nE);

	input wire A;
	output wire nZ;
	input wire nE;

endmodule // vdp_noif0

module vdp_nor8 (  Z, B, A, C, D, F, E, G, H);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;

endmodule // vdp_nor8

module vdp_aon21_sr (  Q, A1, A2, B, nC2, nC1, C2, C1);

	output wire Q;
	input wire A1;
	input wire A2;
	input wire B;
	input wire nC2;
	input wire nC1;
	input wire C2;
	input wire C1;

endmodule // vdp_aon21_sr

module vdp_or9 (  Z, B, A, C, D, F, E, G, H, I);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;
	input wire I;

endmodule // vdp_or9

module vdp_V_PLA (  o[0], o[1], o[2], o[3], o[4], o[5], o[6], o[7], o[8], o[9], o[10], o[11], o[12], o[13], o[14], o[15], o[16], o[17], o[18], o[19], o[20], o[21], o[22], o[23], o[24], o[25], o[26], o[27], o[28], o[29], o[30], o[31], o[32], o[33], o[34], o[35], o[36], o[37], o[38], o[39], o[40], o[41], o[42], o[43], o[44], o[45], o[46], o[47], Vcnt[0], Vcnt[1], Vcnt[2], Vcnt[3], Vcnt[4], Vcnt[5], Vcnt[6], Vcnt[7], Vcnt[8], ODD_EVEN, LS0, PAL, nPAL, 2, 3, M5);

	output wire o[0];
	output wire o[1];
	output wire o[2];
	output wire o[3];
	output wire o[4];
	output wire o[5];
	output wire o[6];
	output wire o[7];
	output wire o[8];
	output wire o[9];
	output wire o[10];
	output wire o[11];
	output wire o[12];
	output wire o[13];
	output wire o[14];
	output wire o[15];
	output wire o[16];
	output wire o[17];
	output wire o[18];
	output wire o[19];
	output wire o[20];
	output wire o[21];
	output wire o[22];
	output wire o[23];
	output wire o[24];
	output wire o[25];
	output wire o[26];
	output wire o[27];
	output wire o[28];
	output wire o[29];
	output wire o[30];
	output wire o[31];
	output wire o[32];
	output wire o[33];
	output wire o[34];
	output wire o[35];
	output wire o[36];
	output wire o[37];
	output wire o[38];
	output wire o[39];
	output wire o[40];
	output wire o[41];
	output wire o[42];
	output wire o[43];
	output wire o[44];
	output wire o[45];
	output wire o[46];
	output wire o[47];
	input wire Vcnt[0];
	input wire Vcnt[1];
	input wire Vcnt[2];
	input wire Vcnt[3];
	input wire Vcnt[4];
	input wire Vcnt[5];
	input wire Vcnt[6];
	input wire Vcnt[7];
	input wire Vcnt[8];
	input wire ODD_EVEN;
	input wire LS0;
	input wire PAL;
	input wire nPAL;
	input wire 2;
	input wire 3;
	input wire M5;

endmodule // vdp_V_PLA

module vdp_cram (  q[8], D[8], q[7], D[7], q[6], D[6], q[5], D[5], q[4], D[4], q[3], D[3], q[2], D[2], q[1], D[1], q[0], D[0], A[0], A[1], CLK, A[2], A[3], A[4], A[5], B, A);

	output wire q[8];
	input wire D[8];
	output wire q[7];
	input wire D[7];
	output wire q[6];
	input wire D[6];
	output wire q[5];
	input wire D[5];
	output wire q[4];
	input wire D[4];
	output wire q[3];
	input wire D[3];
	output wire q[2];
	input wire D[2];
	output wire q[1];
	input wire D[1];
	output wire q[0];
	input wire D[0];
	input wire A[0];
	input wire A[1];
	input wire CLK;
	input wire A[2];
	input wire A[3];
	input wire A[4];
	input wire A[5];
	input wire B;
	input wire A;

endmodule // vdp_cram

module vdp_linebuf_ram (  q[0], D[0], q[1], D[1], q[2], D[2], q[3], D[3], q[4], D[4], q[5], D[5], q[6], D[6], q[7], D[7], q[8], D[8], q[9], D[9], q[10], D[10], q[11], D[11], q[12], D[12], q[13], D[13], q[14], D[14], q[15], D[15], q[16], D[16], q[17], D[17], q[18], D[18], q[19], D[19], q[20], D[20], q[21], D[21], q[22], D[22], q[23], D[23], q[24], D[24], q[25], D[25], q[26], D[26], q[27], D[27], CLK, A[5], A[4], A[3], A[2], A[1], A[0], A, B, C, D);

	output wire q[0];
	input wire D[0];
	output wire q[1];
	input wire D[1];
	output wire q[2];
	input wire D[2];
	output wire q[3];
	input wire D[3];
	output wire q[4];
	input wire D[4];
	output wire q[5];
	input wire D[5];
	output wire q[6];
	input wire D[6];
	output wire q[7];
	input wire D[7];
	output wire q[8];
	input wire D[8];
	output wire q[9];
	input wire D[9];
	output wire q[10];
	input wire D[10];
	output wire q[11];
	input wire D[11];
	output wire q[12];
	input wire D[12];
	output wire q[13];
	input wire D[13];
	output wire q[14];
	input wire D[14];
	output wire q[15];
	input wire D[15];
	output wire q[16];
	input wire D[16];
	output wire q[17];
	input wire D[17];
	output wire q[18];
	input wire D[18];
	output wire q[19];
	input wire D[19];
	output wire q[20];
	input wire D[20];
	output wire q[21];
	input wire D[21];
	output wire q[22];
	input wire D[22];
	output wire q[23];
	input wire D[23];
	output wire q[24];
	input wire D[24];
	output wire q[25];
	input wire D[25];
	output wire q[26];
	input wire D[26];
	output wire q[27];
	input wire D[27];
	input wire CLK;
	input wire A[5];
	input wire A[4];
	input wire A[3];
	input wire A[2];
	input wire A[1];
	input wire A[0];
	input wire A;
	input wire B;
	input wire C;
	input wire D;

endmodule // vdp_linebuf_ram

module vdp_att_cashe_ram2 (  q[0], D[0], q[1], D[1], q[2], D[2], q[3], D[3], q[4], D[4], q[5], D[5], q[6], D[6], q[7], D[7], q[8], D[8], q[9], D[9], q[10], D[10], CLK, A[6], A[5], A[1], A[0], A[4], A[3], A[2], A, B);

	output wire q[0];
	input wire D[0];
	output wire q[1];
	input wire D[1];
	output wire q[2];
	input wire D[2];
	output wire q[3];
	input wire D[3];
	output wire q[4];
	input wire D[4];
	output wire q[5];
	input wire D[5];
	output wire q[6];
	input wire D[6];
	output wire q[7];
	input wire D[7];
	output wire q[8];
	input wire D[8];
	output wire q[9];
	input wire D[9];
	output wire q[10];
	input wire D[10];
	input wire CLK;
	input wire A[6];
	input wire A[5];
	input wire A[1];
	input wire A[0];
	input wire A[4];
	input wire A[3];
	input wire A[2];
	input wire A;
	input wire B;

endmodule // vdp_att_cashe_ram2

module vdp_att_cashe_ram1 (  q[0], D[0], q[1], D[1], q[2], D[2], q[3], D[3], q[4], D[4], q[5], D[5], q[6], D[6], q[7], D[7], q[8], D[8], q[9], D[9], CLK, A[0], A[1], A[2], A[3], A[4], A[5], A[6], A, B);

	output wire q[0];
	input wire D[0];
	output wire q[1];
	input wire D[1];
	output wire q[2];
	input wire D[2];
	output wire q[3];
	input wire D[3];
	output wire q[4];
	input wire D[4];
	output wire q[5];
	input wire D[5];
	output wire q[6];
	input wire D[6];
	output wire q[7];
	input wire D[7];
	output wire q[8];
	input wire D[8];
	output wire q[9];
	input wire D[9];
	input wire CLK;
	input wire A[0];
	input wire A[1];
	input wire A[2];
	input wire A[3];
	input wire A[4];
	input wire A[5];
	input wire A[6];
	input wire A;
	input wire B;

endmodule // vdp_att_cashe_ram1

module vdp_att_temp_ram (  A[4], A[0], A[1], A[2], A[3], q[0], D[0], q[1], D[1], q[2], D[2], q[3], D[3], q[4], D[4], q[5], D[5], q[6], D[6], q[7], D[7], q[8], D[8], q[9], D[9], q[10], D[10], q[11], D[11], q[12], D[12], q[13], D[13], q[14], D[14], q[15], D[15], q[16], D[16], q[17], D[17], q[18], D[18], q[19], D[19], q[20], D[20], q[21], D[21], q[22], D[22], q[23], D[23], q[24], D[24], q[25], D[25], q[26], D[26], q[26], D[26], q[27], D[27], q[28], D[28], q[29], D[29], q[30], D[30], q[31], D[31], q[32], D[32], CLK, A, B, C);

	input wire A[4];
	input wire A[0];
	input wire A[1];
	input wire A[2];
	input wire A[3];
	output wire q[0];
	input wire D[0];
	output wire q[1];
	input wire D[1];
	output wire q[2];
	input wire D[2];
	output wire q[3];
	input wire D[3];
	output wire q[4];
	input wire D[4];
	output wire q[5];
	input wire D[5];
	output wire q[6];
	input wire D[6];
	output wire q[7];
	input wire D[7];
	output wire q[8];
	input wire D[8];
	output wire q[9];
	input wire D[9];
	output wire q[10];
	input wire D[10];
	output wire q[11];
	input wire D[11];
	output wire q[12];
	input wire D[12];
	output wire q[13];
	input wire D[13];
	output wire q[14];
	input wire D[14];
	output wire q[15];
	input wire D[15];
	output wire q[16];
	input wire D[16];
	output wire q[17];
	input wire D[17];
	output wire q[18];
	input wire D[18];
	output wire q[19];
	input wire D[19];
	output wire q[20];
	input wire D[20];
	output wire q[21];
	input wire D[21];
	output wire q[22];
	input wire D[22];
	output wire q[23];
	input wire D[23];
	output wire q[24];
	input wire D[24];
	output wire q[25];
	input wire D[25];
	output wire q[26];
	input wire D[26];
	output wire q[26];
	input wire D[26];
	output wire q[27];
	input wire D[27];
	output wire q[28];
	input wire D[28];
	output wire q[29];
	input wire D[29];
	output wire q[30];
	input wire D[30];
	output wire q[31];
	input wire D[31];
	output wire q[32];
	input wire D[32];
	input wire CLK;
	input wire A;
	input wire B;
	input wire C;

endmodule // vdp_att_temp_ram

module vdp_vsram (  CLK, D[10], q[10], D[9], q[9], D[8], q[8], D[7], q[7], D[6], q[6], D[5], q[5], D[4], q[4], D[3], q[3], D[2], q[2], D[1], q[1], D[0], q[0], A[1], A[2], A[3], A[4], A[5], A[0], A, B);

	input wire CLK;
	input wire D[10];
	output wire q[10];
	input wire D[9];
	output wire q[9];
	input wire D[8];
	output wire q[8];
	input wire D[7];
	output wire q[7];
	input wire D[6];
	output wire q[6];
	input wire D[5];
	output wire q[5];
	input wire D[4];
	output wire q[4];
	input wire D[3];
	output wire q[3];
	input wire D[2];
	output wire q[2];
	input wire D[1];
	output wire q[1];
	input wire D[0];
	output wire q[0];
	input wire A[1];
	input wire A[2];
	input wire A[3];
	input wire A[4];
	input wire A[5];
	input wire A[0];
	input wire A;
	input wire B;

endmodule // vdp_vsram

module vdp_H_PLA (  HPLA[0], HPLA[1], HPLA[2], HPLA[3], HPLA[4], HPLA[5], HPLA[7], HPLA[8], HPLA[9], HPLA[6], HPLA[10], HPLA[11], HPLA[16], HPLA[15], HPLA[14], HPLA[13], HPLA[12], i0, HPLA[17], HPLA[18], HPLA[19], HPLA[20], HPLA[21], HPLA[22], Hcnt[0], Hcnt[1], Hcnt[2], Hcnt[3], Hcnt[4], Hcnt[5], Hcnt[6], Hcnt[7], Hcnt[8], H40, M5, B, C, A, HPLA[23], HPLA[24], HPLA[25], HPLA[26], HPLA[27], HPLA[28], HPLA[29], HPLA[30], HPLA[31], HPLA[32], HPLA[33], 3, HPLA[35], HPLA[36], HPLA[34]);

	output wire HPLA[0];
	output wire HPLA[1];
	output wire HPLA[2];
	output wire HPLA[3];
	output wire HPLA[4];
	output wire HPLA[5];
	output wire HPLA[7];
	output wire HPLA[8];
	output wire HPLA[9];
	output wire HPLA[6];
	output wire HPLA[10];
	output wire HPLA[11];
	output wire HPLA[16];
	output wire HPLA[15];
	output wire HPLA[14];
	output wire HPLA[13];
	output wire HPLA[12];
	input wire i0;
	output wire HPLA[17];
	output wire HPLA[18];
	output wire HPLA[19];
	output wire HPLA[20];
	output wire HPLA[21];
	output wire HPLA[22];
	input wire Hcnt[0];
	input wire Hcnt[1];
	input wire Hcnt[2];
	input wire Hcnt[3];
	input wire Hcnt[4];
	input wire Hcnt[5];
	input wire Hcnt[6];
	input wire Hcnt[7];
	input wire Hcnt[8];
	input wire H40;
	input wire M5;
	input wire B;
	input wire C;
	input wire A;
	output wire HPLA[23];
	output wire HPLA[24];
	output wire HPLA[25];
	output wire HPLA[26];
	output wire HPLA[27];
	output wire HPLA[28];
	output wire HPLA[29];
	output wire HPLA[30];
	output wire HPLA[31];
	output wire HPLA[32];
	output wire HPLA[33];
	input wire 3;
	output wire HPLA[35];
	output wire HPLA[36];
	output wire HPLA[34];

endmodule // vdp_H_PLA



// ERROR: conflicting wire VRAMA[8]
// WARNING: wire not driving anything w128
// ERROR: conflicting wire AD_DATA[7]
// ERROR: conflicting wire AD_DATA[6]
// ERROR: conflicting wire AD_DATA[4]
// ERROR: conflicting wire RD_DATA[2]
// ERROR: conflicting wire RD_DATA[1]
// ERROR: conflicting wire RD_DATA[0]
// ERROR: conflicting wire AD_DATA[5]
// ERROR: conflicting wire DB[0]
// ERROR: conflicting wire DB[1]
// ERROR: conflicting wire DB[2]
// ERROR: conflicting wire w156
// ERROR: conflicting wire DB[4]
// ERROR: conflicting wire DB[5]
// ERROR: conflicting wire DB[6]
// ERROR: conflicting wire w160
// ERROR: conflicting wire DB[8]
// ERROR: conflicting wire DB[9]
// ERROR: conflicting wire AD_DATA[3]
// ERROR: conflicting wire AD_DATA[2]
// ERROR: conflicting wire AD_DATA[1]
// ERROR: conflicting wire AD_DATA[0]
// ERROR: conflicting wire DB[14]
// ERROR: conflicting wire DB[13]
// ERROR: conflicting wire DB[12]
// ERROR: conflicting wire w170
// ERROR: conflicting wire DB[10]
// ERROR: floating wire w172
// ERROR: floating wire w190
// ERROR: conflicting wire RD_DATA[4]
// ERROR: floating wire w221
// ERROR: conflicting wire RD_DATA[6]
// ERROR: floating wire w237
// ERROR: conflicting wire w239
// ERROR: conflicting wire w247
// ERROR: conflicting wire w256
// ERROR: conflicting wire w264
// ERROR: conflicting wire w281
// ERROR: conflicting wire w290
// ERROR: conflicting wire w291
// ERROR: conflicting wire w300
// ERROR: conflicting wire w308
// ERROR: conflicting wire w324
// ERROR: conflicting wire w325
// ERROR: floating wire w338
// ERROR: conflicting wire RD_DATA[5]
// ERROR: floating wire w354
// ERROR: conflicting wire w358
// ERROR: conflicting wire w359
// ERROR: floating wire w462
// ERROR: conflicting wire VRAMA[0]
// ERROR: floating wire w578
// ERROR: conflicting wire VRAMA[7]
// ERROR: conflicting wire VRAMA[9]
// ERROR: conflicting wire VRAMA[10]
// ERROR: conflicting wire VRAMA[6]
// ERROR: conflicting wire VRAMA[5]
// ERROR: conflicting wire VRAMA[11]
// ERROR: conflicting wire VRAMA[12]
// ERROR: conflicting wire VRAMA[4]
// ERROR: conflicting wire VRAMA[13]
// ERROR: conflicting wire VRAMA[3]
// ERROR: conflicting wire VRAMA[14]
// ERROR: conflicting wire VRAMA[2]
// ERROR: conflicting wire CA[14]
// ERROR: conflicting wire VRAMA[15]
// ERROR: conflicting wire VRAMA[1]
// ERROR: conflicting wire VRAMA[16]
// ERROR: floating wire w801
// ERROR: floating wire w803
// ERROR: floating wire w816
// ERROR: floating wire w817
// ERROR: floating wire w834
// ERROR: floating wire w930
// ERROR: floating wire w932
// ERROR: floating wire w1001
// ERROR: floating wire w1078
// ERROR: floating wire w1084
// ERROR: conflicting wire COL[0]
// ERROR: conflicting wire COL[1]
// ERROR: conflicting wire COL[2]
// ERROR: conflicting wire COL[3]
// ERROR: conflicting wire COL[4]
// ERROR: conflicting wire COL[5]
// ERROR: conflicting wire COL[6]
// ERROR: floating wire w1101
// ERROR: floating wire w1102
// ERROR: floating wire w1190
// ERROR: floating wire w1211
// ERROR: floating wire w1230
// ERROR: floating wire w1304
// ERROR: floating wire w1311
// ERROR: floating wire w1319
// ERROR: floating wire w1336
// ERROR: floating wire w1367
// ERROR: floating wire w1391
// ERROR: floating wire w1516
// ERROR: floating wire w1611
// ERROR: floating wire w1688
// ERROR: floating wire w1698
// ERROR: floating wire w1709
// ERROR: floating wire w1727
// ERROR: floating wire w1749
// WARNING: wire not driving anything w1777
// ERROR: floating wire w1793
// ERROR: conflicting wire w1798
// ERROR: floating wire w1834
// ERROR: floating wire w1844
// ERROR: conflicting wire w1887
// WARNING: wire not driving anything w1917
// ERROR: floating wire w1918
// ERROR: floating wire w1941
// ERROR: floating wire w1953
// ERROR: floating wire w1996
// ERROR: floating wire w2085
// ERROR: floating wire w2170
// ERROR: floating wire w2271
// ERROR: floating wire w2306
// ERROR: floating wire w2496
// ERROR: floating wire w2575
// ERROR: floating wire w2645
// ERROR: floating wire w2651
// ERROR: floating wire w2719
// WARNING: wire not driving anything w2734
// ERROR: floating wire w2816
// ERROR: floating wire w3070
// ERROR: floating wire w3137
// ERROR: floating wire w3143
// ERROR: floating wire w3225
// ERROR: floating wire w3335
// WARNING: wire not driving anything w3344
// ERROR: floating wire w3387
// WARNING: wire not driving anything w3396
// ERROR: floating wire w3480
// ERROR: floating wire w3550
// ERROR: conflicting wire w3557
// ERROR: floating wire w3630
// ERROR: floating wire w3687
// ERROR: floating wire w3697
// ERROR: floating wire w3698
// ERROR: floating wire w3730
// ERROR: floating wire w3773
// ERROR: floating wire w3778
// ERROR: floating wire w3832
// ERROR: floating wire w3834
// ERROR: floating wire w3910
// ERROR: floating wire w3936
// ERROR: floating wire w3991
// ERROR: floating wire w4110
// ERROR: floating wire w4443
// ERROR: floating wire w4455
// ERROR: floating wire w4528
// ERROR: floating wire w4613
// ERROR: floating wire w4682
// ERROR: floating wire w4687
// ERROR: floating wire w4725
// ERROR: floating wire w4728
// ERROR: floating wire w4783
// ERROR: floating wire w4788
// ERROR: floating wire w4817
// ERROR: floating wire w4861
// ERROR: floating wire w4919
// ERROR: floating wire w4934
// ERROR: floating wire w4941
// ERROR: floating wire w4943
// ERROR: floating wire w4982
// ERROR: floating wire w5175
// ERROR: floating wire w5232
// ERROR: floating wire w5370
// ERROR: floating wire w5385
// ERROR: floating wire w5389
// ERROR: floating wire w5397
// ERROR: floating wire w5427
// ERROR: floating wire w5477
// ERROR: floating wire w5486
// ERROR: floating wire w5492
// ERROR: floating wire w5518
// ERROR: floating wire w5549
// WARNING: wire not driving anything w5563
// ERROR: conflicting wire w5590
// ERROR: floating wire w5598
// ERROR: floating wire w5670
// ERROR: floating wire w5682
// ERROR: floating wire w5699
// ERROR: floating wire w5738
// ERROR: floating wire w5792
// ERROR: floating wire w5856
// ERROR: conflicting wire w5876
// ERROR: floating wire w5937
// ERROR: floating wire w5939
// ERROR: floating wire w5952
// ERROR: conflicting wire w5961
// ERROR: floating wire w5990
// ERROR: floating wire w6021
// ERROR: floating wire w6038
// ERROR: floating wire w6182
// ERROR: floating wire w6198
// ERROR: floating wire w6229
// ERROR: floating wire w6275
// ERROR: floating wire w6321
// ERROR: floating wire w6322
// ERROR: conflicting wire w6411
// ERROR: floating wire w6630
// ERROR: floating wire w6745
// ERROR: floating wire w6747
// ERROR: floating wire w6748
// WARNING: Cell vdp_fa:g385 port CO not connected.
// WARNING: Cell vdp_and:g527 port Z not connected.
// WARNING: Cell vdp_cnt_bit_load:g871 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g873 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g1405 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g1406 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1407 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1408 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1409 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1410 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1411 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1412 port Q not connected.
// WARNING: Cell vdp_or:g1576 port Z not connected.
// WARNING: Cell vdp_cnt_bit_load:g1959 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g1960 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2145 port CO not connected.
// WARNING: Cell vdp_ha:g2278 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2280 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2282 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2284 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2286 port CO not connected.
// WARNING: Cell vdp_rs_ff:g2380 port nQ not connected.
// WARNING: Cell vdp_rs_ff:g2381 port nQ not connected.
// WARNING: Cell vdp_comp_we:g2612 port nZ not connected.
// WARNING: Cell vdp_fa:g3842 port CO not connected.
// WARNING: Cell vdp_fa:g4058 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g4437 port CO not connected.
// WARNING: Cell vdp_fa:g4453 port CO not connected.
// WARNING: Cell vdp_fa:g4463 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g5851 port CO not connected.
// WARNING: Cell vdp_fa:g5862 port CO not connected.
// WARNING: Cell vdp_fa:g5888 port CO not connected.
// WARNING: Cell vdp_fa:g5892 port CO not connected.
// WARNING: Cell vdp_fa:g6086 port CO not connected.
// WARNING: Cell vdp_ha:g6137 port CO not connected.
// WARNING: Cell vdp_sr_bit:g6146 port Q not connected.
// WARNING: Cell vdp_fa:g6150 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g6216 port CO not connected.
