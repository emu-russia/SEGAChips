// TOP описание процессора Z80 сэги

module Z80 ();

endmodule // Z80
