module VDP (  CH0_EN, CH0VOL[0], CH0VOL[1], CH1_EN, CH1VOL[0], CH1VOL[1], CH2_EN, CH2VOL[0], CH2VOL[1], CH3_EN, CH3VOL[0], CH3VOL[1], PSGDAC0[0], PSGDAC0[1], PSGDAC0[2], PSGDAC0[3], PSGDAC0[4], PSGDAC0[5], PSGDAC0[6], PSGDAC0[7], PSGDAC1[0], PSGDAC1[1], PSGDAC1[2], PSGDAC1[3], PSGDAC1[4], PSGDAC1[5], PSGDAC1[6], PSGDAC1[7], PSGDAC2[0], PSGDAC2[1], PSGDAC2[2], PSGDAC2[3], PSGDAC2[4], PSGDAC2[5], PSGDAC2[6], PSGDAC2[7], PSGDAC3[0], PSGDAC3[1], PSGDAC3[2], PSGDAC3[3], PSGDAC3[4], PSGDAC3[5], PSGDAC3[6], PSGDAC3[7], CAi[22], CAo[22], CA[19], DTACK_OUT, Z80_INT, RA[7], RA[6], RA[5], RA[4], RA[2], RA[1], RA[0], nRAS0, RA[3], nCAS0, nOE0, nLWR, nUWR, DTACK_IN, RnW, nLDS, nUDS, nAS, nM1, nWR, nRD, nIORQ, nILP2, nILP1, nINTAK, nMREQ, nBG, BGACK_OUT, BGACK_IN, nBR, VSYNC, nCSYNC, nCSYNC_IN, nHSYNC, nHSYNC_IN, DB[15], DB[14], DB[13], DB[12], DB[11], DB[10], DB[9], DB[8], DB[7], DB[6], DB[5], DB[4], DB[3], DB[2], DB[1], DB[0], CA[0], CA[1], CA[2], CA[3], CA[4], CA[5], CA[6], CA[7], CA[8], CA[9], CA[10], CA[11], CA[12], CA[13], CA[14], CA[15], CA[16], CA[17], CA[18], CA[20], CA[21], R_DAC[0], R_DAC[1], R_DAC[2], R_DAC[3], R_DAC[4], R_DAC[5], R_DAC[6], R_DAC[7], R_DAC[8], G_DAC[0], G_DAC[1], G_DAC[2], G_DAC[3], G_DAC[4], G_DAC[5], G_DAC[6], G_DAC[7], G_DAC[8], R_DAC[9], R_DAC[10], R_DAC[11], R_DAC[12], R_DAC[13], R_DAC[14], R_DAC[15], R_DAC[16], B_DAC[0], B_DAC[1], B_DAC[2], B_DAC[3], B_DAC[4], B_DAC[5], B_DAC[6], B_DAC[7], B_DAC[8], G_DAC[9], G_DAC[10], G_DAC[11], G_DAC[12], G_DAC[13], G_DAC[14], G_DAC[15], G_DAC[16], B_DAC[9], B_DAC[10], B_DAC[11], B_DAC[12], B_DAC[13], B_DAC[14], B_DAC[15], B_DAC[16], nOE1, nWE0, nWE1, nCAS1, nRAS1, AD_RD_DIR, nYS, nSC, nSE0_1, ADo[7], ADo[6], ADo[5], ADo[4], ADo[3], ADo[2], ADo[1], ADo[0], RDo[6], RDo[5], RDo[4], RDo[3], RDo[2], RDo[1], RDo[0], RDi[6], RDi[7], RDi[4], RDi[5], RDi[2], RDi[3], RDi[0], RDi[1], ADi[6], ADi[7], ADi[4], ADi[5], ADi[2], ADi[3], ADi[0], ADi[1], RDo[7], SD[7], SD[6], SD[5], SD[4], SD[3], SD[2], SD[1], SD[0], CLK1, CLK0, EDCLKi, EDCLKo, MCLK, SUB_CLK, nRES_PAD, 68kCLKi, EDCLKd, CA_PAD_DIR, DB_PAD_DIR, SEL0_M3, nPAL, nHL, SPA/Bo, SPA/Bi);

	output wire CH0_EN;
	output wire CH0VOL[0];
	output wire CH0VOL[1];
	output wire CH1_EN;
	output wire CH1VOL[0];
	output wire CH1VOL[1];
	output wire CH2_EN;
	output wire CH2VOL[0];
	output wire CH2VOL[1];
	output wire CH3_EN;
	output wire CH3VOL[0];
	output wire CH3VOL[1];
	output wire PSGDAC0[0];
	output wire PSGDAC0[1];
	output wire PSGDAC0[2];
	output wire PSGDAC0[3];
	output wire PSGDAC0[4];
	output wire PSGDAC0[5];
	output wire PSGDAC0[6];
	output wire PSGDAC0[7];
	output wire PSGDAC1[0];
	output wire PSGDAC1[1];
	output wire PSGDAC1[2];
	output wire PSGDAC1[3];
	output wire PSGDAC1[4];
	output wire PSGDAC1[5];
	output wire PSGDAC1[6];
	output wire PSGDAC1[7];
	output wire PSGDAC2[0];
	output wire PSGDAC2[1];
	output wire PSGDAC2[2];
	output wire PSGDAC2[3];
	output wire PSGDAC2[4];
	output wire PSGDAC2[5];
	output wire PSGDAC2[6];
	output wire PSGDAC2[7];
	output wire PSGDAC3[0];
	output wire PSGDAC3[1];
	output wire PSGDAC3[2];
	output wire PSGDAC3[3];
	output wire PSGDAC3[4];
	output wire PSGDAC3[5];
	output wire PSGDAC3[6];
	output wire PSGDAC3[7];
	input wire CAi[22];
	output wire CAo[22];
	output wire CA[19];
	output wire DTACK_OUT;
	output wire Z80_INT;
	output wire RA[7];
	output wire RA[6];
	output wire RA[5];
	output wire RA[4];
	output wire RA[2];
	output wire RA[1];
	output wire RA[0];
	output wire nRAS0;
	output wire RA[3];
	output wire nCAS0;
	output wire nOE0;
	output wire nLWR;
	output wire nUWR;
	input wire DTACK_IN;
	input wire RnW;
	input wire nLDS;
	input wire nUDS;
	input wire nAS;
	input wire nM1;
	input wire nWR;
	input wire nRD;
	input wire nIORQ;
	output wire nILP2;
	output wire nILP1;
	input wire nINTAK;
	input wire nMREQ;
	input wire nBG;
	output wire BGACK_OUT;
	input wire BGACK_IN;
	output wire nBR;
	output wire VSYNC;
	output wire nCSYNC;
	input wire nCSYNC_IN;
	output wire nHSYNC;
	input wire nHSYNC_IN;
	inout wire DB[15];
	inout wire DB[14];
	inout wire DB[13];
	inout wire DB[12];
	inout wire DB[11];
	inout wire DB[10];
	inout wire DB[9];
	inout wire DB[8];
	inout wire DB[7];
	inout wire DB[6];
	inout wire DB[5];
	inout wire DB[4];
	inout wire DB[3];
	inout wire DB[2];
	inout wire DB[1];
	inout wire DB[0];
	inout wire CA[0];
	inout wire CA[1];
	inout wire CA[2];
	inout wire CA[3];
	inout wire CA[4];
	inout wire CA[5];
	inout wire CA[6];
	inout wire CA[7];
	inout wire CA[8];
	inout wire CA[9];
	inout wire CA[10];
	inout wire CA[11];
	inout wire CA[12];
	inout wire CA[13];
	inout wire CA[14];
	inout wire CA[15];
	inout wire CA[16];
	inout wire CA[17];
	output wire CA[18];
	inout wire CA[20];
	inout wire CA[21];
	output wire R_DAC[0];
	output wire R_DAC[1];
	output wire R_DAC[2];
	output wire R_DAC[3];
	output wire R_DAC[4];
	output wire R_DAC[5];
	output wire R_DAC[6];
	output wire R_DAC[7];
	output wire R_DAC[8];
	output wire G_DAC[0];
	output wire G_DAC[1];
	output wire G_DAC[2];
	output wire G_DAC[3];
	output wire G_DAC[4];
	output wire G_DAC[5];
	output wire G_DAC[6];
	output wire G_DAC[7];
	output wire G_DAC[8];
	output wire R_DAC[9];
	output wire R_DAC[10];
	output wire R_DAC[11];
	output wire R_DAC[12];
	output wire R_DAC[13];
	output wire R_DAC[14];
	output wire R_DAC[15];
	output wire R_DAC[16];
	output wire B_DAC[0];
	output wire B_DAC[1];
	output wire B_DAC[2];
	output wire B_DAC[3];
	output wire B_DAC[4];
	output wire B_DAC[5];
	output wire B_DAC[6];
	output wire B_DAC[7];
	output wire B_DAC[8];
	output wire G_DAC[9];
	output wire G_DAC[10];
	output wire G_DAC[11];
	output wire G_DAC[12];
	output wire G_DAC[13];
	output wire G_DAC[14];
	output wire G_DAC[15];
	output wire G_DAC[16];
	output wire B_DAC[9];
	output wire B_DAC[10];
	output wire B_DAC[11];
	output wire B_DAC[12];
	output wire B_DAC[13];
	output wire B_DAC[14];
	output wire B_DAC[15];
	output wire B_DAC[16];
	output wire nOE1;
	output wire nWE0;
	output wire nWE1;
	output wire nCAS1;
	output wire nRAS1;
	output wire AD_RD_DIR;
	output wire nYS;
	output wire nSC;
	output wire nSE0_1;
	output wire ADo[7];
	output wire ADo[6];
	output wire ADo[5];
	output wire ADo[4];
	output wire ADo[3];
	output wire ADo[2];
	output wire ADo[1];
	output wire ADo[0];
	output wire RDo[6];
	output wire RDo[5];
	output wire RDo[4];
	output wire RDo[3];
	output wire RDo[2];
	output wire RDo[1];
	output wire RDo[0];
	input wire RDi[6];
	input wire RDi[7];
	input wire RDi[4];
	input wire RDi[5];
	input wire RDi[2];
	input wire RDi[3];
	input wire RDi[0];
	input wire RDi[1];
	input wire ADi[6];
	input wire ADi[7];
	input wire ADi[4];
	input wire ADi[5];
	input wire ADi[2];
	input wire ADi[3];
	input wire ADi[0];
	input wire ADi[1];
	output wire RDo[7];
	input wire SD[7];
	input wire SD[6];
	input wire SD[5];
	input wire SD[4];
	input wire SD[3];
	input wire SD[2];
	input wire SD[1];
	input wire SD[0];
	output wire CLK1;
	output wire CLK0;
	input wire EDCLKi;
	output wire EDCLKo;
	input wire MCLK;
	output wire SUB_CLK;
	input wire nRES_PAD;
	input wire 68kCLKi;
	output wire EDCLKd;
	output wire CA_PAD_DIR;
	output wire DB_PAD_DIR;
	input wire SEL0_M3;
	input wire nPAL;
	input wire nHL;
	output wire SPA/Bo;
	input wire SPA/Bi;

	// Wires

	wire w1;
	wire H40;
	wire w3;
	wire w4;
	wire w5;
	wire w6;
	wire w7;
	wire w8;
	wire w9;
	wire w10;
	wire w11;
	wire w12;
	wire w13;
	wire w14;
	wire w15;
	wire w16;
	wire w17;
	wire w18;
	wire w19;
	wire w20;
	wire w21;
	wire w22;
	wire w23;
	wire w24;
	wire w25;
	wire w26;
	wire w27;
	wire w28;
	wire w29;
	wire w30;
	wire w31;
	wire w32;
	wire w33;
	wire w34;
	wire w35;
	wire w36;
	wire w37;
	wire w38;
	wire w39;
	wire w40;
	wire w41;
	wire w42;
	wire w43;
	wire w44;
	wire w45;
	wire w46;
	wire w47;
	wire w48;
	wire ODD/EVEN;
	wire w50;
	wire w51;
	wire w52;
	wire w53;
	wire w54;
	wire w55;
	wire w56;
	wire w57;
	wire w58;
	wire w59;
	wire FIFOo[7];
	wire FIFOo[6];
	wire FIFOo[5];
	wire FIFOo[4];
	wire FIFOo[3];
	wire FIFOo[2];
	wire FIFOo[1];
	wire FIFOo[0];
	wire w68;
	wire w69;
	wire w70;
	wire w71;
	wire w72;
	wire w73;
	wire w74;
	wire w75;
	wire w76;
	wire w77;
	wire w78;
	wire w79;
	wire w80;
	wire w81;
	wire w82;
	wire w83;
	wire VRAMA[8];
	wire w85;
	wire w86;
	wire w87;
	wire w88;
	wire w89;
	wire w90;
	wire w91;
	wire w92;
	wire w93;
	wire w94;
	wire w95;
	wire w96;
	wire w97;
	wire w98;
	wire w99;
	wire w100;
	wire w101;
	wire VPOS[9];
	wire w103;
	wire w104;
	wire w105;
	wire w106;
	wire HPOS[0];
	wire w108;
	wire w109;
	wire w110;
	wire w111;
	wire w112;
	wire w113;
	wire w114;
	wire w115;
	wire w116;
	wire VPOS[8];
	wire w118;
	wire w119;
	wire w120;
	wire w121;
	wire w122;
	wire w123;
	wire w124;
	wire w125;
	wire w126;
	wire w127;
	wire w128;
	wire w129;
	wire w130;
	wire w131;
	wire w132;
	wire w133;
	wire w134;
	wire AD_DATA[7];
	wire AD_DATA[6];
	wire AD_DATA[4];
	wire RD_DATA[2];
	wire RD_DATA[1];
	wire RD_DATA[0];
	wire AD_DATA[5];
	wire w142;
	wire w143;
	wire DCLK1;
	wire DCLK2;
	wire nDCLK1;
	wire nDCLK2;
	wire HCLK1;
	wire HCLK2;
	wire nHCLK1;
	wire nHCLK2;
	wire SYSRES;
	wire DB[0];
	wire DB[1];
	wire DB[2];
	wire DB[3];
	wire DB[4];
	wire DB[5];
	wire DB[6];
	wire DB[7];
	wire DB[8];
	wire DB[9];
	wire AD_DATA[3];
	wire AD_DATA[2];
	wire AD_DATA[1];
	wire AD_DATA[0];
	wire DB[14];
	wire DB[13];
	wire DB[12];
	wire DB[11];
	wire DB[10];
	wire w172;
	wire M5;
	wire w174;
	wire w175;
	wire w176;
	wire HPOS[1];
	wire w178;
	wire w179;
	wire w180;
	wire w181;
	wire w182;
	wire w183;
	wire w184;
	wire w185;
	wire w186;
	wire w187;
	wire w188;
	wire w189;
	wire w190;
	wire VPOS[2];
	wire HPOS[3];
	wire w193;
	wire w194;
	wire w195;
	wire w196;
	wire w197;
	wire w198;
	wire w199;
	wire w200;
	wire w201;
	wire w202;
	wire w203;
	wire w204;
	wire w205;
	wire VPOS[4];
	wire HPOS[5];
	wire w208;
	wire RD_DATA[4];
	wire w210;
	wire w211;
	wire w212;
	wire w213;
	wire w214;
	wire w215;
	wire w216;
	wire w217;
	wire w218;
	wire w219;
	wire w220;
	wire w221;
	wire HPOS[7];
	wire w223;
	wire RD_DATA[6];
	wire w225;
	wire w226;
	wire w227;
	wire w228;
	wire w229;
	wire w230;
	wire w231;
	wire w232;
	wire w233;
	wire w234;
	wire w235;
	wire w236;
	wire w237;
	wire w238;
	wire w239;
	wire w240;
	wire w241;
	wire w242;
	wire w243;
	wire w244;
	wire w245;
	wire w246;
	wire w247;
	wire w248;
	wire w249;
	wire w250;
	wire w251;
	wire w252;
	wire w253;
	wire w254;
	wire w255;
	wire w256;
	wire w257;
	wire w258;
	wire w259;
	wire w260;
	wire w261;
	wire w262;
	wire w263;
	wire w264;
	wire w265;
	wire w266;
	wire w267;
	wire w268;
	wire w269;
	wire w270;
	wire w271;
	wire w272;
	wire w273;
	wire w274;
	wire w275;
	wire w276;
	wire w277;
	wire w278;
	wire w279;
	wire w280;
	wire w281;
	wire w282;
	wire w283;
	wire w284;
	wire w285;
	wire w286;
	wire w287;
	wire w288;
	wire w289;
	wire w290;
	wire w291;
	wire w292;
	wire w293;
	wire w294;
	wire w295;
	wire w296;
	wire w297;
	wire w298;
	wire w299;
	wire w300;
	wire w301;
	wire w302;
	wire w303;
	wire w304;
	wire w305;
	wire w306;
	wire w307;
	wire w308;
	wire w309;
	wire HPOS[2];
	wire VPOS[1];
	wire w312;
	wire w313;
	wire w314;
	wire w315;
	wire w316;
	wire w317;
	wire w318;
	wire w319;
	wire w320;
	wire w321;
	wire w322;
	wire VPOS[3];
	wire w324;
	wire HPOS[4];
	wire w326;
	wire w327;
	wire w328;
	wire w329;
	wire w330;
	wire w331;
	wire w332;
	wire w333;
	wire w334;
	wire w335;
	wire w336;
	wire w337;
	wire w338;
	wire HPOS[6];
	wire VPOS[5];
	wire RD_DATA[5];
	wire w342;
	wire w343;
	wire w344;
	wire w345;
	wire w346;
	wire w347;
	wire w348;
	wire w349;
	wire w350;
	wire w351;
	wire w352;
	wire w353;
	wire w354;
	wire HPOS[8];
	wire VPOS[7];
	wire DB[15];
	wire w358;
	wire w359;
	wire w360;
	wire w361;
	wire w362;
	wire w363;
	wire w364;
	wire w365;
	wire w366;
	wire w367;
	wire w368;
	wire w369;
	wire w370;
	wire w371;
	wire w372;
	wire w373;
	wire w374;
	wire w375;
	wire w376;
	wire w377;
	wire w378;
	wire w379;
	wire w380;
	wire w381;
	wire w382;
	wire w383;
	wire w384;
	wire w385;
	wire w386;
	wire w387;
	wire w388;
	wire w389;
	wire w390;
	wire w391;
	wire w392;
	wire w393;
	wire w394;
	wire w395;
	wire w396;
	wire w397;
	wire w398;
	wire w399;
	wire w400;
	wire w401;
	wire w402;
	wire w403;
	wire w404;
	wire w405;
	wire w406;
	wire w407;
	wire w408;
	wire w409;
	wire w410;
	wire w411;
	wire w412;
	wire w413;
	wire w414;
	wire w415;
	wire w416;
	wire w417;
	wire w418;
	wire w419;
	wire w420;
	wire w421;
	wire w422;
	wire w423;
	wire w424;
	wire w425;
	wire w426;
	wire w427;
	wire w428;
	wire w429;
	wire w430;
	wire w431;
	wire w432;
	wire w433;
	wire w434;
	wire w435;
	wire w436;
	wire 128k;
	wire w438;
	wire w439;
	wire w440;
	wire w441;
	wire w442;
	wire w443;
	wire w444;
	wire w445;
	wire w446;
	wire w447;
	wire w448;
	wire w449;
	wire w450;
	wire w451;
	wire w452;
	wire w453;
	wire w454;
	wire w455;
	wire w456;
	wire w457;
	wire w458;
	wire w459;
	wire w460;
	wire w461;
	wire w462;
	wire w463;
	wire w464;
	wire w465;
	wire w466;
	wire w467;
	wire w468;
	wire w469;
	wire w470;
	wire w471;
	wire w472;
	wire w473;
	wire CA[0];
	wire w475;
	wire w476;
	wire w477;
	wire w478;
	wire w479;
	wire w480;
	wire w481;
	wire w482;
	wire w483;
	wire w484;
	wire w485;
	wire w486;
	wire w487;
	wire w488;
	wire w489;
	wire w490;
	wire w491;
	wire w492;
	wire w493;
	wire w494;
	wire w495;
	wire w496;
	wire w497;
	wire w498;
	wire w499;
	wire w500;
	wire w501;
	wire w502;
	wire w503;
	wire w504;
	wire w505;
	wire w506;
	wire w507;
	wire w508;
	wire w509;
	wire w510;
	wire w511;
	wire w512;
	wire w513;
	wire w514;
	wire w515;
	wire w516;
	wire w517;
	wire w518;
	wire w519;
	wire w520;
	wire w521;
	wire w522;
	wire w523;
	wire w524;
	wire w525;
	wire w526;
	wire w527;
	wire w528;
	wire w529;
	wire w530;
	wire w531;
	wire w532;
	wire w533;
	wire w534;
	wire w535;
	wire w536;
	wire w537;
	wire w538;
	wire w539;
	wire w540;
	wire w541;
	wire w542;
	wire w543;
	wire w544;
	wire w545;
	wire w546;
	wire w547;
	wire w548;
	wire w549;
	wire w550;
	wire w551;
	wire w552;
	wire w553;
	wire w554;
	wire w555;
	wire w556;
	wire w557;
	wire w558;
	wire w559;
	wire w560;
	wire w561;
	wire w562;
	wire w563;
	wire w564;
	wire VRAMA[0];
	wire w566;
	wire w567;
	wire w568;
	wire w569;
	wire w570;
	wire w571;
	wire w572;
	wire w573;
	wire w574;
	wire w575;
	wire w576;
	wire w577;
	wire w578;
	wire w579;
	wire w580;
	wire w581;
	wire w582;
	wire w583;
	wire w584;
	wire w585;
	wire w586;
	wire w587;
	wire w588;
	wire w589;
	wire w590;
	wire w591;
	wire w592;
	wire w593;
	wire w594;
	wire w595;
	wire w596;
	wire w597;
	wire w598;
	wire w599;
	wire w600;
	wire w601;
	wire DMA_BUSY;
	wire w603;
	wire w604;
	wire w605;
	wire w606;
	wire w607;
	wire w608;
	wire w609;
	wire REG_BUS[0];
	wire w611;
	wire w612;
	wire w613;
	wire w614;
	wire REG_BUS[7];
	wire w616;
	wire w617;
	wire w618;
	wire w619;
	wire w620;
	wire w621;
	wire w622;
	wire w623;
	wire w624;
	wire w625;
	wire w626;
	wire w627;
	wire w628;
	wire w629;
	wire w630;
	wire w631;
	wire w632;
	wire w633;
	wire w634;
	wire w635;
	wire w636;
	wire w637;
	wire w638;
	wire w639;
	wire CA[8];
	wire CA[7];
	wire w642;
	wire w643;
	wire w644;
	wire w645;
	wire w646;
	wire w647;
	wire w648;
	wire w649;
	wire w650;
	wire w651;
	wire w652;
	wire w653;
	wire w654;
	wire CA[9];
	wire w656;
	wire VRAMA[7];
	wire w658;
	wire REG_BUS[6];
	wire VRAMA[9];
	wire w661;
	wire CA[6];
	wire w663;
	wire w664;
	wire w665;
	wire w666;
	wire w667;
	wire w668;
	wire w669;
	wire w670;
	wire w671;
	wire w672;
	wire w673;
	wire w674;
	wire w675;
	wire w676;
	wire w677;
	wire REG_BUS[5];
	wire VRAMA[10];
	wire VRAMA[6];
	wire w681;
	wire REG_BUS[1];
	wire w683;
	wire w684;
	wire w685;
	wire w686;
	wire CA[10];
	wire w688;
	wire w689;
	wire w690;
	wire w691;
	wire w692;
	wire w693;
	wire w694;
	wire REG_BUS[2];
	wire w696;
	wire CA[11];
	wire w698;
	wire w699;
	wire w700;
	wire w701;
	wire w702;
	wire w703;
	wire w704;
	wire w705;
	wire w706;
	wire w707;
	wire VRAMA[5];
	wire w709;
	wire w710;
	wire VRAMA[11];
	wire CA[5];
	wire w713;
	wire w714;
	wire w715;
	wire REG_BUS[3];
	wire VRAMA[12];
	wire VRAMA[4];
	wire w719;
	wire w720;
	wire w721;
	wire REG_BUS[4];
	wire w723;
	wire CA[12];
	wire w725;
	wire w726;
	wire CA[4];
	wire w728;
	wire w729;
	wire w730;
	wire w731;
	wire CA[19];
	wire w733;
	wire w734;
	wire w735;
	wire w736;
	wire w737;
	wire VRAMA[13];
	wire w739;
	wire w740;
	wire w741;
	wire VRAMA[3];
	wire CA[3];
	wire w744;
	wire w745;
	wire CA[13];
	wire CA[20];
	wire w748;
	wire w749;
	wire w750;
	wire w751;
	wire w752;
	wire w753;
	wire VRAMA[14];
	wire VRAMA[2];
	wire w756;
	wire w757;
	wire w758;
	wire w759;
	wire w760;
	wire CA[2];
	wire w762;
	wire w763;
	wire w764;
	wire CA[21];
	wire w766;
	wire w767;
	wire w768;
	wire w769;
	wire w770;
	wire CA[14];
	wire w772;
	wire w773;
	wire VRAMA[15];
	wire CA[15];
	wire VRAMA[1];
	wire w777;
	wire w778;
	wire w779;
	wire w780;
	wire w781;
	wire w782;
	wire w783;
	wire w784;
	wire w785;
	wire w786;
	wire w787;
	wire CA[17];
	wire CA[1];
	wire VRAMA[16];
	wire w791;
	wire w792;
	wire CA[16];
	wire w794;
	wire w795;
	wire w796;
	wire w797;
	wire w798;
	wire w799;
	wire w800;
	wire w801;
	wire w802;
	wire w803;
	wire w804;
	wire w805;
	wire w806;
	wire w807;
	wire w808;
	wire w809;
	wire w810;
	wire w811;
	wire w812;
	wire w813;
	wire w814;
	wire w815;
	wire w816;
	wire w817;
	wire w818;
	wire w819;
	wire w820;
	wire w821;
	wire w822;
	wire w823;
	wire w824;
	wire w825;
	wire w826;
	wire w827;
	wire w828;
	wire w829;
	wire w830;
	wire w831;
	wire w832;
	wire w833;
	wire w834;
	wire w835;
	wire w836;
	wire w837;
	wire w838;
	wire w839;
	wire w840;
	wire w841;
	wire w842;
	wire w843;
	wire w844;
	wire w845;
	wire w846;
	wire w847;
	wire w848;
	wire w849;
	wire w850;
	wire w851;
	wire w852;
	wire w853;
	wire w854;
	wire w855;
	wire w856;
	wire w857;
	wire w858;
	wire w859;
	wire w860;
	wire w861;
	wire w862;
	wire w863;
	wire w864;
	wire w865;
	wire w866;
	wire w867;
	wire w868;
	wire w869;
	wire w870;
	wire w871;
	wire w872;
	wire w873;
	wire w874;
	wire w875;
	wire w876;
	wire w877;
	wire w878;
	wire w879;
	wire w880;
	wire w881;
	wire w882;
	wire w883;
	wire w884;
	wire w885;
	wire w886;
	wire w887;
	wire w888;
	wire w889;
	wire w890;
	wire w891;
	wire w892;
	wire w893;
	wire w894;
	wire w895;
	wire w896;
	wire w897;
	wire w898;
	wire w899;
	wire w900;
	wire w901;
	wire w902;
	wire w903;
	wire w904;
	wire w905;
	wire w906;
	wire w907;
	wire w908;
	wire w909;
	wire w910;
	wire w911;
	wire w912;
	wire w913;
	wire w914;
	wire w915;
	wire w916;
	wire w917;
	wire w918;
	wire w919;
	wire w920;
	wire w921;
	wire w922;
	wire w923;
	wire w924;
	wire w925;
	wire w926;
	wire w927;
	wire w928;
	wire w929;
	wire w930;
	wire w931;
	wire w932;
	wire w933;
	wire w934;
	wire w935;
	wire w936;
	wire w937;
	wire w938;
	wire w939;
	wire w940;
	wire w941;
	wire w942;
	wire w943;
	wire w944;
	wire w945;
	wire w946;
	wire w947;
	wire w948;
	wire w949;
	wire w950;
	wire w951;
	wire w952;
	wire w953;
	wire w954;
	wire w955;
	wire w956;
	wire w957;
	wire w958;
	wire w959;
	wire w960;
	wire w961;
	wire w962;
	wire w963;
	wire w964;
	wire w965;
	wire w966;
	wire w967;
	wire w968;
	wire w969;
	wire w970;
	wire w971;
	wire w972;
	wire w973;
	wire w974;
	wire w975;
	wire w976;
	wire w977;
	wire w978;
	wire w979;
	wire w980;
	wire w981;
	wire w982;
	wire w983;
	wire w984;
	wire w985;
	wire w986;
	wire w987;
	wire w988;
	wire w989;
	wire w990;
	wire w991;
	wire w992;
	wire w993;
	wire w994;
	wire w995;
	wire w996;
	wire w997;
	wire w998;
	wire w999;
	wire w1000;
	wire w1001;
	wire w1002;
	wire w1003;
	wire w1004;
	wire w1005;
	wire w1006;
	wire w1007;
	wire w1008;
	wire w1009;
	wire w1010;
	wire w1011;
	wire w1012;
	wire w1013;
	wire w1014;
	wire w1015;
	wire w1016;
	wire w1017;
	wire w1018;
	wire w1019;
	wire w1020;
	wire w1021;
	wire w1022;
	wire w1023;
	wire w1024;
	wire w1025;
	wire w1026;
	wire w1027;
	wire w1028;
	wire w1029;
	wire w1030;
	wire w1031;
	wire w1032;
	wire w1033;
	wire w1034;
	wire w1035;
	wire w1036;
	wire w1037;
	wire w1038;
	wire w1039;
	wire w1040;
	wire w1041;
	wire w1042;
	wire w1043;
	wire w1044;
	wire w1045;
	wire w1046;
	wire w1047;
	wire w1048;
	wire w1049;
	wire w1050;
	wire w1051;
	wire w1052;
	wire w1053;
	wire w1054;
	wire w1055;
	wire w1056;
	wire w1057;
	wire w1058;
	wire LS0;
	wire w1060;
	wire VPOS[0];
	wire w1062;
	wire w1063;
	wire w1064;
	wire w1065;
	wire w1066;
	wire w1067;
	wire w1068;
	wire w1069;
	wire w1070;
	wire w1071;
	wire w1072;
	wire w1073;
	wire w1074;
	wire w1075;
	wire w1076;
	wire w1077;
	wire w1078;
	wire w1079;
	wire w1080;
	wire w1081;
	wire w1082;
	wire w1083;
	wire COL[0];
	wire COL[1];
	wire COL[2];
	wire COL[3];
	wire COL[4];
	wire COL[5];
	wire COL[6];
	wire w1091;
	wire w1092;
	wire w1093;
	wire w1094;
	wire w1095;
	wire w1096;
	wire w1097;
	wire w1098;
	wire w1099;
	wire w1100;
	wire w1101;
	wire w1102;
	wire w1103;
	wire w1104;
	wire w1105;
	wire w1106;
	wire w1107;
	wire w1108;
	wire w1109;
	wire w1110;
	wire w1111;
	wire w1112;
	wire w1113;
	wire w1114;
	wire w1115;
	wire w1116;
	wire w1117;
	wire w1118;
	wire w1119;
	wire w1120;
	wire w1121;
	wire w1122;
	wire w1123;
	wire w1124;
	wire w1125;
	wire w1126;
	wire w1127;
	wire w1128;
	wire w1129;
	wire w1130;
	wire w1131;
	wire w1132;
	wire w1133;
	wire w1134;
	wire w1135;
	wire w1136;
	wire w1137;
	wire w1138;
	wire w1139;
	wire w1140;
	wire w1141;
	wire w1142;
	wire w1143;
	wire w1144;
	wire w1145;
	wire w1146;
	wire w1147;
	wire w1148;
	wire PSG_TEST_OE;
	wire w1150;
	wire w1151;
	wire w1152;
	wire w1153;
	wire w1154;
	wire w1155;
	wire w1156;
	wire w1157;
	wire w1158;
	wire w1159;
	wire w1160;
	wire w1161;
	wire w1162;
	wire w1163;
	wire w1164;
	wire w1165;
	wire w1166;
	wire w1167;
	wire w1168;
	wire w1169;
	wire w1170;
	wire w1171;
	wire w1172;
	wire w1173;
	wire w1174;
	wire w1175;
	wire w1176;
	wire w1177;
	wire w1178;
	wire w1179;
	wire w1180;
	wire w1181;
	wire w1182;
	wire w1183;
	wire w1184;
	wire w1185;
	wire w1186;
	wire w1187;
	wire w1188;
	wire w1189;
	wire w1190;
	wire w1191;
	wire w1192;
	wire w1193;
	wire w1194;
	wire w1195;
	wire w1196;
	wire w1197;
	wire w1198;
	wire w1199;
	wire w1200;
	wire w1201;
	wire PAL;
	wire w1203;
	wire w1204;
	wire w1205;
	wire w1206;
	wire w1207;
	wire w1208;
	wire w1209;
	wire w1210;
	wire w1211;
	wire w1212;
	wire w1213;
	wire w1214;
	wire w1215;
	wire w1216;
	wire w1217;
	wire w1218;
	wire w1219;
	wire w1220;
	wire w1221;
	wire w1222;
	wire w1223;
	wire w1224;
	wire w1225;
	wire w1226;
	wire w1227;
	wire w1228;
	wire w1229;
	wire w1230;
	wire w1231;
	wire w1232;
	wire w1233;
	wire w1234;
	wire w1235;
	wire w1236;
	wire w1237;
	wire w1238;
	wire w1239;
	wire w1240;
	wire w1241;
	wire w1242;
	wire w1243;
	wire w1244;
	wire w1245;
	wire w1246;
	wire w1247;
	wire w1248;
	wire w1249;
	wire w1250;
	wire w1251;
	wire w1252;
	wire w1253;
	wire w1254;
	wire w1255;
	wire w1256;
	wire w1257;
	wire w1258;
	wire w1259;
	wire w1260;
	wire w1261;
	wire w1262;
	wire w1263;
	wire w1264;
	wire w1265;
	wire w1266;
	wire w1267;
	wire w1268;
	wire w1269;
	wire w1270;
	wire w1271;
	wire w1272;
	wire w1273;
	wire w1274;
	wire w1275;
	wire w1276;
	wire w1277;
	wire w1278;
	wire w1279;
	wire w1280;
	wire w1281;
	wire w1282;
	wire w1283;
	wire w1284;
	wire w1285;
	wire w1286;
	wire w1287;
	wire w1288;
	wire w1289;
	wire w1290;
	wire w1291;
	wire w1292;
	wire w1293;
	wire w1294;
	wire w1295;
	wire w1296;
	wire w1297;
	wire w1298;
	wire w1299;
	wire w1300;
	wire w1301;
	wire w1302;
	wire w1303;
	wire w1304;
	wire w1305;
	wire w1306;
	wire w1307;
	wire w1308;
	wire w1309;
	wire w1310;
	wire w1311;
	wire w1312;
	wire w1313;
	wire w1314;
	wire w1315;
	wire w1316;
	wire w1317;
	wire w1318;
	wire w1319;
	wire w1320;
	wire w1321;
	wire w1322;
	wire w1323;
	wire w1324;
	wire w1325;
	wire w1326;
	wire w1327;
	wire w1328;
	wire w1329;
	wire w1330;
	wire w1331;
	wire w1332;
	wire w1333;
	wire w1334;
	wire w1335;
	wire w1336;
	wire w1337;
	wire w1338;
	wire w1339;
	wire w1340;
	wire w1341;
	wire w1342;
	wire w1343;
	wire w1344;
	wire w1345;
	wire w1346;
	wire w1347;
	wire w1348;
	wire w1349;
	wire w1350;
	wire w1351;
	wire w1352;
	wire w1353;
	wire w1354;
	wire w1355;
	wire w1356;
	wire w1357;
	wire w1358;
	wire w1359;
	wire w1360;
	wire w1361;
	wire w1362;
	wire w1363;
	wire w1364;
	wire w1365;
	wire w1366;
	wire w1367;
	wire w1368;
	wire w1369;
	wire w1370;
	wire w1371;
	wire w1372;
	wire w1373;
	wire w1374;
	wire w1375;
	wire w1376;
	wire w1377;
	wire w1378;
	wire w1379;
	wire w1380;
	wire w1381;
	wire w1382;
	wire w1383;
	wire w1384;
	wire w1385;
	wire w1386;
	wire w1387;
	wire w1388;
	wire w1389;
	wire w1390;
	wire w1391;
	wire w1392;
	wire w1393;
	wire w1394;
	wire VRAM_REFRESH;
	wire w1396;
	wire w1397;
	wire w1398;
	wire w1399;
	wire w1400;
	wire w1401;
	wire w1402;
	wire w1403;
	wire w1404;
	wire w1405;
	wire w1406;
	wire w1407;
	wire w1408;
	wire w1409;
	wire w1410;
	wire w1411;
	wire w1412;
	wire w1413;
	wire w1414;
	wire w1415;
	wire w1416;
	wire w1417;
	wire w1418;
	wire w1419;
	wire w1420;
	wire w1421;
	wire w1422;
	wire w1423;
	wire w1424;
	wire w1425;
	wire w1426;
	wire w1427;
	wire w1428;
	wire w1429;
	wire w1430;
	wire w1431;
	wire w1432;
	wire w1433;
	wire w1434;
	wire w1435;
	wire w1436;
	wire w1437;
	wire w1438;
	wire w1439;
	wire w1440;
	wire w1441;
	wire w1442;
	wire w1443;
	wire w1444;
	wire w1445;
	wire w1446;
	wire w1447;
	wire w1448;
	wire w1449;
	wire w1450;
	wire w1451;
	wire w1452;
	wire w1453;
	wire w1454;
	wire w1455;
	wire w1456;
	wire w1457;
	wire w1458;
	wire w1459;
	wire w1460;
	wire w1461;
	wire w1462;
	wire w1463;
	wire w1464;
	wire w1465;
	wire w1466;
	wire w1467;
	wire w1468;
	wire w1469;
	wire w1470;
	wire w1471;
	wire w1472;
	wire w1473;
	wire w1474;
	wire w1475;
	wire w1476;
	wire w1477;
	wire w1478;
	wire w1479;
	wire w1480;
	wire w1481;
	wire w1482;
	wire w1483;
	wire w1484;
	wire w1485;
	wire w1486;
	wire w1487;
	wire w1488;
	wire w1489;
	wire w1490;
	wire w1491;
	wire w1492;
	wire w1493;
	wire w1494;
	wire w1495;
	wire w1496;
	wire w1497;
	wire w1498;
	wire w1499;
	wire w1500;
	wire w1501;
	wire w1502;
	wire w1503;
	wire w1504;
	wire w1505;
	wire w1506;
	wire w1507;
	wire CA[18];
	wire w1509;
	wire w1510;
	wire w1511;
	wire w1512;
	wire w1513;
	wire w1514;
	wire w1515;
	wire w1516;
	wire w1517;
	wire w1518;
	wire w1519;
	wire w1520;
	wire w1521;
	wire w1522;
	wire w1523;
	wire w1524;
	wire w1525;
	wire w1526;
	wire w1527;
	wire w1528;
	wire w1529;
	wire w1530;
	wire w1531;
	wire w1532;
	wire w1533;
	wire w1534;
	wire w1535;
	wire w1536;
	wire w1537;
	wire w1538;
	wire w1539;
	wire w1540;
	wire w1541;
	wire w1542;
	wire w1543;
	wire w1544;
	wire w1545;
	wire w1546;
	wire w1547;
	wire w1548;
	wire w1549;
	wire w1550;
	wire w1551;
	wire w1552;
	wire w1553;
	wire w1554;
	wire w1555;
	wire w1556;
	wire w1557;
	wire w1558;
	wire w1559;
	wire w1560;
	wire w1561;
	wire w1562;
	wire w1563;
	wire w1564;
	wire w1565;
	wire w1566;
	wire w1567;
	wire w1568;
	wire w1569;
	wire VPOS[6];
	wire w1571;
	wire w1572;
	wire w1573;
	wire w1574;
	wire w1575;
	wire w1576;
	wire w1577;
	wire w1578;
	wire w1579;
	wire w1580;
	wire w1581;
	wire w1582;
	wire w1583;
	wire w1584;
	wire w1585;
	wire w1586;
	wire w1587;
	wire w1588;
	wire w1589;
	wire w1590;
	wire w1591;
	wire w1592;
	wire w1593;
	wire w1594;
	wire w1595;
	wire w1596;
	wire w1597;
	wire w1598;
	wire w1599;
	wire w1600;
	wire w1601;
	wire w1602;
	wire w1603;
	wire w1604;
	wire w1605;
	wire w1606;
	wire w1607;
	wire w1608;
	wire w1609;
	wire w1610;
	wire w1611;
	wire w1612;
	wire w1613;
	wire w1614;
	wire w1615;
	wire w1616;
	wire w1617;
	wire w1618;
	wire w1619;
	wire w1620;
	wire w1621;
	wire w1622;
	wire w1623;
	wire w1624;
	wire w1625;
	wire w1626;
	wire w1627;
	wire w1628;
	wire w1629;
	wire w1630;
	wire w1631;
	wire w1632;
	wire w1633;
	wire w1634;
	wire w1635;
	wire w1636;
	wire w1637;
	wire w1638;
	wire w1639;
	wire w1640;
	wire w1641;
	wire w1642;
	wire w1643;
	wire w1644;
	wire w1645;
	wire w1646;
	wire w1647;
	wire w1648;
	wire w1649;
	wire w1650;
	wire w1651;
	wire w1652;
	wire w1653;
	wire w1654;
	wire w1655;
	wire w1656;
	wire w1657;
	wire w1658;
	wire w1659;
	wire w1660;
	wire w1661;
	wire w1662;
	wire w1663;
	wire w1664;
	wire w1665;
	wire w1666;
	wire w1667;
	wire w1668;
	wire w1669;
	wire w1670;
	wire w1671;
	wire w1672;
	wire w1673;
	wire w1674;
	wire w1675;
	wire w1676;
	wire w1677;
	wire w1678;
	wire w1679;
	wire w1680;
	wire w1681;
	wire w1682;
	wire w1683;
	wire w1684;
	wire w1685;
	wire w1686;
	wire w1687;
	wire w1688;
	wire w1689;
	wire w1690;
	wire w1691;
	wire w1692;
	wire w1693;
	wire w1694;
	wire w1695;
	wire w1696;
	wire w1697;
	wire w1698;
	wire w1699;
	wire w1700;
	wire w1701;
	wire w1702;
	wire w1703;
	wire w1704;
	wire w1705;
	wire w1706;
	wire w1707;
	wire w1708;
	wire w1709;
	wire w1710;
	wire w1711;
	wire w1712;
	wire w1713;
	wire w1714;
	wire w1715;
	wire w1716;
	wire w1717;
	wire w1718;
	wire w1719;
	wire w1720;
	wire w1721;
	wire w1722;
	wire w1723;
	wire w1724;
	wire w1725;
	wire w1726;
	wire w1727;
	wire w1728;
	wire w1729;
	wire w1730;
	wire w1731;
	wire w1732;
	wire w1733;
	wire w1734;
	wire w1735;
	wire w1736;
	wire w1737;
	wire w1738;
	wire w1739;
	wire w1740;
	wire w1741;
	wire w1742;
	wire w1743;
	wire w1744;
	wire w1745;
	wire w1746;
	wire w1747;
	wire w1748;
	wire w1749;
	wire w1750;
	wire w1751;
	wire w1752;
	wire w1753;
	wire w1754;
	wire w1755;
	wire w1756;
	wire w1757;
	wire w1758;
	wire w1759;
	wire w1760;
	wire w1761;
	wire w1762;
	wire w1763;
	wire w1764;
	wire w1765;
	wire w1766;
	wire w1767;
	wire w1768;
	wire w1769;
	wire w1770;
	wire w1771;
	wire w1772;
	wire w1773;
	wire w1774;
	wire w1775;
	wire w1776;
	wire w1777;
	wire w1778;
	wire w1779;
	wire w1780;
	wire w1781;
	wire w1782;
	wire w1783;
	wire w1784;
	wire w1785;
	wire w1786;
	wire w1787;
	wire w1788;
	wire w1789;
	wire w1790;
	wire w1791;
	wire w1792;
	wire w1793;
	wire w1794;
	wire w1795;
	wire w1796;
	wire w1797;
	wire w1798;
	wire w1799;
	wire w1800;
	wire w1801;
	wire w1802;
	wire w1803;
	wire w1804;
	wire w1805;
	wire w1806;
	wire w1807;
	wire w1808;
	wire w1809;
	wire w1810;
	wire w1811;
	wire w1812;
	wire w1813;
	wire w1814;
	wire w1815;
	wire w1816;
	wire w1817;
	wire w1818;
	wire w1819;
	wire w1820;
	wire w1821;
	wire w1822;
	wire w1823;
	wire w1824;
	wire w1825;
	wire w1826;
	wire w1827;
	wire w1828;
	wire w1829;
	wire w1830;
	wire w1831;
	wire w1832;
	wire w1833;
	wire w1834;
	wire w1835;
	wire w1836;
	wire w1837;
	wire w1838;
	wire w1839;
	wire w1840;
	wire w1841;
	wire w1842;
	wire w1843;
	wire w1844;
	wire w1845;
	wire w1846;
	wire w1847;
	wire w1848;
	wire w1849;
	wire w1850;
	wire w1851;
	wire w1852;
	wire w1853;
	wire w1854;
	wire w1855;
	wire w1856;
	wire w1857;
	wire w1858;
	wire w1859;
	wire w1860;
	wire w1861;
	wire w1862;
	wire w1863;
	wire w1864;
	wire w1865;
	wire w1866;
	wire w1867;
	wire w1868;
	wire w1869;
	wire w1870;
	wire w1871;
	wire w1872;
	wire w1873;
	wire w1874;
	wire w1875;
	wire w1876;
	wire w1877;
	wire w1878;
	wire w1879;
	wire w1880;
	wire w1881;
	wire w1882;
	wire w1883;
	wire w1884;
	wire w1885;
	wire w1886;
	wire w1887;
	wire w1888;
	wire w1889;
	wire w1890;
	wire w1891;
	wire w1892;
	wire w1893;
	wire w1894;
	wire w1895;
	wire w1896;
	wire w1897;
	wire w1898;
	wire w1899;
	wire w1900;
	wire w1901;
	wire w1902;
	wire w1903;
	wire w1904;
	wire w1905;
	wire w1906;
	wire w1907;
	wire w1908;
	wire w1909;
	wire w1910;
	wire w1911;
	wire w1912;
	wire w1913;
	wire w1914;
	wire w1915;
	wire w1916;
	wire w1917;
	wire w1918;
	wire w1919;
	wire w1920;
	wire w1921;
	wire w1922;
	wire w1923;
	wire w1924;
	wire w1925;
	wire w1926;
	wire w1927;
	wire w1928;
	wire w1929;
	wire w1930;
	wire w1931;
	wire w1932;
	wire w1933;
	wire w1934;
	wire w1935;
	wire w1936;
	wire w1937;
	wire w1938;
	wire w1939;
	wire w1940;
	wire w1941;
	wire w1942;
	wire w1943;
	wire w1944;
	wire w1945;
	wire w1946;
	wire w1947;
	wire w1948;
	wire w1949;
	wire w1950;
	wire w1951;
	wire w1952;
	wire w1953;
	wire w1954;
	wire w1955;
	wire w1956;
	wire w1957;
	wire w1958;
	wire w1959;
	wire w1960;
	wire w1961;
	wire w1962;
	wire w1963;
	wire w1964;
	wire w1965;
	wire w1966;
	wire w1967;
	wire w1968;
	wire w1969;
	wire w1970;
	wire w1971;
	wire w1972;
	wire w1973;
	wire w1974;
	wire w1975;
	wire w1976;
	wire w1977;
	wire w1978;
	wire w1979;
	wire w1980;
	wire w1981;
	wire w1982;
	wire w1983;
	wire w1984;
	wire w1985;
	wire w1986;
	wire w1987;
	wire w1988;
	wire w1989;
	wire w1990;
	wire w1991;
	wire w1992;
	wire w1993;
	wire w1994;
	wire w1995;
	wire w1996;
	wire w1997;
	wire w1998;
	wire w1999;
	wire w2000;
	wire w2001;
	wire w2002;
	wire w2003;
	wire w2004;
	wire w2005;
	wire w2006;
	wire w2007;
	wire w2008;
	wire w2009;
	wire w2010;
	wire w2011;
	wire w2012;
	wire w2013;
	wire w2014;
	wire w2015;
	wire w2016;
	wire w2017;
	wire w2018;
	wire w2019;
	wire w2020;
	wire w2021;
	wire w2022;
	wire w2023;
	wire w2024;
	wire w2025;
	wire w2026;
	wire w2027;
	wire w2028;
	wire w2029;
	wire w2030;
	wire w2031;
	wire w2032;
	wire w2033;
	wire w2034;
	wire w2035;
	wire w2036;
	wire w2037;
	wire w2038;
	wire w2039;
	wire w2040;
	wire w2041;
	wire w2042;
	wire w2043;
	wire w2044;
	wire w2045;
	wire w2046;
	wire w2047;
	wire w2048;
	wire w2049;
	wire w2050;
	wire w2051;
	wire w2052;
	wire w2053;
	wire w2054;
	wire w2055;
	wire w2056;
	wire w2057;
	wire w2058;
	wire w2059;
	wire w2060;
	wire w2061;
	wire w2062;
	wire w2063;
	wire w2064;
	wire w2065;
	wire w2066;
	wire w2067;
	wire w2068;
	wire w2069;
	wire w2070;
	wire w2071;
	wire w2072;
	wire w2073;
	wire w2074;
	wire w2075;
	wire w2076;
	wire w2077;
	wire w2078;
	wire w2079;
	wire w2080;
	wire w2081;
	wire w2082;
	wire w2083;
	wire w2084;
	wire w2085;
	wire w2086;
	wire w2087;
	wire w2088;
	wire w2089;
	wire w2090;
	wire w2091;
	wire w2092;
	wire w2093;
	wire w2094;
	wire w2095;
	wire w2096;
	wire w2097;
	wire w2098;
	wire w2099;
	wire w2100;
	wire w2101;
	wire w2102;
	wire w2103;
	wire w2104;
	wire w2105;
	wire w2106;
	wire w2107;
	wire w2108;
	wire w2109;
	wire w2110;
	wire w2111;
	wire w2112;
	wire w2113;
	wire w2114;
	wire w2115;
	wire w2116;
	wire w2117;
	wire w2118;
	wire w2119;
	wire w2120;
	wire w2121;
	wire w2122;
	wire w2123;
	wire w2124;
	wire w2125;
	wire w2126;
	wire w2127;
	wire w2128;
	wire w2129;
	wire w2130;
	wire w2131;
	wire w2132;
	wire w2133;
	wire w2134;
	wire w2135;
	wire w2136;
	wire w2137;
	wire w2138;
	wire w2139;
	wire w2140;
	wire w2141;
	wire w2142;
	wire w2143;
	wire w2144;
	wire w2145;
	wire w2146;
	wire w2147;
	wire w2148;
	wire w2149;
	wire w2150;
	wire w2151;
	wire w2152;
	wire w2153;
	wire w2154;
	wire w2155;
	wire w2156;
	wire w2157;
	wire w2158;
	wire w2159;
	wire w2160;
	wire w2161;
	wire w2162;
	wire w2163;
	wire w2164;
	wire w2165;
	wire w2166;
	wire w2167;
	wire w2168;
	wire w2169;
	wire w2170;
	wire w2171;
	wire w2172;
	wire w2173;
	wire w2174;
	wire w2175;
	wire w2176;
	wire w2177;
	wire w2178;
	wire w2179;
	wire w2180;
	wire w2181;
	wire w2182;
	wire w2183;
	wire w2184;
	wire w2185;
	wire w2186;
	wire w2187;
	wire w2188;
	wire w2189;
	wire w2190;
	wire w2191;
	wire w2192;
	wire w2193;
	wire w2194;
	wire w2195;
	wire w2196;
	wire w2197;
	wire w2198;
	wire w2199;
	wire w2200;
	wire w2201;
	wire w2202;
	wire w2203;
	wire w2204;
	wire w2205;
	wire w2206;
	wire w2207;
	wire w2208;
	wire w2209;
	wire w2210;
	wire w2211;
	wire w2212;
	wire w2213;
	wire w2214;
	wire w2215;
	wire w2216;
	wire w2217;
	wire w2218;
	wire w2219;
	wire w2220;
	wire w2221;
	wire w2222;
	wire w2223;
	wire w2224;
	wire w2225;
	wire w2226;
	wire w2227;
	wire w2228;
	wire w2229;
	wire w2230;
	wire w2231;
	wire w2232;
	wire w2233;
	wire w2234;
	wire w2235;
	wire w2236;
	wire w2237;
	wire w2238;
	wire w2239;
	wire w2240;
	wire w2241;
	wire w2242;
	wire w2243;
	wire w2244;
	wire w2245;
	wire w2246;
	wire w2247;
	wire w2248;
	wire w2249;
	wire w2250;
	wire w2251;
	wire w2252;
	wire w2253;
	wire w2254;
	wire w2255;
	wire w2256;
	wire w2257;
	wire w2258;
	wire w2259;
	wire w2260;
	wire w2261;
	wire w2262;
	wire w2263;
	wire w2264;
	wire w2265;
	wire w2266;
	wire w2267;
	wire w2268;
	wire w2269;
	wire w2270;
	wire w2271;
	wire w2272;
	wire w2273;
	wire w2274;
	wire w2275;
	wire w2276;
	wire w2277;
	wire w2278;
	wire w2279;
	wire w2280;
	wire w2281;
	wire w2282;
	wire w2283;
	wire w2284;
	wire w2285;
	wire w2286;
	wire w2287;
	wire w2288;
	wire w2289;
	wire w2290;
	wire w2291;
	wire w2292;
	wire w2293;
	wire w2294;
	wire w2295;
	wire w2296;
	wire w2297;
	wire w2298;
	wire w2299;
	wire w2300;
	wire w2301;
	wire w2302;
	wire w2303;
	wire w2304;
	wire w2305;
	wire w2306;
	wire w2307;
	wire w2308;
	wire w2309;
	wire w2310;
	wire w2311;
	wire w2312;
	wire w2313;
	wire w2314;
	wire w2315;
	wire w2316;
	wire w2317;
	wire w2318;
	wire w2319;
	wire w2320;
	wire w2321;
	wire w2322;
	wire w2323;
	wire w2324;
	wire w2325;
	wire w2326;
	wire w2327;
	wire w2328;
	wire w2329;
	wire w2330;
	wire w2331;
	wire w2332;
	wire w2333;
	wire w2334;
	wire w2335;
	wire w2336;
	wire w2337;
	wire w2338;
	wire w2339;
	wire w2340;
	wire w2341;
	wire w2342;
	wire w2343;
	wire w2344;
	wire w2345;
	wire w2346;
	wire w2347;
	wire w2348;
	wire w2349;
	wire w2350;
	wire w2351;
	wire w2352;
	wire w2353;
	wire w2354;
	wire w2355;
	wire w2356;
	wire w2357;
	wire w2358;
	wire w2359;
	wire w2360;
	wire w2361;
	wire w2362;
	wire w2363;
	wire w2364;
	wire w2365;
	wire w2366;
	wire w2367;
	wire w2368;
	wire w2369;
	wire w2370;
	wire w2371;
	wire w2372;
	wire w2373;
	wire w2374;
	wire w2375;
	wire w2376;
	wire w2377;
	wire w2378;
	wire w2379;
	wire w2380;
	wire w2381;
	wire w2382;
	wire w2383;
	wire w2384;
	wire w2385;
	wire w2386;
	wire w2387;
	wire w2388;
	wire w2389;
	wire w2390;
	wire w2391;
	wire w2392;
	wire w2393;
	wire w2394;
	wire w2395;
	wire w2396;
	wire w2397;
	wire w2398;
	wire w2399;
	wire w2400;
	wire w2401;
	wire w2402;
	wire w2403;
	wire w2404;
	wire w2405;
	wire w2406;
	wire w2407;
	wire w2408;
	wire w2409;
	wire w2410;
	wire w2411;
	wire w2412;
	wire w2413;
	wire w2414;
	wire w2415;
	wire w2416;
	wire w2417;
	wire w2418;
	wire w2419;
	wire w2420;
	wire w2421;
	wire w2422;
	wire w2423;
	wire w2424;
	wire w2425;
	wire w2426;
	wire w2427;
	wire w2428;
	wire w2429;
	wire w2430;
	wire w2431;
	wire w2432;
	wire w2433;
	wire w2434;
	wire w2435;
	wire w2436;
	wire w2437;
	wire w2438;
	wire w2439;
	wire w2440;
	wire w2441;
	wire w2442;
	wire w2443;
	wire w2444;
	wire w2445;
	wire w2446;
	wire w2447;
	wire w2448;
	wire w2449;
	wire w2450;
	wire w2451;
	wire w2452;
	wire w2453;
	wire w2454;
	wire w2455;
	wire w2456;
	wire w2457;
	wire w2458;
	wire w2459;
	wire w2460;
	wire w2461;
	wire w2462;
	wire w2463;
	wire w2464;
	wire w2465;
	wire w2466;
	wire w2467;
	wire w2468;
	wire w2469;
	wire w2470;
	wire w2471;
	wire w2472;
	wire w2473;
	wire w2474;
	wire w2475;
	wire w2476;
	wire w2477;
	wire w2478;
	wire w2479;
	wire w2480;
	wire w2481;
	wire w2482;
	wire w2483;
	wire w2484;
	wire w2485;
	wire w2486;
	wire w2487;
	wire w2488;
	wire w2489;
	wire w2490;
	wire w2491;
	wire w2492;
	wire w2493;
	wire w2494;
	wire w2495;
	wire w2496;
	wire w2497;
	wire w2498;
	wire w2499;
	wire w2500;
	wire w2501;
	wire w2502;
	wire w2503;
	wire w2504;
	wire w2505;
	wire w2506;
	wire w2507;
	wire w2508;
	wire w2509;
	wire w2510;
	wire w2511;
	wire w2512;
	wire w2513;
	wire w2514;
	wire w2515;
	wire w2516;
	wire w2517;
	wire w2518;
	wire w2519;
	wire w2520;
	wire w2521;
	wire w2522;
	wire w2523;
	wire w2524;
	wire w2525;
	wire w2526;
	wire w2527;
	wire w2528;
	wire w2529;
	wire w2530;
	wire w2531;
	wire w2532;
	wire w2533;
	wire w2534;
	wire w2535;
	wire w2536;
	wire w2537;
	wire w2538;
	wire w2539;
	wire w2540;
	wire w2541;
	wire w2542;
	wire w2543;
	wire w2544;
	wire w2545;
	wire w2546;
	wire w2547;
	wire w2548;
	wire w2549;
	wire w2550;
	wire w2551;
	wire w2552;
	wire w2553;
	wire w2554;
	wire w2555;
	wire w2556;
	wire w2557;
	wire w2558;
	wire w2559;
	wire w2560;
	wire w2561;
	wire w2562;
	wire w2563;
	wire w2564;
	wire w2565;
	wire w2566;
	wire w2567;
	wire w2568;
	wire w2569;
	wire w2570;
	wire w2571;
	wire w2572;
	wire w2573;
	wire w2574;
	wire w2575;
	wire w2576;
	wire w2577;
	wire w2578;
	wire w2579;
	wire w2580;
	wire w2581;
	wire w2582;
	wire w2583;
	wire w2584;
	wire w2585;
	wire w2586;
	wire w2587;
	wire w2588;
	wire w2589;
	wire w2590;
	wire w2591;
	wire w2592;
	wire w2593;
	wire w2594;
	wire w2595;
	wire w2596;
	wire w2597;
	wire w2598;
	wire w2599;
	wire w2600;
	wire w2601;
	wire w2602;
	wire w2603;
	wire w2604;
	wire w2605;
	wire w2606;
	wire w2607;
	wire w2608;
	wire w2609;
	wire w2610;
	wire w2611;
	wire w2612;
	wire w2613;
	wire w2614;
	wire w2615;
	wire w2616;
	wire w2617;
	wire w2618;
	wire w2619;
	wire w2620;
	wire w2621;
	wire w2622;
	wire w2623;
	wire w2624;
	wire w2625;
	wire w2626;
	wire w2627;
	wire w2628;
	wire w2629;
	wire w2630;
	wire w2631;
	wire RES;
	wire w2633;
	wire w2634;
	wire w2635;
	wire w2636;
	wire EDCLK_O;
	wire nYS;
	wire w2639;
	wire w2640;
	wire w2641;
	wire w2642;
	wire w2643;
	wire w2644;
	wire w2645;
	wire w2646;
	wire w2647;
	wire w2648;
	wire w2649;
	wire w2650;
	wire w2651;
	wire w2652;
	wire w2653;
	wire w2654;
	wire w2655;
	wire w2656;
	wire w2657;
	wire w2658;
	wire w2659;
	wire w2660;
	wire w2661;
	wire w2662;
	wire w2663;
	wire w2664;
	wire w2665;
	wire w2666;
	wire w2667;
	wire w2668;
	wire w2669;
	wire w2670;
	wire w2671;
	wire w2672;
	wire w2673;
	wire w2674;
	wire w2675;
	wire w2676;
	wire w2677;
	wire w2678;
	wire w2679;
	wire w2680;
	wire w2681;
	wire w2682;
	wire w2683;
	wire w2684;
	wire w2685;
	wire w2686;
	wire w2687;
	wire w2688;
	wire w2689;
	wire w2690;
	wire w2691;
	wire w2692;
	wire w2693;
	wire w2694;
	wire w2695;
	wire w2696;
	wire w2697;
	wire w2698;
	wire w2699;
	wire w2700;
	wire w2701;
	wire w2702;
	wire w2703;
	wire SPR_PRIO;
	wire w2705;
	wire w2706;
	wire w2707;
	wire w2708;
	wire w2709;
	wire w2710;
	wire w2711;
	wire w2712;
	wire w2713;
	wire w2714;
	wire w2715;
	wire w2716;
	wire w2717;
	wire w2718;
	wire w2719;
	wire w2720;
	wire w2721;
	wire w2722;
	wire w2723;
	wire w2724;
	wire w2725;
	wire w2726;
	wire w2727;
	wire w2728;
	wire w2729;
	wire w2730;
	wire w2731;
	wire w2732;
	wire w2733;
	wire w2734;
	wire w2735;
	wire w2736;
	wire w2737;
	wire w2738;
	wire w2739;
	wire w2740;
	wire w2741;
	wire w2742;
	wire w2743;
	wire w2744;
	wire w2745;
	wire w2746;
	wire w2747;
	wire w2748;
	wire w2749;
	wire w2750;
	wire w2751;
	wire w2752;
	wire w2753;
	wire w2754;
	wire w2755;
	wire w2756;
	wire w2757;
	wire w2758;
	wire w2759;
	wire w2760;
	wire w2761;
	wire w2762;
	wire w2763;
	wire w2764;
	wire w2765;
	wire w2766;
	wire w2767;
	wire w2768;
	wire w2769;
	wire w2770;
	wire w2771;
	wire w2772;
	wire w2773;
	wire PLANE_A_PRIO;
	wire PLANE_B_PRIO;
	wire w2776;
	wire w2777;
	wire w2778;
	wire w2779;
	wire w2780;
	wire w2781;
	wire w2782;
	wire w2783;
	wire w2784;
	wire w2785;
	wire w2786;
	wire w2787;
	wire w2788;
	wire w2789;
	wire w2790;
	wire w2791;
	wire w2792;
	wire w2793;
	wire w2794;
	wire w2795;
	wire w2796;
	wire w2797;
	wire w2798;
	wire w2799;
	wire w2800;
	wire w2801;
	wire w2802;
	wire w2803;
	wire w2804;
	wire w2805;
	wire w2806;
	wire w2807;
	wire w2808;
	wire w2809;
	wire w2810;
	wire w2811;
	wire w2812;
	wire w2813;
	wire w2814;
	wire w2815;
	wire w2816;
	wire w2817;
	wire w2818;
	wire w2819;
	wire w2820;
	wire w2821;
	wire w2822;
	wire w2823;
	wire w2824;
	wire w2825;
	wire w2826;
	wire w2827;
	wire w2828;
	wire w2829;
	wire w2830;
	wire w2831;
	wire w2832;
	wire w2833;
	wire w2834;
	wire w2835;
	wire w2836;
	wire w2837;
	wire w2838;
	wire w2839;
	wire w2840;
	wire w2841;
	wire w2842;
	wire w2843;
	wire w2844;
	wire w2845;
	wire w2846;
	wire w2847;
	wire w2848;
	wire w2849;
	wire w2850;
	wire w2851;
	wire w2852;
	wire w2853;
	wire w2854;
	wire w2855;
	wire w2856;
	wire w2857;
	wire w2858;
	wire w2859;
	wire w2860;
	wire w2861;
	wire w2862;
	wire w2863;
	wire w2864;
	wire w2865;
	wire w2866;
	wire w2867;
	wire w2868;
	wire w2869;
	wire w2870;
	wire w2871;
	wire w2872;
	wire w2873;
	wire w2874;
	wire w2875;
	wire w2876;
	wire w2877;
	wire w2878;
	wire w2879;
	wire w2880;
	wire w2881;
	wire w2882;
	wire w2883;
	wire w2884;
	wire w2885;
	wire w2886;
	wire w2887;
	wire w2888;
	wire w2889;
	wire w2890;
	wire w2891;
	wire w2892;
	wire w2893;
	wire w2894;
	wire w2895;
	wire w2896;
	wire w2897;
	wire w2898;
	wire w2899;
	wire w2900;
	wire w2901;
	wire w2902;
	wire w2903;
	wire w2904;
	wire w2905;
	wire w2906;
	wire w2907;
	wire w2908;
	wire w2909;
	wire w2910;
	wire w2911;
	wire w2912;
	wire w2913;
	wire w2914;
	wire w2915;
	wire w2916;
	wire w2917;
	wire w2918;
	wire w2919;
	wire w2920;
	wire w2921;
	wire w2922;
	wire w2923;
	wire w2924;
	wire w2925;
	wire w2926;
	wire w2927;
	wire w2928;
	wire w2929;
	wire w2930;
	wire w2931;
	wire w2932;
	wire w2933;
	wire w2934;
	wire w2935;
	wire w2936;
	wire w2937;
	wire w2938;
	wire w2939;
	wire w2940;
	wire w2941;
	wire w2942;
	wire w2943;
	wire w2944;
	wire w2945;
	wire w2946;
	wire w2947;
	wire w2948;
	wire w2949;
	wire w2950;
	wire w2951;
	wire w2952;
	wire w2953;
	wire w2954;
	wire w2955;
	wire w2956;
	wire w2957;
	wire w2958;
	wire w2959;
	wire w2960;
	wire w2961;
	wire w2962;
	wire w2963;
	wire w2964;
	wire w2965;
	wire w2966;
	wire w2967;
	wire w2968;
	wire w2969;
	wire w2970;
	wire w2971;
	wire w2972;
	wire w2973;
	wire w2974;
	wire w2975;
	wire w2976;
	wire w2977;
	wire w2978;
	wire w2979;
	wire w2980;
	wire w2981;
	wire w2982;
	wire w2983;
	wire w2984;
	wire w2985;
	wire w2986;
	wire w2987;
	wire w2988;
	wire w2989;
	wire w2990;
	wire w2991;
	wire w2992;
	wire w2993;
	wire w2994;
	wire w2995;
	wire w2996;
	wire w2997;
	wire w2998;
	wire w2999;
	wire w3000;
	wire w3001;
	wire w3002;
	wire w3003;
	wire w3004;
	wire w3005;
	wire w3006;
	wire w3007;
	wire w3008;
	wire w3009;
	wire w3010;
	wire w3011;
	wire w3012;
	wire w3013;
	wire w3014;
	wire w3015;
	wire w3016;
	wire w3017;
	wire w3018;
	wire w3019;
	wire w3020;
	wire w3021;
	wire w3022;
	wire w3023;
	wire w3024;
	wire w3025;
	wire w3026;
	wire w3027;
	wire w3028;
	wire w3029;
	wire w3030;
	wire w3031;
	wire w3032;
	wire w3033;
	wire w3034;
	wire w3035;
	wire w3036;
	wire w3037;
	wire w3038;
	wire w3039;
	wire w3040;
	wire w3041;
	wire w3042;
	wire w3043;
	wire w3044;
	wire w3045;
	wire w3046;
	wire w3047;
	wire w3048;
	wire w3049;
	wire w3050;
	wire w3051;
	wire w3052;
	wire w3053;
	wire w3054;
	wire w3055;
	wire w3056;
	wire S[3];
	wire w3058;
	wire w3059;
	wire S[7];
	wire S[2];
	wire w3062;
	wire w3063;
	wire w3064;
	wire w3065;
	wire w3066;
	wire w3067;
	wire S[6];
	wire S[1];
	wire S[5];
	wire S[0];
	wire S[4];
	wire w3073;
	wire w3074;
	wire w3075;
	wire w3076;
	wire w3077;
	wire w3078;
	wire w3079;
	wire w3080;
	wire w3081;
	wire w3082;
	wire w3083;
	wire w3084;
	wire w3085;
	wire w3086;
	wire w3087;
	wire w3088;
	wire w3089;
	wire w3090;
	wire w3091;
	wire w3092;
	wire w3093;
	wire w3094;
	wire w3095;
	wire w3096;
	wire w3097;
	wire w3098;
	wire w3099;
	wire w3100;
	wire w3101;
	wire w3102;
	wire w3103;
	wire w3104;
	wire w3105;
	wire w3106;
	wire w3107;
	wire w3108;
	wire w3109;
	wire w3110;
	wire w3111;
	wire w3112;
	wire w3113;
	wire w3114;
	wire w3115;
	wire w3116;
	wire w3117;
	wire w3118;
	wire w3119;
	wire w3120;
	wire w3121;
	wire w3122;
	wire w3123;
	wire w3124;
	wire w3125;
	wire w3126;
	wire w3127;
	wire w3128;
	wire w3129;
	wire w3130;
	wire w3131;
	wire w3132;
	wire w3133;
	wire w3134;
	wire w3135;
	wire w3136;
	wire w3137;
	wire w3138;
	wire w3139;
	wire w3140;
	wire w3141;
	wire w3142;
	wire w3143;
	wire w3144;
	wire w3145;
	wire w3146;
	wire w3147;
	wire w3148;
	wire w3149;
	wire w3150;
	wire w3151;
	wire w3152;
	wire w3153;
	wire w3154;
	wire w3155;
	wire w3156;
	wire w3157;
	wire w3158;
	wire w3159;
	wire w3160;
	wire w3161;
	wire w3162;
	wire w3163;
	wire w3164;
	wire w3165;
	wire w3166;
	wire w3167;
	wire w3168;
	wire w3169;
	wire w3170;
	wire w3171;
	wire w3172;
	wire w3173;
	wire w3174;
	wire w3175;
	wire w3176;
	wire w3177;
	wire w3178;
	wire w3179;
	wire w3180;
	wire w3181;
	wire w3182;
	wire w3183;
	wire w3184;
	wire w3185;
	wire w3186;
	wire w3187;
	wire w3188;
	wire w3189;
	wire w3190;
	wire w3191;
	wire w3192;
	wire w3193;
	wire w3194;
	wire w3195;
	wire w3196;
	wire w3197;
	wire w3198;
	wire w3199;
	wire w3200;
	wire w3201;
	wire w3202;
	wire w3203;
	wire w3204;
	wire w3205;
	wire w3206;
	wire w3207;
	wire w3208;
	wire w3209;
	wire w3210;
	wire w3211;
	wire w3212;
	wire w3213;
	wire w3214;
	wire w3215;
	wire w3216;
	wire w3217;
	wire w3218;
	wire w3219;
	wire w3220;
	wire w3221;
	wire w3222;
	wire w3223;
	wire w3224;
	wire w3225;
	wire w3226;
	wire w3227;
	wire w3228;
	wire w3229;
	wire w3230;
	wire w3231;
	wire w3232;
	wire w3233;
	wire w3234;
	wire w3235;
	wire w3236;
	wire w3237;
	wire w3238;
	wire w3239;
	wire w3240;
	wire w3241;
	wire w3242;
	wire w3243;
	wire w3244;
	wire w3245;
	wire w3246;
	wire w3247;
	wire w3248;
	wire w3249;
	wire w3250;
	wire w3251;
	wire w3252;
	wire w3253;
	wire w3254;
	wire w3255;
	wire w3256;
	wire w3257;
	wire w3258;
	wire w3259;
	wire w3260;
	wire w3261;
	wire w3262;
	wire w3263;
	wire w3264;
	wire w3265;
	wire w3266;
	wire w3267;
	wire w3268;
	wire w3269;
	wire w3270;
	wire w3271;
	wire w3272;
	wire w3273;
	wire w3274;
	wire w3275;
	wire w3276;
	wire w3277;
	wire w3278;
	wire w3279;
	wire w3280;
	wire w3281;
	wire w3282;
	wire w3283;
	wire w3284;
	wire w3285;
	wire w3286;
	wire w3287;
	wire w3288;
	wire w3289;
	wire w3290;
	wire w3291;
	wire w3292;
	wire w3293;
	wire w3294;
	wire w3295;
	wire w3296;
	wire w3297;
	wire w3298;
	wire w3299;
	wire w3300;
	wire w3301;
	wire w3302;
	wire w3303;
	wire w3304;
	wire w3305;
	wire w3306;
	wire w3307;
	wire w3308;
	wire w3309;
	wire w3310;
	wire w3311;
	wire w3312;
	wire w3313;
	wire w3314;
	wire w3315;
	wire w3316;
	wire w3317;
	wire w3318;
	wire w3319;
	wire w3320;
	wire w3321;
	wire w3322;
	wire w3323;
	wire w3324;
	wire w3325;
	wire w3326;
	wire w3327;
	wire w3328;
	wire w3329;
	wire w3330;
	wire w3331;
	wire w3332;
	wire w3333;
	wire w3334;
	wire w3335;
	wire w3336;
	wire w3337;
	wire w3338;
	wire w3339;
	wire w3340;
	wire w3341;
	wire w3342;
	wire w3343;
	wire w3344;
	wire w3345;
	wire w3346;
	wire w3347;
	wire w3348;
	wire w3349;
	wire w3350;
	wire w3351;
	wire w3352;
	wire w3353;
	wire w3354;
	wire w3355;
	wire w3356;
	wire w3357;
	wire w3358;
	wire w3359;
	wire w3360;
	wire w3361;
	wire w3362;
	wire w3363;
	wire w3364;
	wire w3365;
	wire w3366;
	wire w3367;
	wire w3368;
	wire w3369;
	wire w3370;
	wire w3371;
	wire w3372;
	wire w3373;
	wire w3374;
	wire w3375;
	wire w3376;
	wire w3377;
	wire w3378;
	wire w3379;
	wire w3380;
	wire w3381;
	wire w3382;
	wire w3383;
	wire w3384;
	wire w3385;
	wire w3386;
	wire w3387;
	wire w3388;
	wire w3389;
	wire w3390;
	wire w3391;
	wire w3392;
	wire w3393;
	wire w3394;
	wire w3395;
	wire w3396;
	wire w3397;
	wire w3398;
	wire w3399;
	wire w3400;
	wire w3401;
	wire w3402;
	wire w3403;
	wire w3404;
	wire w3405;
	wire w3406;
	wire w3407;
	wire w3408;
	wire w3409;
	wire w3410;
	wire w3411;
	wire w3412;
	wire w3413;
	wire w3414;
	wire w3415;
	wire w3416;
	wire w3417;
	wire w3418;
	wire w3419;
	wire w3420;
	wire w3421;
	wire w3422;
	wire w3423;
	wire w3424;
	wire w3425;
	wire w3426;
	wire w3427;
	wire w3428;
	wire w3429;
	wire w3430;
	wire w3431;
	wire w3432;
	wire w3433;
	wire w3434;
	wire w3435;
	wire w3436;
	wire w3437;
	wire w3438;
	wire w3439;
	wire w3440;
	wire w3441;
	wire w3442;
	wire w3443;
	wire w3444;
	wire w3445;
	wire w3446;
	wire w3447;
	wire w3448;
	wire w3449;
	wire w3450;
	wire w3451;
	wire w3452;
	wire w3453;
	wire w3454;
	wire w3455;
	wire w3456;
	wire w3457;
	wire w3458;
	wire w3459;
	wire w3460;
	wire w3461;
	wire w3462;
	wire w3463;
	wire w3464;
	wire w3465;
	wire w3466;
	wire w3467;
	wire w3468;
	wire w3469;
	wire w3470;
	wire w3471;
	wire w3472;
	wire w3473;
	wire w3474;
	wire w3475;
	wire w3476;
	wire w3477;
	wire w3478;
	wire w3479;
	wire w3480;
	wire w3481;
	wire w3482;
	wire w3483;
	wire w3484;
	wire w3485;
	wire w3486;
	wire w3487;
	wire w3488;
	wire w3489;
	wire w3490;
	wire w3491;
	wire w3492;
	wire w3493;
	wire w3494;
	wire w3495;
	wire w3496;
	wire w3497;
	wire w3498;
	wire w3499;
	wire w3500;
	wire w3501;
	wire w3502;
	wire w3503;
	wire w3504;
	wire w3505;
	wire w3506;
	wire w3507;
	wire w3508;
	wire w3509;
	wire w3510;
	wire w3511;
	wire w3512;
	wire w3513;
	wire w3514;
	wire w3515;
	wire w3516;
	wire w3517;
	wire w3518;
	wire w3519;
	wire w3520;
	wire w3521;
	wire w3522;
	wire w3523;
	wire w3524;
	wire w3525;
	wire w3526;
	wire w3527;
	wire w3528;
	wire w3529;
	wire w3530;
	wire w3531;
	wire w3532;
	wire w3533;
	wire w3534;
	wire w3535;
	wire w3536;
	wire w3537;
	wire w3538;
	wire w3539;
	wire w3540;
	wire w3541;
	wire w3542;
	wire w3543;
	wire w3544;
	wire w3545;
	wire w3546;
	wire w3547;
	wire w3548;
	wire w3549;
	wire w3550;
	wire w3551;
	wire w3552;
	wire w3553;
	wire w3554;
	wire w3555;
	wire w3556;
	wire w3557;
	wire w3558;
	wire w3559;
	wire w3560;
	wire w3561;
	wire w3562;
	wire w3563;
	wire w3564;
	wire w3565;
	wire w3566;
	wire w3567;
	wire w3568;
	wire w3569;
	wire w3570;
	wire w3571;
	wire w3572;
	wire w3573;
	wire w3574;
	wire w3575;
	wire w3576;
	wire w3577;
	wire w3578;
	wire w3579;
	wire w3580;
	wire w3581;
	wire w3582;
	wire w3583;
	wire w3584;
	wire w3585;
	wire w3586;
	wire w3587;
	wire w3588;
	wire w3589;
	wire w3590;
	wire w3591;
	wire w3592;
	wire w3593;
	wire w3594;
	wire w3595;
	wire w3596;
	wire w3597;
	wire w3598;
	wire w3599;
	wire w3600;
	wire w3601;
	wire w3602;
	wire w3603;
	wire w3604;
	wire w3605;
	wire w3606;
	wire w3607;
	wire w3608;
	wire w3609;
	wire w3610;
	wire w3611;
	wire w3612;
	wire w3613;
	wire w3614;
	wire w3615;
	wire w3616;
	wire w3617;
	wire w3618;
	wire w3619;
	wire w3620;
	wire w3621;
	wire w3622;
	wire w3623;
	wire w3624;
	wire w3625;
	wire w3626;
	wire w3627;
	wire w3628;
	wire w3629;
	wire w3630;
	wire w3631;
	wire w3632;
	wire w3633;
	wire w3634;
	wire w3635;
	wire w3636;
	wire w3637;
	wire w3638;
	wire w3639;
	wire w3640;
	wire w3641;
	wire w3642;
	wire w3643;
	wire w3644;
	wire w3645;
	wire w3646;
	wire w3647;
	wire w3648;
	wire w3649;
	wire w3650;
	wire w3651;
	wire w3652;
	wire w3653;
	wire w3654;
	wire w3655;
	wire w3656;
	wire w3657;
	wire w3658;
	wire w3659;
	wire w3660;
	wire w3661;
	wire w3662;
	wire w3663;
	wire w3664;
	wire w3665;
	wire w3666;
	wire w3667;
	wire w3668;
	wire w3669;
	wire w3670;
	wire w3671;
	wire w3672;
	wire w3673;
	wire w3674;
	wire w3675;
	wire w3676;
	wire w3677;
	wire w3678;
	wire w3679;
	wire w3680;
	wire w3681;
	wire w3682;
	wire w3683;
	wire w3684;
	wire w3685;
	wire w3686;
	wire w3687;
	wire w3688;
	wire w3689;
	wire w3690;
	wire w3691;
	wire w3692;
	wire w3693;
	wire w3694;
	wire w3695;
	wire w3696;
	wire w3697;
	wire w3698;
	wire w3699;
	wire w3700;
	wire w3701;
	wire w3702;
	wire w3703;
	wire w3704;
	wire w3705;
	wire w3706;
	wire w3707;
	wire w3708;
	wire w3709;
	wire w3710;
	wire w3711;
	wire w3712;
	wire w3713;
	wire w3714;
	wire w3715;
	wire w3716;
	wire w3717;
	wire w3718;
	wire w3719;
	wire w3720;
	wire w3721;
	wire w3722;
	wire w3723;
	wire w3724;
	wire w3725;
	wire w3726;
	wire w3727;
	wire w3728;
	wire w3729;
	wire w3730;
	wire w3731;
	wire w3732;
	wire w3733;
	wire w3734;
	wire w3735;
	wire w3736;
	wire w3737;
	wire w3738;
	wire w3739;
	wire w3740;
	wire w3741;
	wire w3742;
	wire w3743;
	wire w3744;
	wire w3745;
	wire w3746;
	wire w3747;
	wire w3748;
	wire w3749;
	wire w3750;
	wire w3751;
	wire w3752;
	wire w3753;
	wire w3754;
	wire w3755;
	wire w3756;
	wire w3757;
	wire w3758;
	wire w3759;
	wire w3760;
	wire w3761;
	wire w3762;
	wire w3763;
	wire w3764;
	wire w3765;
	wire w3766;
	wire w3767;
	wire w3768;
	wire w3769;
	wire w3770;
	wire w3771;
	wire w3772;
	wire w3773;
	wire w3774;
	wire w3775;
	wire w3776;
	wire w3777;
	wire w3778;
	wire w3779;
	wire w3780;
	wire w3781;
	wire w3782;
	wire w3783;
	wire w3784;
	wire w3785;
	wire w3786;
	wire w3787;
	wire w3788;
	wire w3789;
	wire w3790;
	wire w3791;
	wire w3792;
	wire w3793;
	wire w3794;
	wire w3795;
	wire w3796;
	wire w3797;
	wire w3798;
	wire w3799;
	wire w3800;
	wire w3801;
	wire w3802;
	wire w3803;
	wire w3804;
	wire w3805;
	wire w3806;
	wire w3807;
	wire w3808;
	wire w3809;
	wire w3810;
	wire w3811;
	wire w3812;
	wire w3813;
	wire w3814;
	wire w3815;
	wire w3816;
	wire w3817;
	wire w3818;
	wire w3819;
	wire w3820;
	wire w3821;
	wire w3822;
	wire w3823;
	wire w3824;
	wire w3825;
	wire w3826;
	wire w3827;
	wire w3828;
	wire w3829;
	wire w3830;
	wire w3831;
	wire w3832;
	wire w3833;
	wire w3834;
	wire w3835;
	wire w3836;
	wire w3837;
	wire w3838;
	wire w3839;
	wire w3840;
	wire w3841;
	wire w3842;
	wire w3843;
	wire w3844;
	wire w3845;
	wire w3846;
	wire w3847;
	wire w3848;
	wire w3849;
	wire w3850;
	wire w3851;
	wire w3852;
	wire w3853;
	wire w3854;
	wire w3855;
	wire w3856;
	wire w3857;
	wire w3858;
	wire w3859;
	wire w3860;
	wire w3861;
	wire w3862;
	wire w3863;
	wire w3864;
	wire w3865;
	wire w3866;
	wire w3867;
	wire w3868;
	wire w3869;
	wire w3870;
	wire w3871;
	wire w3872;
	wire w3873;
	wire w3874;
	wire w3875;
	wire w3876;
	wire w3877;
	wire w3878;
	wire w3879;
	wire w3880;
	wire w3881;
	wire w3882;
	wire w3883;
	wire w3884;
	wire w3885;
	wire w3886;
	wire w3887;
	wire w3888;
	wire w3889;
	wire w3890;
	wire w3891;
	wire w3892;
	wire w3893;
	wire w3894;
	wire w3895;
	wire w3896;
	wire w3897;
	wire w3898;
	wire w3899;
	wire w3900;
	wire w3901;
	wire w3902;
	wire w3903;
	wire w3904;
	wire w3905;
	wire w3906;
	wire w3907;
	wire w3908;
	wire w3909;
	wire w3910;
	wire w3911;
	wire w3912;
	wire w3913;
	wire w3914;
	wire w3915;
	wire w3916;
	wire w3917;
	wire w3918;
	wire w3919;
	wire w3920;
	wire w3921;
	wire w3922;
	wire w3923;
	wire w3924;
	wire w3925;
	wire w3926;
	wire w3927;
	wire w3928;
	wire w3929;
	wire w3930;
	wire w3931;
	wire w3932;
	wire w3933;
	wire w3934;
	wire w3935;
	wire w3936;
	wire w3937;
	wire w3938;
	wire w3939;
	wire w3940;
	wire w3941;
	wire w3942;
	wire w3943;
	wire w3944;
	wire w3945;
	wire w3946;
	wire w3947;
	wire w3948;
	wire w3949;
	wire w3950;
	wire w3951;
	wire w3952;
	wire w3953;
	wire w3954;
	wire w3955;
	wire w3956;
	wire w3957;
	wire w3958;
	wire w3959;
	wire w3960;
	wire w3961;
	wire w3962;
	wire w3963;
	wire w3964;
	wire w3965;
	wire w3966;
	wire w3967;
	wire w3968;
	wire w3969;
	wire w3970;
	wire w3971;
	wire w3972;
	wire w3973;
	wire w3974;
	wire w3975;
	wire w3976;
	wire w3977;
	wire w3978;
	wire w3979;
	wire w3980;
	wire w3981;
	wire w3982;
	wire w3983;
	wire w3984;
	wire w3985;
	wire w3986;
	wire w3987;
	wire w3988;
	wire w3989;
	wire w3990;
	wire w3991;
	wire w3992;
	wire w3993;
	wire w3994;
	wire w3995;
	wire w3996;
	wire w3997;
	wire w3998;
	wire w3999;
	wire w4000;
	wire w4001;
	wire w4002;
	wire w4003;
	wire w4004;
	wire w4005;
	wire w4006;
	wire w4007;
	wire w4008;
	wire w4009;
	wire w4010;
	wire w4011;
	wire w4012;
	wire w4013;
	wire w4014;
	wire w4015;
	wire w4016;
	wire w4017;
	wire w4018;
	wire w4019;
	wire w4020;
	wire w4021;
	wire w4022;
	wire w4023;
	wire w4024;
	wire w4025;
	wire w4026;
	wire w4027;
	wire w4028;
	wire w4029;
	wire w4030;
	wire w4031;
	wire w4032;
	wire w4033;
	wire w4034;
	wire w4035;
	wire w4036;
	wire w4037;
	wire w4038;
	wire w4039;
	wire w4040;
	wire w4041;
	wire w4042;
	wire w4043;
	wire w4044;
	wire w4045;
	wire w4046;
	wire w4047;
	wire w4048;
	wire w4049;
	wire w4050;
	wire w4051;
	wire w4052;
	wire w4053;
	wire w4054;
	wire w4055;
	wire w4056;
	wire w4057;
	wire w4058;
	wire w4059;
	wire w4060;
	wire w4061;
	wire w4062;
	wire w4063;
	wire w4064;
	wire w4065;
	wire w4066;
	wire w4067;
	wire w4068;
	wire w4069;
	wire w4070;
	wire w4071;
	wire w4072;
	wire w4073;
	wire w4074;
	wire w4075;
	wire w4076;
	wire w4077;
	wire w4078;
	wire w4079;
	wire w4080;
	wire w4081;
	wire w4082;
	wire w4083;
	wire w4084;
	wire w4085;
	wire w4086;
	wire w4087;
	wire w4088;
	wire w4089;
	wire w4090;
	wire w4091;
	wire w4092;
	wire w4093;
	wire w4094;
	wire w4095;
	wire w4096;
	wire w4097;
	wire w4098;
	wire w4099;
	wire w4100;
	wire w4101;
	wire w4102;
	wire w4103;
	wire w4104;
	wire w4105;
	wire w4106;
	wire w4107;
	wire w4108;
	wire w4109;
	wire w4110;
	wire w4111;
	wire w4112;
	wire w4113;
	wire w4114;
	wire w4115;
	wire w4116;
	wire w4117;
	wire w4118;
	wire w4119;
	wire w4120;
	wire w4121;
	wire w4122;
	wire w4123;
	wire w4124;
	wire w4125;
	wire w4126;
	wire w4127;
	wire w4128;
	wire w4129;
	wire w4130;
	wire w4131;
	wire w4132;
	wire w4133;
	wire w4134;
	wire w4135;
	wire w4136;
	wire w4137;
	wire w4138;
	wire w4139;
	wire w4140;
	wire w4141;
	wire w4142;
	wire w4143;
	wire w4144;
	wire w4145;
	wire w4146;
	wire w4147;
	wire w4148;
	wire w4149;
	wire w4150;
	wire w4151;
	wire w4152;
	wire w4153;
	wire w4154;
	wire w4155;
	wire w4156;
	wire w4157;
	wire w4158;
	wire w4159;
	wire w4160;
	wire w4161;
	wire w4162;
	wire w4163;
	wire w4164;
	wire w4165;
	wire w4166;
	wire w4167;
	wire w4168;
	wire w4169;
	wire w4170;
	wire w4171;
	wire w4172;
	wire w4173;
	wire w4174;
	wire w4175;
	wire w4176;
	wire w4177;
	wire w4178;
	wire w4179;
	wire w4180;
	wire w4181;
	wire w4182;
	wire w4183;
	wire w4184;
	wire w4185;
	wire w4186;
	wire w4187;
	wire w4188;
	wire w4189;
	wire w4190;
	wire w4191;
	wire w4192;
	wire w4193;
	wire w4194;
	wire w4195;
	wire w4196;
	wire w4197;
	wire w4198;
	wire w4199;
	wire w4200;
	wire w4201;
	wire w4202;
	wire w4203;
	wire w4204;
	wire w4205;
	wire w4206;
	wire w4207;
	wire w4208;
	wire w4209;
	wire w4210;
	wire w4211;
	wire w4212;
	wire w4213;
	wire w4214;
	wire w4215;
	wire w4216;
	wire w4217;
	wire w4218;
	wire w4219;
	wire w4220;
	wire w4221;
	wire w4222;
	wire w4223;
	wire w4224;
	wire w4225;
	wire w4226;
	wire w4227;
	wire w4228;
	wire w4229;
	wire w4230;
	wire w4231;
	wire w4232;
	wire w4233;
	wire w4234;
	wire w4235;
	wire w4236;
	wire w4237;
	wire w4238;
	wire w4239;
	wire w4240;
	wire w4241;
	wire w4242;
	wire w4243;
	wire w4244;
	wire w4245;
	wire w4246;
	wire w4247;
	wire w4248;
	wire w4249;
	wire w4250;
	wire w4251;
	wire w4252;
	wire w4253;
	wire w4254;
	wire w4255;
	wire w4256;
	wire w4257;
	wire w4258;
	wire w4259;
	wire w4260;
	wire w4261;
	wire w4262;
	wire w4263;
	wire w4264;
	wire w4265;
	wire w4266;
	wire w4267;
	wire w4268;
	wire w4269;
	wire w4270;
	wire w4271;
	wire w4272;
	wire w4273;
	wire w4274;
	wire w4275;
	wire w4276;
	wire w4277;
	wire w4278;
	wire w4279;
	wire w4280;
	wire w4281;
	wire w4282;
	wire w4283;
	wire w4284;
	wire w4285;
	wire w4286;
	wire w4287;
	wire w4288;
	wire w4289;
	wire w4290;
	wire w4291;
	wire w4292;
	wire w4293;
	wire w4294;
	wire w4295;
	wire w4296;
	wire w4297;
	wire w4298;
	wire w4299;
	wire w4300;
	wire w4301;
	wire w4302;
	wire w4303;
	wire w4304;
	wire w4305;
	wire w4306;
	wire w4307;
	wire w4308;
	wire w4309;
	wire w4310;
	wire w4311;
	wire w4312;
	wire w4313;
	wire w4314;
	wire w4315;
	wire w4316;
	wire w4317;
	wire w4318;
	wire w4319;
	wire w4320;
	wire w4321;
	wire w4322;
	wire w4323;
	wire w4324;
	wire w4325;
	wire w4326;
	wire w4327;
	wire w4328;
	wire w4329;
	wire w4330;
	wire w4331;
	wire w4332;
	wire w4333;
	wire w4334;
	wire w4335;
	wire w4336;
	wire w4337;
	wire w4338;
	wire w4339;
	wire w4340;
	wire w4341;
	wire w4342;
	wire w4343;
	wire w4344;
	wire w4345;
	wire w4346;
	wire w4347;
	wire w4348;
	wire w4349;
	wire w4350;
	wire w4351;
	wire w4352;
	wire w4353;
	wire w4354;
	wire w4355;
	wire w4356;
	wire w4357;
	wire w4358;
	wire w4359;
	wire w4360;
	wire w4361;
	wire w4362;
	wire w4363;
	wire w4364;
	wire w4365;
	wire w4366;
	wire w4367;
	wire w4368;
	wire w4369;
	wire w4370;
	wire w4371;
	wire w4372;
	wire w4373;
	wire w4374;
	wire w4375;
	wire w4376;
	wire w4377;
	wire w4378;
	wire w4379;
	wire w4380;
	wire w4381;
	wire w4382;
	wire w4383;
	wire w4384;
	wire w4385;
	wire w4386;
	wire w4387;
	wire w4388;
	wire w4389;
	wire w4390;
	wire w4391;
	wire w4392;
	wire w4393;
	wire w4394;
	wire w4395;
	wire w4396;
	wire w4397;
	wire w4398;
	wire w4399;
	wire w4400;
	wire w4401;
	wire w4402;
	wire w4403;
	wire w4404;
	wire w4405;
	wire w4406;
	wire w4407;
	wire w4408;
	wire w4409;
	wire w4410;
	wire w4411;
	wire w4412;
	wire w4413;
	wire w4414;
	wire w4415;
	wire w4416;
	wire w4417;
	wire w4418;
	wire w4419;
	wire w4420;
	wire w4421;
	wire w4422;
	wire w4423;
	wire w4424;
	wire w4425;
	wire w4426;
	wire w4427;
	wire w4428;
	wire w4429;
	wire w4430;
	wire w4431;
	wire w4432;
	wire w4433;
	wire w4434;
	wire w4435;
	wire w4436;
	wire w4437;
	wire w4438;
	wire w4439;
	wire w4440;
	wire w4441;
	wire w4442;
	wire w4443;
	wire w4444;
	wire w4445;
	wire w4446;
	wire w4447;
	wire w4448;
	wire w4449;
	wire w4450;
	wire w4451;
	wire 68K CPU CLOCK;
	wire w4453;
	wire w4454;
	wire w4455;
	wire w4456;
	wire w4457;
	wire w4458;
	wire w4459;
	wire w4460;
	wire w4461;
	wire w4462;
	wire w4463;
	wire w4464;
	wire w4465;
	wire w4466;
	wire w4467;
	wire w4468;
	wire w4469;
	wire w4470;
	wire w4471;
	wire w4472;
	wire w4473;
	wire w4474;
	wire w4475;
	wire w4476;
	wire w4477;
	wire w4478;
	wire w4479;
	wire w4480;
	wire w4481;
	wire w4482;
	wire w4483;
	wire w4484;
	wire w4485;
	wire w4486;
	wire w4487;
	wire w4488;
	wire w4489;
	wire w4490;
	wire w4491;
	wire w4492;
	wire w4493;
	wire w4494;
	wire w4495;
	wire w4496;
	wire nRAS1;
	wire nCAS1;
	wire nWE1;
	wire nWE0;
	wire nOE1;
	wire AD_RD_DIR;
	wire w4503;
	wire w4504;
	wire w4505;
	wire w4506;
	wire w4507;
	wire w4508;
	wire w4509;
	wire w4510;
	wire w4511;
	wire w4512;
	wire w4513;
	wire w4514;
	wire w4515;
	wire w4516;
	wire w4517;
	wire w4518;
	wire w4519;
	wire w4520;
	wire w4521;
	wire w4522;
	wire w4523;
	wire w4524;
	wire w4525;
	wire w4526;
	wire w4527;
	wire w4528;
	wire w4529;
	wire w4530;
	wire w4531;
	wire w4532;
	wire w4533;
	wire w4534;
	wire w4535;
	wire w4536;
	wire w4537;
	wire w4538;
	wire w4539;
	wire w4540;
	wire w4541;
	wire w4542;
	wire w4543;
	wire w4544;
	wire w4545;
	wire w4546;
	wire w4547;
	wire w4548;
	wire w4549;
	wire w4550;
	wire w4551;
	wire w4552;
	wire w4553;
	wire w4554;
	wire w4555;
	wire w4556;
	wire w4557;
	wire w4558;
	wire w4559;
	wire w4560;
	wire w4561;
	wire w4562;
	wire w4563;
	wire w4564;
	wire w4565;
	wire w4566;
	wire w4567;
	wire w4568;
	wire w4569;
	wire w4570;
	wire w4571;
	wire w4572;
	wire w4573;
	wire w4574;
	wire w4575;
	wire w4576;
	wire w4577;
	wire w4578;
	wire w4579;
	wire w4580;
	wire w4581;
	wire w4582;
	wire w4583;
	wire w4584;
	wire w4585;
	wire w4586;
	wire w4587;
	wire w4588;
	wire w4589;
	wire w4590;
	wire w4591;
	wire w4592;
	wire w4593;
	wire w4594;
	wire w4595;
	wire w4596;
	wire w4597;
	wire w4598;
	wire w4599;
	wire w4600;
	wire w4601;
	wire w4602;
	wire w4603;
	wire w4604;
	wire w4605;
	wire w4606;
	wire w4607;
	wire w4608;
	wire w4609;
	wire w4610;
	wire w4611;
	wire w4612;
	wire w4613;
	wire w4614;
	wire w4615;
	wire w4616;
	wire w4617;
	wire w4618;
	wire w4619;
	wire w4620;
	wire w4621;
	wire w4622;
	wire w4623;
	wire w4624;
	wire w4625;
	wire w4626;
	wire w4627;
	wire w4628;
	wire w4629;
	wire w4630;
	wire w4631;
	wire w4632;
	wire w4633;
	wire w4634;
	wire w4635;
	wire w4636;
	wire w4637;
	wire w4638;
	wire w4639;
	wire w4640;
	wire w4641;
	wire w4642;
	wire w4643;
	wire w4644;
	wire w4645;
	wire w4646;
	wire w4647;
	wire w4648;
	wire w4649;
	wire w4650;
	wire w4651;
	wire w4652;
	wire w4653;
	wire w4654;
	wire w4655;
	wire w4656;
	wire w4657;
	wire w4658;
	wire w4659;
	wire w4660;
	wire w4661;
	wire w4662;
	wire w4663;
	wire w4664;
	wire w4665;
	wire w4666;
	wire w4667;
	wire w4668;
	wire w4669;
	wire w4670;
	wire w4671;
	wire w4672;
	wire w4673;
	wire w4674;
	wire w4675;
	wire w4676;
	wire w4677;
	wire w4678;
	wire w4679;
	wire w4680;
	wire w4681;
	wire w4682;
	wire w4683;
	wire w4684;
	wire w4685;
	wire w4686;
	wire w4687;
	wire w4688;
	wire w4689;
	wire w4690;
	wire w4691;
	wire w4692;
	wire w4693;
	wire w4694;
	wire w4695;
	wire w4696;
	wire w4697;
	wire w4698;
	wire w4699;
	wire w4700;
	wire w4701;
	wire w4702;
	wire w4703;
	wire w4704;
	wire w4705;
	wire w4706;
	wire w4707;
	wire w4708;
	wire w4709;
	wire w4710;
	wire w4711;
	wire w4712;
	wire w4713;
	wire w4714;
	wire w4715;
	wire w4716;
	wire w4717;
	wire w4718;
	wire w4719;
	wire w4720;
	wire w4721;
	wire w4722;
	wire w4723;
	wire w4724;
	wire w4725;
	wire w4726;
	wire w4727;
	wire w4728;
	wire w4729;
	wire w4730;
	wire w4731;
	wire w4732;
	wire w4733;
	wire w4734;
	wire w4735;
	wire w4736;
	wire w4737;
	wire w4738;
	wire w4739;
	wire w4740;
	wire w4741;
	wire w4742;
	wire w4743;
	wire w4744;
	wire w4745;
	wire w4746;
	wire w4747;
	wire w4748;
	wire w4749;
	wire w4750;
	wire w4751;
	wire w4752;
	wire w4753;
	wire w4754;
	wire w4755;
	wire w4756;
	wire w4757;
	wire w4758;
	wire w4759;
	wire w4760;
	wire w4761;
	wire w4762;
	wire w4763;
	wire w4764;
	wire w4765;
	wire w4766;
	wire w4767;
	wire w4768;
	wire w4769;
	wire w4770;
	wire w4771;
	wire w4772;
	wire w4773;
	wire w4774;
	wire w4775;
	wire w4776;
	wire w4777;
	wire w4778;
	wire w4779;
	wire w4780;
	wire w4781;
	wire w4782;
	wire w4783;
	wire w4784;
	wire w4785;
	wire w4786;
	wire w4787;
	wire w4788;
	wire w4789;
	wire w4790;
	wire w4791;
	wire w4792;
	wire w4793;
	wire w4794;
	wire w4795;
	wire w4796;
	wire w4797;
	wire w4798;
	wire w4799;
	wire w4800;
	wire w4801;
	wire w4802;
	wire w4803;
	wire w4804;
	wire w4805;
	wire w4806;
	wire w4807;
	wire w4808;
	wire w4809;
	wire w4810;
	wire w4811;
	wire w4812;
	wire w4813;
	wire w4814;
	wire w4815;
	wire w4816;
	wire w4817;
	wire w4818;
	wire w4819;
	wire w4820;
	wire w4821;
	wire w4822;
	wire w4823;
	wire w4824;
	wire w4825;
	wire w4826;
	wire w4827;
	wire w4828;
	wire w4829;
	wire w4830;
	wire w4831;
	wire w4832;
	wire w4833;
	wire w4834;
	wire w4835;
	wire w4836;
	wire w4837;
	wire w4838;
	wire w4839;
	wire w4840;
	wire w4841;
	wire w4842;
	wire w4843;
	wire w4844;
	wire w4845;
	wire w4846;
	wire w4847;
	wire w4848;
	wire w4849;
	wire w4850;
	wire w4851;
	wire w4852;
	wire w4853;
	wire w4854;
	wire w4855;
	wire w4856;
	wire w4857;
	wire w4858;
	wire w4859;
	wire w4860;
	wire w4861;
	wire w4862;
	wire w4863;
	wire w4864;
	wire w4865;
	wire w4866;
	wire w4867;
	wire w4868;
	wire w4869;
	wire w4870;
	wire w4871;
	wire w4872;
	wire w4873;
	wire w4874;
	wire w4875;
	wire w4876;
	wire w4877;
	wire w4878;
	wire w4879;
	wire w4880;
	wire w4881;
	wire w4882;
	wire w4883;
	wire w4884;
	wire w4885;
	wire w4886;
	wire w4887;
	wire w4888;
	wire w4889;
	wire w4890;
	wire w4891;
	wire w4892;
	wire w4893;
	wire w4894;
	wire w4895;
	wire w4896;
	wire w4897;
	wire w4898;
	wire w4899;
	wire w4900;
	wire w4901;
	wire w4902;
	wire w4903;
	wire w4904;
	wire w4905;
	wire w4906;
	wire w4907;
	wire w4908;
	wire w4909;
	wire w4910;
	wire w4911;
	wire w4912;
	wire w4913;
	wire w4914;
	wire w4915;
	wire w4916;
	wire w4917;
	wire w4918;
	wire w4919;
	wire w4920;
	wire w4921;
	wire w4922;
	wire w4923;
	wire w4924;
	wire w4925;
	wire w4926;
	wire w4927;
	wire w4928;
	wire w4929;
	wire w4930;
	wire w4931;
	wire w4932;
	wire w4933;
	wire w4934;
	wire w4935;
	wire w4936;
	wire w4937;
	wire w4938;
	wire w4939;
	wire w4940;
	wire w4941;
	wire w4942;
	wire w4943;
	wire w4944;
	wire w4945;
	wire w4946;
	wire w4947;
	wire w4948;
	wire w4949;
	wire w4950;
	wire w4951;
	wire w4952;
	wire w4953;
	wire w4954;
	wire w4955;
	wire w4956;
	wire w4957;
	wire w4958;
	wire w4959;
	wire w4960;
	wire w4961;
	wire w4962;
	wire w4963;
	wire w4964;
	wire w4965;
	wire w4966;
	wire w4967;
	wire w4968;
	wire w4969;
	wire w4970;
	wire w4971;
	wire w4972;
	wire w4973;
	wire w4974;
	wire w4975;
	wire w4976;
	wire w4977;
	wire w4978;
	wire w4979;
	wire w4980;
	wire w4981;
	wire w4982;
	wire w4983;
	wire w4984;
	wire w4985;
	wire w4986;
	wire w4987;
	wire w4988;
	wire w4989;
	wire w4990;
	wire w4991;
	wire w4992;
	wire w4993;
	wire w4994;
	wire w4995;
	wire w4996;
	wire w4997;
	wire w4998;
	wire w4999;
	wire w5000;
	wire w5001;
	wire w5002;
	wire w5003;
	wire w5004;
	wire w5005;
	wire w5006;
	wire w5007;
	wire w5008;
	wire w5009;
	wire w5010;
	wire w5011;
	wire w5012;
	wire w5013;
	wire w5014;
	wire w5015;
	wire w5016;
	wire w5017;
	wire w5018;
	wire w5019;
	wire w5020;
	wire w5021;
	wire w5022;
	wire w5023;
	wire w5024;
	wire w5025;
	wire w5026;
	wire w5027;
	wire w5028;
	wire w5029;
	wire w5030;
	wire w5031;
	wire w5032;
	wire w5033;
	wire w5034;
	wire w5035;
	wire w5036;
	wire w5037;
	wire w5038;
	wire w5039;
	wire w5040;
	wire w5041;
	wire w5042;
	wire w5043;
	wire w5044;
	wire w5045;
	wire w5046;
	wire w5047;
	wire w5048;
	wire w5049;
	wire w5050;
	wire w5051;
	wire w5052;
	wire w5053;
	wire w5054;
	wire w5055;
	wire w5056;
	wire w5057;
	wire w5058;
	wire w5059;
	wire w5060;
	wire w5061;
	wire w5062;
	wire w5063;
	wire w5064;
	wire w5065;
	wire w5066;
	wire w5067;
	wire w5068;
	wire w5069;
	wire w5070;
	wire w5071;
	wire w5072;
	wire w5073;
	wire w5074;
	wire w5075;
	wire w5076;
	wire w5077;
	wire w5078;
	wire w5079;
	wire w5080;
	wire w5081;
	wire w5082;
	wire w5083;
	wire w5084;
	wire w5085;
	wire w5086;
	wire w5087;
	wire w5088;
	wire w5089;
	wire w5090;
	wire w5091;
	wire w5092;
	wire w5093;
	wire w5094;
	wire w5095;
	wire w5096;
	wire w5097;
	wire w5098;
	wire w5099;
	wire w5100;
	wire w5101;
	wire w5102;
	wire w5103;
	wire w5104;
	wire w5105;
	wire w5106;
	wire w5107;
	wire w5108;
	wire w5109;
	wire w5110;
	wire w5111;
	wire w5112;
	wire w5113;
	wire w5114;
	wire w5115;
	wire w5116;
	wire w5117;
	wire w5118;
	wire w5119;
	wire w5120;
	wire w5121;
	wire w5122;
	wire w5123;
	wire w5124;
	wire w5125;
	wire w5126;
	wire w5127;
	wire w5128;
	wire w5129;
	wire w5130;
	wire w5131;
	wire w5132;
	wire w5133;
	wire w5134;
	wire w5135;
	wire w5136;
	wire w5137;
	wire w5138;
	wire w5139;
	wire w5140;
	wire w5141;
	wire w5142;
	wire w5143;
	wire w5144;
	wire w5145;
	wire w5146;
	wire w5147;
	wire w5148;
	wire w5149;
	wire w5150;
	wire w5151;
	wire w5152;
	wire w5153;
	wire w5154;
	wire w5155;
	wire w5156;
	wire w5157;
	wire w5158;
	wire w5159;
	wire w5160;
	wire w5161;
	wire w5162;
	wire w5163;
	wire w5164;
	wire w5165;
	wire w5166;
	wire w5167;
	wire w5168;
	wire w5169;
	wire w5170;
	wire w5171;
	wire w5172;
	wire w5173;
	wire w5174;
	wire w5175;
	wire w5176;
	wire w5177;
	wire w5178;
	wire w5179;
	wire w5180;
	wire w5181;
	wire w5182;
	wire w5183;
	wire w5184;
	wire w5185;
	wire w5186;
	wire w5187;
	wire w5188;
	wire w5189;
	wire w5190;
	wire w5191;
	wire w5192;
	wire w5193;
	wire w5194;
	wire w5195;
	wire w5196;
	wire w5197;
	wire w5198;
	wire w5199;
	wire w5200;
	wire w5201;
	wire w5202;
	wire w5203;
	wire w5204;
	wire w5205;
	wire w5206;
	wire w5207;
	wire w5208;
	wire w5209;
	wire w5210;
	wire w5211;
	wire w5212;
	wire w5213;
	wire w5214;
	wire w5215;
	wire w5216;
	wire w5217;
	wire w5218;
	wire w5219;
	wire w5220;
	wire w5221;
	wire w5222;
	wire w5223;
	wire w5224;
	wire w5225;
	wire w5226;
	wire w5227;
	wire w5228;
	wire w5229;
	wire w5230;
	wire w5231;
	wire w5232;
	wire w5233;
	wire w5234;
	wire w5235;
	wire w5236;
	wire w5237;
	wire w5238;
	wire w5239;
	wire w5240;
	wire w5241;
	wire w5242;
	wire w5243;
	wire w5244;
	wire w5245;
	wire w5246;
	wire w5247;
	wire w5248;
	wire w5249;
	wire w5250;
	wire w5251;
	wire w5252;
	wire w5253;
	wire w5254;
	wire w5255;
	wire w5256;
	wire w5257;
	wire w5258;
	wire w5259;
	wire w5260;
	wire w5261;
	wire w5262;
	wire w5263;
	wire w5264;
	wire w5265;
	wire w5266;
	wire w5267;
	wire w5268;
	wire w5269;
	wire w5270;
	wire w5271;
	wire w5272;
	wire w5273;
	wire w5274;
	wire w5275;
	wire w5276;
	wire w5277;
	wire w5278;
	wire w5279;
	wire w5280;
	wire w5281;
	wire w5282;
	wire w5283;
	wire w5284;
	wire w5285;
	wire w5286;
	wire w5287;
	wire w5288;
	wire w5289;
	wire w5290;
	wire w5291;
	wire w5292;
	wire w5293;
	wire w5294;
	wire w5295;
	wire w5296;
	wire w5297;
	wire w5298;
	wire w5299;
	wire w5300;
	wire w5301;
	wire w5302;
	wire w5303;
	wire w5304;
	wire w5305;
	wire w5306;
	wire w5307;
	wire w5308;
	wire w5309;
	wire w5310;
	wire w5311;
	wire w5312;
	wire w5313;
	wire w5314;
	wire w5315;
	wire w5316;
	wire w5317;
	wire w5318;
	wire w5319;
	wire w5320;
	wire w5321;
	wire w5322;
	wire w5323;
	wire w5324;
	wire w5325;
	wire w5326;
	wire w5327;
	wire w5328;
	wire w5329;
	wire w5330;
	wire w5331;
	wire w5332;
	wire w5333;
	wire w5334;
	wire w5335;
	wire w5336;
	wire w5337;
	wire w5338;
	wire w5339;
	wire w5340;
	wire w5341;
	wire w5342;
	wire w5343;
	wire w5344;
	wire w5345;
	wire w5346;
	wire w5347;
	wire w5348;
	wire w5349;
	wire w5350;
	wire w5351;
	wire w5352;
	wire w5353;
	wire w5354;
	wire w5355;
	wire w5356;
	wire w5357;
	wire w5358;
	wire w5359;
	wire w5360;
	wire w5361;
	wire w5362;
	wire w5363;
	wire w5364;
	wire w5365;
	wire w5366;
	wire w5367;
	wire w5368;
	wire w5369;
	wire w5370;
	wire w5371;
	wire w5372;
	wire w5373;
	wire w5374;
	wire w5375;
	wire w5376;
	wire w5377;
	wire w5378;
	wire w5379;
	wire w5380;
	wire w5381;
	wire w5382;
	wire w5383;
	wire w5384;
	wire w5385;
	wire w5386;
	wire w5387;
	wire w5388;
	wire w5389;
	wire w5390;
	wire w5391;
	wire w5392;
	wire w5393;
	wire w5394;
	wire w5395;
	wire w5396;
	wire w5397;
	wire w5398;
	wire w5399;
	wire w5400;
	wire w5401;
	wire w5402;
	wire w5403;
	wire w5404;
	wire w5405;
	wire w5406;
	wire w5407;
	wire w5408;
	wire w5409;
	wire w5410;
	wire w5411;
	wire w5412;
	wire w5413;
	wire w5414;
	wire w5415;
	wire w5416;
	wire w5417;
	wire w5418;
	wire w5419;
	wire w5420;
	wire w5421;
	wire w5422;
	wire w5423;
	wire w5424;
	wire w5425;
	wire w5426;
	wire w5427;
	wire w5428;
	wire w5429;
	wire w5430;
	wire w5431;
	wire w5432;
	wire w5433;
	wire w5434;
	wire w5435;
	wire w5436;
	wire w5437;
	wire w5438;
	wire w5439;
	wire w5440;
	wire w5441;
	wire w5442;
	wire w5443;
	wire w5444;
	wire w5445;
	wire w5446;
	wire w5447;
	wire w5448;
	wire w5449;
	wire w5450;
	wire w5451;
	wire w5452;
	wire w5453;
	wire w5454;
	wire w5455;
	wire w5456;
	wire w5457;
	wire w5458;
	wire w5459;
	wire w5460;
	wire w5461;
	wire w5462;
	wire w5463;
	wire w5464;
	wire w5465;
	wire w5466;
	wire w5467;
	wire w5468;
	wire w5469;
	wire w5470;
	wire w5471;
	wire w5472;
	wire w5473;
	wire w5474;
	wire w5475;
	wire w5476;
	wire w5477;
	wire w5478;
	wire w5479;
	wire w5480;
	wire w5481;
	wire w5482;
	wire w5483;
	wire w5484;
	wire w5485;
	wire w5486;
	wire w5487;
	wire w5488;
	wire w5489;
	wire w5490;
	wire w5491;
	wire w5492;
	wire w5493;
	wire w5494;
	wire w5495;
	wire w5496;
	wire w5497;
	wire w5498;
	wire w5499;
	wire w5500;
	wire w5501;
	wire w5502;
	wire w5503;
	wire w5504;
	wire w5505;
	wire w5506;
	wire w5507;
	wire w5508;
	wire w5509;
	wire w5510;
	wire w5511;
	wire w5512;
	wire w5513;
	wire w5514;
	wire w5515;
	wire w5516;
	wire w5517;
	wire w5518;
	wire w5519;
	wire w5520;
	wire w5521;
	wire w5522;
	wire w5523;
	wire w5524;
	wire w5525;
	wire w5526;
	wire w5527;
	wire w5528;
	wire w5529;
	wire w5530;
	wire w5531;
	wire w5532;
	wire w5533;
	wire w5534;
	wire w5535;
	wire w5536;
	wire w5537;
	wire w5538;
	wire w5539;
	wire w5540;
	wire w5541;
	wire w5542;
	wire w5543;
	wire w5544;
	wire w5545;
	wire w5546;
	wire w5547;
	wire w5548;
	wire w5549;
	wire w5550;
	wire w5551;
	wire w5552;
	wire w5553;
	wire w5554;
	wire w5555;
	wire w5556;
	wire w5557;
	wire w5558;
	wire w5559;
	wire w5560;
	wire w5561;
	wire w5562;
	wire w5563;
	wire w5564;
	wire w5565;
	wire w5566;
	wire w5567;
	wire w5568;
	wire w5569;
	wire w5570;
	wire w5571;
	wire w5572;
	wire w5573;
	wire w5574;
	wire w5575;
	wire w5576;
	wire w5577;
	wire w5578;
	wire w5579;
	wire w5580;
	wire w5581;
	wire w5582;
	wire w5583;
	wire w5584;
	wire w5585;
	wire w5586;
	wire w5587;
	wire w5588;
	wire w5589;
	wire w5590;
	wire w5591;
	wire w5592;
	wire w5593;
	wire w5594;
	wire w5595;
	wire w5596;
	wire w5597;
	wire w5598;
	wire w5599;
	wire w5600;
	wire w5601;
	wire w5602;
	wire w5603;
	wire w5604;
	wire w5605;
	wire w5606;
	wire w5607;
	wire w5608;
	wire w5609;
	wire w5610;
	wire w5611;
	wire w5612;
	wire w5613;
	wire w5614;
	wire w5615;
	wire w5616;
	wire w5617;
	wire w5618;
	wire w5619;
	wire w5620;
	wire w5621;
	wire w5622;
	wire w5623;
	wire w5624;
	wire w5625;
	wire w5626;
	wire w5627;
	wire w5628;
	wire w5629;
	wire w5630;
	wire w5631;
	wire w5632;
	wire w5633;
	wire w5634;
	wire w5635;
	wire w5636;
	wire w5637;
	wire w5638;
	wire w5639;
	wire w5640;
	wire w5641;
	wire w5642;
	wire w5643;
	wire w5644;
	wire w5645;
	wire w5646;
	wire w5647;
	wire w5648;
	wire w5649;
	wire w5650;
	wire w5651;
	wire w5652;
	wire w5653;
	wire w5654;
	wire w5655;
	wire w5656;
	wire w5657;
	wire w5658;
	wire w5659;
	wire w5660;
	wire w5661;
	wire w5662;
	wire w5663;
	wire w5664;
	wire w5665;
	wire w5666;
	wire w5667;
	wire w5668;
	wire w5669;
	wire w5670;
	wire w5671;
	wire w5672;
	wire w5673;
	wire w5674;
	wire w5675;
	wire w5676;
	wire w5677;
	wire w5678;
	wire w5679;
	wire w5680;
	wire w5681;
	wire w5682;
	wire w5683;
	wire w5684;
	wire w5685;
	wire w5686;
	wire w5687;
	wire w5688;
	wire w5689;
	wire w5690;
	wire w5691;
	wire w5692;
	wire w5693;
	wire w5694;
	wire w5695;
	wire w5696;
	wire w5697;
	wire w5698;
	wire w5699;
	wire w5700;
	wire w5701;
	wire w5702;
	wire w5703;
	wire w5704;
	wire w5705;
	wire w5706;
	wire w5707;
	wire w5708;
	wire w5709;
	wire w5710;
	wire w5711;
	wire w5712;
	wire w5713;
	wire w5714;
	wire w5715;
	wire w5716;
	wire w5717;
	wire w5718;
	wire w5719;
	wire w5720;
	wire w5721;
	wire w5722;
	wire w5723;
	wire w5724;
	wire w5725;
	wire w5726;
	wire w5727;
	wire w5728;
	wire w5729;
	wire w5730;
	wire w5731;
	wire w5732;
	wire w5733;
	wire w5734;
	wire w5735;
	wire w5736;
	wire w5737;
	wire w5738;
	wire w5739;
	wire w5740;
	wire w5741;
	wire w5742;
	wire w5743;
	wire w5744;
	wire w5745;
	wire w5746;
	wire w5747;
	wire w5748;
	wire w5749;
	wire w5750;
	wire w5751;
	wire w5752;
	wire w5753;
	wire w5754;
	wire w5755;
	wire w5756;
	wire w5757;
	wire w5758;
	wire w5759;
	wire w5760;
	wire w5761;
	wire w5762;
	wire w5763;
	wire w5764;
	wire w5765;
	wire w5766;
	wire w5767;
	wire w5768;
	wire w5769;
	wire w5770;
	wire w5771;
	wire w5772;
	wire w5773;
	wire w5774;
	wire w5775;
	wire w5776;
	wire w5777;
	wire w5778;
	wire w5779;
	wire w5780;
	wire w5781;
	wire w5782;
	wire w5783;
	wire w5784;
	wire w5785;
	wire w5786;
	wire w5787;
	wire w5788;
	wire w5789;
	wire w5790;
	wire w5791;
	wire w5792;
	wire w5793;
	wire w5794;
	wire w5795;
	wire w5796;
	wire w5797;
	wire w5798;
	wire w5799;
	wire w5800;
	wire w5801;
	wire w5802;
	wire w5803;
	wire w5804;
	wire w5805;
	wire w5806;
	wire w5807;
	wire w5808;
	wire w5809;
	wire w5810;
	wire w5811;
	wire w5812;
	wire w5813;
	wire w5814;
	wire w5815;
	wire w5816;
	wire w5817;
	wire w5818;
	wire w5819;
	wire w5820;
	wire w5821;
	wire w5822;
	wire w5823;
	wire w5824;
	wire w5825;
	wire w5826;
	wire w5827;
	wire w5828;
	wire w5829;
	wire w5830;
	wire w5831;
	wire w5832;
	wire w5833;
	wire w5834;
	wire w5835;
	wire w5836;
	wire w5837;
	wire w5838;
	wire w5839;
	wire w5840;
	wire w5841;
	wire w5842;
	wire w5843;
	wire w5844;
	wire w5845;
	wire w5846;
	wire w5847;
	wire w5848;
	wire w5849;
	wire w5850;
	wire w5851;
	wire w5852;
	wire w5853;
	wire w5854;
	wire w5855;
	wire w5856;
	wire w5857;
	wire w5858;
	wire w5859;
	wire w5860;
	wire w5861;
	wire w5862;
	wire w5863;
	wire w5864;
	wire w5865;
	wire w5866;
	wire w5867;
	wire w5868;
	wire w5869;
	wire w5870;
	wire w5871;
	wire w5872;
	wire w5873;
	wire w5874;
	wire w5875;
	wire w5876;
	wire w5877;
	wire w5878;
	wire w5879;
	wire w5880;
	wire w5881;
	wire w5882;
	wire w5883;
	wire w5884;
	wire w5885;
	wire w5886;
	wire w5887;
	wire w5888;
	wire w5889;
	wire w5890;
	wire w5891;
	wire w5892;
	wire w5893;
	wire w5894;
	wire w5895;
	wire w5896;
	wire w5897;
	wire w5898;
	wire w5899;
	wire w5900;
	wire w5901;
	wire w5902;
	wire w5903;
	wire w5904;
	wire w5905;
	wire w5906;
	wire w5907;
	wire w5908;
	wire w5909;
	wire w5910;
	wire w5911;
	wire w5912;
	wire w5913;
	wire w5914;
	wire w5915;
	wire w5916;
	wire w5917;
	wire w5918;
	wire w5919;
	wire w5920;
	wire w5921;
	wire w5922;
	wire w5923;
	wire w5924;
	wire w5925;
	wire w5926;
	wire w5927;
	wire w5928;
	wire w5929;
	wire w5930;
	wire w5931;
	wire w5932;
	wire w5933;
	wire w5934;
	wire w5935;
	wire w5936;
	wire w5937;
	wire w5938;
	wire w5939;
	wire w5940;
	wire w5941;
	wire w5942;
	wire w5943;
	wire w5944;
	wire w5945;
	wire w5946;
	wire w5947;
	wire w5948;
	wire w5949;
	wire w5950;
	wire w5951;
	wire w5952;
	wire w5953;
	wire w5954;
	wire w5955;
	wire w5956;
	wire w5957;
	wire w5958;
	wire w5959;
	wire w5960;
	wire w5961;
	wire w5962;
	wire w5963;
	wire w5964;
	wire w5965;
	wire w5966;
	wire w5967;
	wire w5968;
	wire w5969;
	wire w5970;
	wire w5971;
	wire w5972;
	wire w5973;
	wire w5974;
	wire w5975;
	wire w5976;
	wire w5977;
	wire w5978;
	wire w5979;
	wire w5980;
	wire w5981;
	wire w5982;
	wire w5983;
	wire w5984;
	wire w5985;
	wire w5986;
	wire w5987;
	wire w5988;
	wire w5989;
	wire w5990;
	wire w5991;
	wire w5992;
	wire w5993;
	wire w5994;
	wire w5995;
	wire w5996;
	wire w5997;
	wire w5998;
	wire w5999;
	wire w6000;
	wire w6001;
	wire w6002;
	wire w6003;
	wire w6004;
	wire w6005;
	wire w6006;
	wire w6007;
	wire w6008;
	wire w6009;
	wire w6010;
	wire w6011;
	wire w6012;
	wire w6013;
	wire w6014;
	wire w6015;
	wire w6016;
	wire w6017;
	wire w6018;
	wire w6019;
	wire w6020;
	wire w6021;
	wire w6022;
	wire w6023;
	wire w6024;
	wire w6025;
	wire w6026;
	wire w6027;
	wire w6028;
	wire w6029;
	wire w6030;
	wire w6031;
	wire w6032;
	wire w6033;
	wire w6034;
	wire w6035;
	wire w6036;
	wire w6037;
	wire w6038;
	wire w6039;
	wire w6040;
	wire w6041;
	wire w6042;
	wire w6043;
	wire w6044;
	wire w6045;
	wire w6046;
	wire w6047;
	wire w6048;
	wire w6049;
	wire w6050;
	wire w6051;
	wire w6052;
	wire w6053;
	wire w6054;
	wire w6055;
	wire w6056;
	wire w6057;
	wire w6058;
	wire w6059;
	wire w6060;
	wire w6061;
	wire w6062;
	wire w6063;
	wire w6064;
	wire w6065;
	wire w6066;
	wire w6067;
	wire w6068;
	wire w6069;
	wire w6070;
	wire w6071;
	wire w6072;
	wire w6073;
	wire w6074;
	wire w6075;
	wire w6076;
	wire w6077;
	wire w6078;
	wire w6079;
	wire w6080;
	wire w6081;
	wire w6082;
	wire w6083;
	wire w6084;
	wire w6085;
	wire w6086;
	wire w6087;
	wire w6088;
	wire w6089;
	wire w6090;
	wire w6091;
	wire w6092;
	wire w6093;
	wire w6094;
	wire w6095;
	wire w6096;
	wire w6097;
	wire w6098;
	wire w6099;
	wire w6100;
	wire w6101;
	wire w6102;
	wire w6103;
	wire w6104;
	wire w6105;
	wire w6106;
	wire w6107;
	wire w6108;
	wire w6109;
	wire w6110;
	wire w6111;
	wire w6112;
	wire w6113;
	wire w6114;
	wire w6115;
	wire w6116;
	wire w6117;
	wire w6118;
	wire w6119;
	wire w6120;
	wire w6121;
	wire w6122;
	wire w6123;
	wire w6124;
	wire w6125;
	wire w6126;
	wire w6127;
	wire w6128;
	wire w6129;
	wire w6130;
	wire w6131;
	wire w6132;
	wire w6133;
	wire w6134;
	wire w6135;
	wire w6136;
	wire w6137;
	wire w6138;
	wire w6139;
	wire w6140;
	wire w6141;
	wire w6142;
	wire w6143;
	wire w6144;
	wire w6145;
	wire w6146;
	wire w6147;
	wire w6148;
	wire w6149;
	wire w6150;
	wire w6151;
	wire w6152;
	wire w6153;
	wire w6154;
	wire w6155;
	wire w6156;
	wire w6157;
	wire w6158;
	wire w6159;
	wire w6160;
	wire w6161;
	wire w6162;
	wire w6163;
	wire w6164;
	wire w6165;
	wire w6166;
	wire w6167;
	wire w6168;
	wire w6169;
	wire w6170;
	wire w6171;
	wire w6172;
	wire w6173;
	wire w6174;
	wire w6175;
	wire w6176;
	wire w6177;
	wire w6178;
	wire w6179;
	wire w6180;
	wire w6181;
	wire w6182;
	wire w6183;
	wire w6184;
	wire w6185;
	wire w6186;
	wire w6187;
	wire w6188;
	wire w6189;
	wire w6190;
	wire w6191;
	wire w6192;
	wire w6193;
	wire w6194;
	wire w6195;
	wire w6196;
	wire w6197;
	wire w6198;
	wire w6199;
	wire w6200;
	wire w6201;
	wire w6202;
	wire w6203;
	wire w6204;
	wire w6205;
	wire w6206;
	wire w6207;
	wire w6208;
	wire w6209;
	wire w6210;
	wire w6211;
	wire w6212;
	wire w6213;
	wire w6214;
	wire w6215;
	wire w6216;
	wire w6217;
	wire w6218;
	wire w6219;
	wire w6220;
	wire w6221;
	wire w6222;
	wire w6223;
	wire w6224;
	wire w6225;
	wire w6226;
	wire w6227;
	wire w6228;
	wire w6229;
	wire w6230;
	wire w6231;
	wire w6232;
	wire w6233;
	wire w6234;
	wire w6235;
	wire w6236;
	wire w6237;
	wire w6238;
	wire w6239;
	wire w6240;
	wire w6241;
	wire w6242;
	wire w6243;
	wire w6244;
	wire w6245;
	wire w6246;
	wire w6247;
	wire w6248;
	wire w6249;
	wire w6250;
	wire w6251;
	wire w6252;
	wire w6253;
	wire w6254;
	wire w6255;
	wire w6256;
	wire w6257;
	wire w6258;
	wire w6259;
	wire w6260;
	wire w6261;
	wire w6262;
	wire w6263;
	wire w6264;
	wire w6265;
	wire w6266;
	wire w6267;
	wire w6268;
	wire w6269;
	wire w6270;
	wire w6271;
	wire w6272;
	wire w6273;
	wire w6274;
	wire w6275;
	wire w6276;
	wire w6277;
	wire w6278;
	wire w6279;
	wire w6280;
	wire w6281;
	wire w6282;
	wire w6283;
	wire w6284;
	wire w6285;
	wire w6286;
	wire w6287;
	wire w6288;
	wire w6289;
	wire w6290;
	wire w6291;
	wire w6292;
	wire w6293;
	wire w6294;
	wire w6295;
	wire w6296;
	wire w6297;
	wire w6298;
	wire w6299;
	wire w6300;
	wire w6301;
	wire w6302;
	wire w6303;
	wire w6304;
	wire w6305;
	wire w6306;
	wire w6307;
	wire w6308;
	wire w6309;
	wire w6310;
	wire w6311;
	wire w6312;
	wire w6313;
	wire w6314;
	wire w6315;
	wire w6316;
	wire w6317;
	wire w6318;
	wire w6319;
	wire w6320;
	wire w6321;
	wire w6322;
	wire w6323;
	wire w6324;
	wire w6325;
	wire w6326;
	wire w6327;
	wire w6328;
	wire w6329;
	wire w6330;
	wire w6331;
	wire w6332;
	wire w6333;
	wire w6334;
	wire w6335;
	wire w6336;
	wire w6337;
	wire w6338;
	wire w6339;
	wire w6340;
	wire w6341;
	wire w6342;
	wire w6343;
	wire w6344;
	wire w6345;
	wire w6346;
	wire w6347;
	wire w6348;
	wire w6349;
	wire w6350;
	wire w6351;
	wire w6352;
	wire w6353;
	wire w6354;
	wire w6355;
	wire w6356;
	wire w6357;
	wire w6358;
	wire w6359;
	wire w6360;
	wire w6361;
	wire w6362;
	wire w6363;
	wire w6364;
	wire w6365;
	wire w6366;
	wire w6367;
	wire w6368;
	wire w6369;
	wire w6370;
	wire w6371;
	wire w6372;
	wire w6373;
	wire w6374;
	wire w6375;
	wire w6376;
	wire w6377;
	wire w6378;
	wire w6379;
	wire w6380;
	wire w6381;
	wire w6382;
	wire w6383;
	wire w6384;
	wire w6385;
	wire w6386;
	wire w6387;
	wire w6388;
	wire w6389;
	wire w6390;
	wire w6391;
	wire w6392;
	wire w6393;
	wire w6394;
	wire w6395;
	wire w6396;
	wire w6397;
	wire w6398;
	wire w6399;
	wire w6400;
	wire w6401;
	wire w6402;
	wire w6403;
	wire w6404;
	wire w6405;
	wire w6406;
	wire w6407;
	wire w6408;
	wire w6409;
	wire w6410;
	wire w6411;
	wire w6412;
	wire w6413;
	wire w6414;
	wire w6415;
	wire w6416;
	wire w6417;
	wire w6418;
	wire w6419;
	wire w6420;
	wire w6421;
	wire w6422;
	wire w6423;
	wire w6424;
	wire w6425;
	wire w6426;
	wire w6427;
	wire w6428;
	wire w6429;
	wire w6430;
	wire w6431;
	wire w6432;
	wire w6433;
	wire w6434;
	wire w6435;
	wire w6436;
	wire w6437;
	wire w6438;
	wire w6439;
	wire w6440;
	wire w6441;
	wire w6442;
	wire w6443;
	wire w6444;
	wire w6445;
	wire w6446;
	wire w6447;
	wire w6448;
	wire w6449;
	wire w6450;
	wire w6451;
	wire w6452;
	wire w6453;
	wire w6454;
	wire w6455;
	wire w6456;
	wire w6457;
	wire w6458;
	wire w6459;
	wire w6460;
	wire w6461;
	wire w6462;
	wire w6463;
	wire w6464;
	wire w6465;
	wire w6466;
	wire w6467;
	wire w6468;
	wire w6469;
	wire w6470;
	wire w6471;
	wire w6472;
	wire w6473;
	wire w6474;
	wire w6475;
	wire w6476;
	wire w6477;
	wire w6478;
	wire w6479;
	wire w6480;
	wire w6481;
	wire w6482;
	wire w6483;
	wire w6484;
	wire w6485;
	wire w6486;
	wire w6487;
	wire w6488;
	wire w6489;
	wire w6490;
	wire w6491;
	wire w6492;
	wire w6493;
	wire w6494;
	wire w6495;
	wire w6496;
	wire w6497;
	wire w6498;
	wire w6499;
	wire w6500;
	wire w6501;
	wire w6502;
	wire w6503;
	wire w6504;
	wire w6505;
	wire w6506;
	wire w6507;
	wire w6508;
	wire w6509;
	wire w6510;
	wire w6511;
	wire w6512;
	wire w6513;
	wire w6514;
	wire w6515;
	wire w6516;
	wire w6517;
	wire w6518;
	wire w6519;
	wire w6520;
	wire w6521;
	wire w6522;
	wire w6523;
	wire w6524;
	wire w6525;
	wire w6526;
	wire w6527;
	wire w6528;
	wire w6529;
	wire w6530;
	wire w6531;
	wire w6532;
	wire w6533;
	wire w6534;
	wire w6535;
	wire w6536;
	wire w6537;
	wire w6538;
	wire w6539;
	wire w6540;
	wire w6541;
	wire w6542;
	wire w6543;
	wire w6544;
	wire w6545;
	wire w6546;
	wire w6547;
	wire w6548;
	wire w6549;
	wire w6550;
	wire w6551;
	wire w6552;
	wire w6553;
	wire w6554;
	wire w6555;
	wire w6556;
	wire w6557;
	wire w6558;
	wire w6559;
	wire w6560;
	wire w6561;
	wire w6562;
	wire w6563;
	wire w6564;
	wire w6565;
	wire w6566;
	wire w6567;
	wire w6568;
	wire w6569;
	wire w6570;
	wire w6571;
	wire w6572;
	wire w6573;
	wire w6574;
	wire w6575;
	wire w6576;
	wire w6577;
	wire w6578;
	wire w6579;
	wire w6580;
	wire w6581;
	wire w6582;
	wire w6583;
	wire w6584;
	wire w6585;
	wire w6586;
	wire w6587;
	wire w6588;
	wire w6589;
	wire w6590;
	wire w6591;
	wire w6592;
	wire w6593;
	wire w6594;
	wire w6595;
	wire w6596;
	wire w6597;
	wire w6598;
	wire w6599;
	wire w6600;
	wire w6601;
	wire w6602;
	wire w6603;
	wire w6604;
	wire w6605;
	wire w6606;
	wire w6607;
	wire w6608;
	wire w6609;
	wire w6610;
	wire w6611;
	wire w6612;
	wire w6613;
	wire w6614;
	wire w6615;
	wire w6616;
	wire w6617;
	wire w6618;
	wire w6619;
	wire w6620;
	wire w6621;
	wire w6622;
	wire w6623;
	wire w6624;
	wire w6625;
	wire w6626;
	wire w6627;
	wire w6628;
	wire w6629;
	wire w6630;
	wire w6631;
	wire w6632;
	wire w6633;
	wire w6634;
	wire w6635;
	wire w6636;
	wire w6637;
	wire w6638;
	wire w6639;
	wire w6640;
	wire w6641;
	wire w6642;
	wire w6643;
	wire w6644;
	wire w6645;
	wire w6646;
	wire w6647;
	wire w6648;
	wire w6649;
	wire w6650;
	wire w6651;
	wire w6652;
	wire w6653;
	wire w6654;
	wire w6655;
	wire w6656;
	wire w6657;
	wire w6658;
	wire w6659;
	wire w6660;
	wire w6661;
	wire w6662;
	wire w6663;
	wire w6664;
	wire w6665;
	wire w6666;
	wire w6667;
	wire w6668;
	wire w6669;
	wire w6670;
	wire w6671;
	wire w6672;
	wire w6673;
	wire w6674;
	wire w6675;
	wire w6676;
	wire w6677;
	wire w6678;
	wire w6679;
	wire w6680;
	wire w6681;
	wire w6682;
	wire w6683;
	wire w6684;
	wire w6685;
	wire w6686;
	wire w6687;
	wire w6688;
	wire w6689;
	wire w6690;
	wire w6691;
	wire w6692;
	wire w6693;
	wire w6694;
	wire w6695;
	wire w6696;
	wire w6697;
	wire w6698;
	wire w6699;
	wire w6700;
	wire w6701;
	wire w6702;
	wire w6703;
	wire w6704;
	wire w6705;
	wire w6706;
	wire w6707;
	wire w6708;
	wire w6709;
	wire w6710;
	wire w6711;
	wire w6712;
	wire w6713;
	wire w6714;
	wire w6715;
	wire w6716;
	wire w6717;
	wire w6718;
	wire w6719;
	wire w6720;
	wire w6721;
	wire w6722;
	wire w6723;
	wire w6724;
	wire w6725;
	wire w6726;
	wire w6727;
	wire w6728;
	wire w6729;
	wire w6730;
	wire w6731;
	wire w6732;
	wire w6733;
	wire w6734;
	wire w6735;
	wire w6736;
	wire w6737;
	wire w6738;
	wire w6739;
	wire w6740;
	wire w6741;
	wire w6742;
	wire w6743;
	wire w6744;
	wire w6745;
	wire w6746;
	wire w6747;
	wire w6748;
	wire w6749;
	wire w6750;
	wire w6751;
	wire w6752;
	wire w6753;
	wire w6754;
	wire w6755;
	wire w6756;
	wire w6757;
	wire w6758;
	wire w6759;
	wire w6760;
	wire w6761;
	wire w6762;
	wire w6763;
	wire w6764;
	wire w6765;
	wire w6766;
	wire w6767;
	wire w6768;
	wire w6769;
	wire w6770;
	wire w6771;
	wire w6772;
	wire w6773;
	wire w6774;
	wire w6775;
	wire w6776;
	wire w6777;
	wire w6778;
	wire w6779;
	wire w6780;
	wire w6781;
	wire w6782;
	wire w6783;
	wire w6784;
	wire w6785;
	wire w6786;
	wire w6787;
	wire w6788;
	wire w6789;
	wire w6790;
	wire w6791;
	wire w6792;
	wire w6793;
	wire w6794;
	wire w6795;
	wire w6796;
	wire w6797;
	wire w6798;
	wire w6799;
	wire w6800;
	wire w6801;
	wire w6802;
	wire w6803;
	wire w6804;
	wire w6805;
	wire w6806;
	wire w6807;
	wire w6808;
	wire w6809;
	wire w6810;
	wire w6811;
	wire w6812;
	wire w6813;
	wire w6814;
	wire w6815;
	wire w6816;
	wire w6817;
	wire w6818;
	wire w6819;
	wire w6820;
	wire w6821;
	wire w6822;
	wire w6823;
	wire w6824;
	wire w6825;

	assign CH0_EN = w2017;
	assign CH0VOL[0] = w2020;
	assign CH0VOL[1] = w2021;
	assign CH1_EN = w2016;
	assign CH1VOL[0] = w2080;
	assign CH1VOL[1] = w2081;
	assign CH2_EN = w2018;
	assign CH2VOL[0] = w2100;
	assign CH2VOL[1] = w2099;
	assign CH3_EN = w2015;
	assign CH3VOL[0] = w2122;
	assign CH3VOL[1] = w2121;
	assign PSGDAC0[0] = w2022;
	assign PSGDAC0[1] = w2023;
	assign PSGDAC0[2] = w2024;
	assign PSGDAC0[3] = w2025;
	assign PSGDAC0[4] = w2026;
	assign PSGDAC0[5] = w2027;
	assign PSGDAC0[6] = w2028;
	assign PSGDAC0[7] = w2029;
	assign PSGDAC1[0] = w2082;
	assign PSGDAC1[1] = w2083;
	assign PSGDAC1[2] = w2084;
	assign PSGDAC1[3] = w2085;
	assign PSGDAC1[4] = w2086;
	assign PSGDAC1[5] = w2087;
	assign PSGDAC1[6] = w2088;
	assign PSGDAC1[7] = w2089;
	assign PSGDAC2[0] = w2111;
	assign PSGDAC2[1] = w2112;
	assign PSGDAC2[2] = w2113;
	assign PSGDAC2[3] = w2114;
	assign PSGDAC2[4] = w2115;
	assign PSGDAC2[5] = w2116;
	assign PSGDAC2[6] = w2117;
	assign PSGDAC2[7] = w2118;
	assign PSGDAC3[0] = w2120;
	assign PSGDAC3[1] = w2119;
	assign PSGDAC3[2] = w2127;
	assign PSGDAC3[3] = w2126;
	assign PSGDAC3[4] = w2125;
	assign PSGDAC3[5] = w2124;
	assign PSGDAC3[6] = w2123;
	assign PSGDAC3[7] = w2128;
	assign w1207 = CAi[22];
	assign CAo[22] = w1366;
	assign CA[19] = CA[19];
	assign DTACK_OUT = w1056;
	assign Z80_INT = w1057;
	assign RA[7] = w1115;
	assign RA[6] = w1114;
	assign RA[5] = w1113;
	assign RA[4] = w1112;
	assign RA[2] = w1110;
	assign RA[1] = w1109;
	assign RA[0] = w1108;
	assign nRAS0 = w1342;
	assign RA[3] = w1111;
	assign nCAS0 = w1415;
	assign nOE0 = w1406;
	assign nLWR = w1407;
	assign nUWR = w1317;
	assign w1394 = DTACK_IN;
	assign w1002 = RnW;
	assign w1386 = nLDS;
	assign w1377 = nUDS;
	assign w1259 = nAS;
	assign w1375 = nM1;
	assign w1376 = nWR;
	assign w1373 = nRD;
	assign w1374 = nIORQ;
	assign nILP2 = w1379;
	assign nILP1 = w1378;
	assign w1240 = nINTAK;
	assign w1372 = nMREQ;
	assign w1242 = nBG;
	assign BGACK_OUT = w1257;
	assign w1393 = BGACK_IN;
	assign nBR = w1436;
	assign VSYNC = w1703;
	assign nCSYNC = w2004;
	assign w1697 = nCSYNC_IN;
	assign nHSYNC = w1762;
	assign w1974 = nHSYNC_IN;
	assign DB[15] = DB[15];
	assign DB[14] = DB[14];
	assign DB[13] = DB[13];
	assign DB[12] = DB[12];
	assign DB[11] = DB[11];
	assign DB[10] = DB[10];
	assign DB[9] = DB[9];
	assign DB[8] = DB[8];
	assign DB[7] = DB[7];
	assign DB[6] = DB[6];
	assign DB[5] = DB[5];
	assign DB[4] = DB[4];
	assign DB[3] = DB[3];
	assign DB[2] = DB[2];
	assign DB[1] = DB[1];
	assign DB[0] = DB[0];
	assign CA[0] = CA[0];
	assign CA[1] = CA[1];
	assign CA[2] = CA[2];
	assign CA[3] = CA[3];
	assign CA[4] = CA[4];
	assign CA[5] = CA[5];
	assign CA[6] = CA[6];
	assign CA[7] = CA[7];
	assign CA[8] = CA[8];
	assign CA[9] = CA[9];
	assign CA[10] = CA[10];
	assign CA[11] = CA[11];
	assign CA[12] = CA[12];
	assign CA[13] = CA[13];
	assign CA[14] = CA[14];
	assign CA[15] = CA[15];
	assign CA[17] = CA[17];
	assign CA[18] = CA[18];
	assign CA[20] = CA[20];
	assign CA[21] = CA[21];
	assign R_DAC[0] = w2953;
	assign R_DAC[1] = w2918;
	assign R_DAC[2] = w2952;
	assign R_DAC[3] = w2917;
	assign R_DAC[4] = w2951;
	assign R_DAC[5] = w2950;
	assign R_DAC[6] = w2949;
	assign R_DAC[7] = w2948;
	assign R_DAC[8] = w2914;
	assign G_DAC[0] = w2946;
	assign G_DAC[1] = w2945;
	assign G_DAC[2] = w2908;
	assign G_DAC[3] = w2907;
	assign G_DAC[4] = w2906;
	assign G_DAC[5] = w2905;
	assign G_DAC[6] = w2904;
	assign G_DAC[7] = w2903;
	assign G_DAC[8] = w2902;
	assign R_DAC[9] = w2915;
	assign R_DAC[10] = w2912;
	assign R_DAC[11] = w2916;
	assign R_DAC[12] = w2911;
	assign R_DAC[13] = w2913;
	assign R_DAC[14] = w2910;
	assign R_DAC[15] = w2909;
	assign R_DAC[16] = w2947;
	assign B_DAC[0] = w2894;
	assign B_DAC[1] = w2944;
	assign B_DAC[2] = w2940;
	assign B_DAC[3] = w2941;
	assign B_DAC[4] = w2942;
	assign B_DAC[5] = w2939;
	assign B_DAC[6] = w2943;
	assign B_DAC[7] = w3001;
	assign B_DAC[8] = w2895;
	assign G_DAC[9] = w2896;
	assign G_DAC[10] = w2901;
	assign G_DAC[11] = w2900;
	assign G_DAC[12] = w2999;
	assign G_DAC[13] = w2899;
	assign G_DAC[14] = w2898;
	assign G_DAC[15] = w2897;
	assign G_DAC[16] = w3000;
	assign B_DAC[9] = w2892;
	assign B_DAC[10] = w2893;
	assign B_DAC[11] = w2938;
	assign B_DAC[12] = w2937;
	assign B_DAC[13] = w2936;
	assign B_DAC[14] = w2935;
	assign B_DAC[15] = w2933;
	assign B_DAC[16] = w2934;
	assign nOE1 = nOE1;
	assign nWE0 = nWE0;
	assign nWE1 = nWE1;
	assign nCAS1 = nCAS1;
	assign nRAS1 = nRAS1;
	assign AD_RD_DIR = AD_RD_DIR;
	assign nYS = nYS;
	assign nSC = w2601;
	assign nSE0_1 = w2494;
	assign ADo[7] = w2454;
	assign ADo[6] = w2462;
	assign ADo[5] = w2639;
	assign ADo[4] = w2469;
	assign ADo[3] = w2579;
	assign ADo[2] = w2578;
	assign ADo[1] = w2530;
	assign ADo[0] = w2693;
	assign RDo[6] = w2640;
	assign RDo[5] = w2670;
	assign RDo[4] = w2645;
	assign RDo[3] = w2644;
	assign RDo[2] = w2672;
	assign RDo[1] = w2694;
	assign RDo[0] = w2501;
	assign w2541 = RDi[6];
	assign w2455 = RDi[7];
	assign w2468 = RDi[4];
	assign w2683 = RDi[5];
	assign w2535 = RDi[2];
	assign w2543 = RDi[3];
	assign w2673 = RDi[0];
	assign w2577 = RDi[1];
	assign w2542 = ADi[6];
	assign w2643 = ADi[7];
	assign w2487 = ADi[4];
	assign w2671 = ADi[5];
	assign w2529 = ADi[2];
	assign w2534 = ADi[3];
	assign w2502 = ADi[0];
	assign w2521 = ADi[1];
	assign RDo[7] = w2642;
	assign w5273 = SD[7];
	assign w5274 = SD[6];
	assign w6702 = SD[5];
	assign w6704 = SD[4];
	assign w5275 = SD[3];
	assign w5272 = SD[2];
	assign w6703 = SD[1];
	assign w5271 = SD[0];
	assign CLK1 = 68K CPU CLOCK;
	assign CLK0 = w1409;
	assign w4475 = EDCLKi;
	assign EDCLKo = EDCLK_O;
	assign w4451 = MCLK;
	assign SUB_CLK = w4440;
	assign w4493 = nRES_PAD;
	assign w1437 = 68kCLKi;
	assign EDCLKd = w1493;
	assign CA_PAD_DIR = w2451;
	assign DB_PAD_DIR = w2452;
	assign w406 = SEL0_M3;
	assign w6708 = nPAL;
	assign w440 = nHL;
	assign SPA/Bo = w2818;
	assign w2761 = SPA/Bi;

	// Instances

	vdp_slatch g1 (.nQ(w354), .D(VPOS[7]), .C(w1564), .nC(w1565) );
	vdp_slatch g2 (.nQ(w1527), .D(HPOS[8]), .C(w375), .nC(w376) );
	vdp_slatch g3 (.nQ(w359), .D(w301), .C(w1466), .nC(w377) );
	vdp_slatch g4 (.D(w302), .C(w1562), .nC(w1563), .nQ(w6810) );
	vdp_slatch g5 (.nQ(w360), .D(w361), .C(w1560), .nC(w1561) );
	vdp_slatch g6 (.nQ(w304), .D(w305), .C(w1558), .nC(w1559) );
	vdp_slatch g7 (.nQ(w362), .D(w361), .C(w378), .nC(w379) );
	vdp_slatch g8 (.nQ(w365), .D(w305), .C(w380), .nC(w381) );
	vdp_slatch g9 (.nQ(w363), .D(w361), .C(w429), .nC(w1463) );
	vdp_slatch g10 (.nQ(w366), .D(w305), .C(w1462), .nC(w386) );
	vdp_slatch g11 (.nQ(w364), .D(w361), .C(w384), .nC(w383) );
	vdp_slatch g12 (.nQ(w307), .D(w305), .C(w382), .nC(w1461) );
	vdp_slatch g13 (.Q(w305), .D(DB[7]), .C(w368), .nC(w367) );
	vdp_slatch g14 (.Q(w361), .D(w931), .C(w371), .nC(w370) );
	vdp_sr_bit g15 (.D(w308), .C2(HCLK2), .C1(HCLK1), .Q(FIFOo[7]), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g16 (.A(1'b1), .nZ(DB[7]), .nE(w1460) );
	vdp_notif0 g17 (.A(w307), .nZ(w308), .nE(w2019) );
	vdp_notif0 g18 (.A(w364), .nZ(w358), .nE(w385) );
	vdp_notif0 g19 (.A(w306), .nZ(AD_DATA[7]), .nE(w1605) );
	vdp_notif0 g20 (.A(w366), .nZ(w308), .nE(w1557) );
	vdp_notif0 g21 (.A(w363), .nZ(w358), .nE(w1604) );
	vdp_notif0 g22 (.A(w1533), .nZ(AD_DATA[7]), .nE(w403) );
	vdp_notif0 g23 (.A(w365), .nZ(w308), .nE(w402) );
	vdp_notif0 g24 (.A(w362), .nZ(w358), .nE(w1464) );
	vdp_notif0 g25 (.A(w1532), .nZ(AD_DATA[7]), .nE(w417) );
	vdp_notif0 g26 (.A(w304), .nZ(w308), .nE(w395) );
	vdp_notif0 g27 (.A(w303), .nZ(AD_DATA[7]), .nE(w415) );
	vdp_notif0 g28 (.A(w359), .nZ(DB[7]), .nE(w1602) );
	vdp_notif0 g29 (.nZ(DB[15]), .nE(w396), .A(w6810) );
	vdp_notif0 g30 (.A(w360), .nZ(w358), .nE(w1603) );
	vdp_notif0 g31 (.A(w354), .nZ(DB[15]), .nE(w1601) );
	vdp_notif0 g32 (.A(w432), .nZ(DB[7]), .nE(w397) );
	vdp_aon22 g33 (.Z(w432), .A1(w1527), .A2(w1566), .B1(w401), .B2(w354) );
	vdp_aon22 g34 (.A2(w399), .B1(w400), .B2(AD_DATA[7]), .A1(w358), .Z(w301) );
	vdp_aon22 g35 (.A2(w6716), .B1(w6717), .B2(w358), .A1(AD_DATA[7]), .Z(w302) );
	vdp_aon22 g36 (.Z(w303), .A2(w398), .B1(w1567), .B2(w304), .A1(w360) );
	vdp_aon22 g37 (.Z(w1532), .A2(w422), .B1(w421), .B2(w362), .A1(w365) );
	vdp_aon22 g38 (.Z(w1533), .A2(w430), .B1(w431), .B2(w363), .A1(w366) );
	vdp_aon22 g39 (.Z(w306), .A2(w6712), .B1(w6713), .B2(w307), .A1(w364) );
	vdp_aon22 g40 (.Z(w931), .A1(DB[15]), .A2(w369), .B1(w373), .B2(DB[7]) );
	vdp_slatch g41 (.nQ(w223), .D(VPOS[6]), .C(w1564), .nC(w1565) );
	vdp_slatch g42 (.nQ(w225), .D(HPOS[7]), .C(w375), .nC(w376) );
	vdp_slatch g43 (.nQ(w227), .D(w263), .C(w1466), .nC(w377) );
	vdp_slatch g44 (.nQ(w265), .D(w1433), .C(w1562), .nC(w1563) );
	vdp_slatch g45 (.nQ(w228), .D(w229), .C(w1560), .nC(w1561) );
	vdp_slatch g46 (.nQ(w267), .D(w268), .C(w1558), .nC(w1559) );
	vdp_slatch g47 (.nQ(w230), .D(w229), .C(w378), .nC(w379) );
	vdp_slatch g48 (.nQ(w232), .D(w268), .C(w380), .nC(w381) );
	vdp_slatch g49 (.nQ(w233), .D(w229), .C(w429), .nC(w1463) );
	vdp_slatch g50 (.nQ(w235), .D(w268), .C(w1462), .nC(w386) );
	vdp_slatch g51 (.nQ(w236), .D(w229), .C(w384), .nC(w383) );
	vdp_slatch g52 (.nQ(w270), .D(w268), .C(w382), .nC(w1461) );
	vdp_slatch g53 (.Q(w268), .D(DB[6]), .C(w368), .nC(w367) );
	vdp_slatch g54 (.Q(w229), .D(w271), .C(w371), .nC(w370) );
	vdp_sr_bit g55 (.D(w264), .Q(FIFOo[6]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g56 (.A(1'b1), .nZ(DB[6]), .nE(w1460) );
	vdp_notif0 g57 (.A(w270), .nZ(w264), .nE(w2019) );
	vdp_notif0 g58 (.A(w236), .nZ(RD_DATA[6]), .nE(w385) );
	vdp_notif0 g59 (.A(w269), .nZ(AD_DATA[6]), .nE(w1605) );
	vdp_notif0 g60 (.A(w235), .nZ(w264), .nE(w1557) );
	vdp_notif0 g61 (.A(w233), .nZ(RD_DATA[6]), .nE(w1604) );
	vdp_notif0 g62 (.A(w234), .nZ(AD_DATA[6]), .nE(w403) );
	vdp_notif0 g63 (.A(w232), .nZ(w264), .nE(w402) );
	vdp_notif0 g64 (.A(w230), .nZ(RD_DATA[6]), .nE(w1464) );
	vdp_notif0 g65 (.A(w231), .nZ(AD_DATA[6]), .nE(w417) );
	vdp_notif0 g66 (.A(w267), .nZ(w264), .nE(w395) );
	vdp_notif0 g67 (.A(w266), .nZ(AD_DATA[6]), .nE(w415) );
	vdp_notif0 g68 (.A(w227), .nZ(DB[6]), .nE(w1602) );
	vdp_notif0 g69 (.A(w265), .nZ(DB[14]), .nE(w396) );
	vdp_notif0 g70 (.A(w228), .nZ(RD_DATA[6]), .nE(w1603) );
	vdp_notif0 g71 (.A(w223), .nZ(DB[14]), .nE(w1601) );
	vdp_notif0 g72 (.A(w226), .nZ(DB[6]), .nE(w397) );
	vdp_aon22 g73 (.A2(w1566), .B1(w401), .B2(w223), .A1(w225), .Z(w226) );
	vdp_aon22 g74 (.Z(w263), .A2(w399), .B1(w400), .B2(AD_DATA[6]), .A1(RD_DATA[6]) );
	vdp_aon22 g75 (.Z(w1433), .A2(w6716), .B1(w6717), .B2(RD_DATA[6]), .A1(AD_DATA[6]) );
	vdp_aon22 g76 (.Z(w266), .A2(w398), .B1(w1567), .B2(w267), .A1(w228) );
	vdp_aon22 g77 (.Z(w231), .A2(w422), .B1(w421), .B2(w232), .A1(w230) );
	vdp_aon22 g78 (.Z(w234), .A2(w430), .B1(w431), .B2(w235), .A1(w233) );
	vdp_aon22 g79 (.Z(w269), .A2(w6712), .B1(w6713), .B2(w270), .A1(w236) );
	vdp_aon22 g80 (.Z(w271), .A1(DB[14]), .A2(w369), .B1(w373), .B2(DB[6]) );
	vdp_slatch g81 (.nQ(w338), .D(VPOS[5]), .C(w1564), .nC(w1565) );
	vdp_slatch g82 (.nQ(w1528), .D(HPOS[6]), .C(w375), .nC(w376) );
	vdp_slatch g83 (.nQ(w343), .D(w292), .C(w1466), .nC(w377) );
	vdp_slatch g84 (.D(w293), .C(w1562), .nC(w1563), .nQ(w6811) );
	vdp_slatch g85 (.nQ(w344), .D(w350), .C(w1560), .nC(w1561) );
	vdp_slatch g86 (.nQ(w295), .D(w296), .C(w1558), .nC(w1559) );
	vdp_slatch g87 (.nQ(w346), .D(w350), .C(w378), .nC(w379) );
	vdp_slatch g88 (.nQ(w345), .D(w296), .C(w380), .nC(w381) );
	vdp_slatch g89 (.nQ(w348), .D(w350), .C(w429), .nC(w1463) );
	vdp_slatch g90 (.nQ(w351), .D(w296), .C(w1462), .nC(w386) );
	vdp_slatch g91 (.nQ(w352), .D(w350), .C(w384), .nC(w383) );
	vdp_slatch g92 (.nQ(w298), .D(w296), .C(w382), .nC(w1461) );
	vdp_slatch g93 (.Q(w296), .D(DB[5]), .C(w368), .nC(w367) );
	vdp_slatch g94 (.Q(w350), .D(w299), .C(w371), .nC(w370) );
	vdp_sr_bit g95 (.D(w300), .Q(FIFOo[5]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g96 (.A(1'b1), .nZ(DB[5]), .nE(w1460) );
	vdp_notif0 g97 (.A(w298), .nZ(w300), .nE(w2019) );
	vdp_notif0 g98 (.A(w352), .nZ(RD_DATA[5]), .nE(w385) );
	vdp_notif0 g99 (.A(w297), .nZ(w291), .nE(w1605) );
	vdp_notif0 g100 (.A(w351), .nZ(w300), .nE(w1557) );
	vdp_notif0 g101 (.A(w348), .nZ(RD_DATA[5]), .nE(w1604) );
	vdp_notif0 g102 (.A(w349), .nZ(w291), .nE(w403) );
	vdp_notif0 g103 (.A(w345), .nZ(w300), .nE(w402) );
	vdp_notif0 g104 (.A(w346), .nZ(RD_DATA[5]), .nE(w1464) );
	vdp_notif0 g105 (.A(w347), .nZ(w291), .nE(w417) );
	vdp_notif0 g106 (.A(w295), .nZ(w300), .nE(w395) );
	vdp_notif0 g107 (.A(w294), .nZ(w291), .nE(w415) );
	vdp_notif0 g108 (.A(w343), .nZ(DB[5]), .nE(w1602) );
	vdp_notif0 g109 (.nZ(DB[13]), .nE(w396), .A(w6811) );
	vdp_notif0 g110 (.A(w344), .nZ(RD_DATA[5]), .nE(w1603) );
	vdp_notif0 g111 (.A(w338), .nZ(DB[13]), .nE(w1601) );
	vdp_notif0 g112 (.A(w342), .nZ(DB[5]), .nE(w397) );
	vdp_aon22 g113 (.Z(w342), .A1(w1528), .A2(w1566), .B1(w401), .B2(w338) );
	vdp_aon22 g114 (.A2(w399), .B1(w400), .B2(w291), .A1(RD_DATA[5]), .Z(w292) );
	vdp_aon22 g115 (.A2(w6716), .B1(w6717), .B2(RD_DATA[5]), .A1(w291), .Z(w293) );
	vdp_aon22 g116 (.Z(w294), .A2(w398), .B1(w1567), .B2(w295), .A1(w344) );
	vdp_aon22 g117 (.Z(w347), .A2(w422), .B1(w421), .B2(w346), .A1(w345) );
	vdp_aon22 g118 (.Z(w349), .A2(w430), .B1(w431), .B2(w348), .A1(w351) );
	vdp_aon22 g119 (.Z(w297), .A2(w6712), .B1(w6713), .B2(w298), .A1(w352) );
	vdp_aon22 g120 (.Z(w299), .A1(DB[13]), .A2(w369), .B1(w373), .B2(DB[5]) );
	vdp_slatch g121 (.nQ(w208), .D(VPOS[4]), .C(w1564), .nC(w1565) );
	vdp_slatch g122 (.nQ(w210), .D(HPOS[5]), .C(w375), .nC(w376) );
	vdp_slatch g123 (.nQ(w1568), .D(w255), .C(w1466), .nC(w377) );
	vdp_slatch g124 (.D(w1531), .C(w1562), .nC(w1563), .nQ(w6812) );
	vdp_slatch g125 (.nQ(w212), .D(w213), .C(w1560), .nC(w1561) );
	vdp_slatch g126 (.nQ(w258), .D(w259), .C(w1558), .nC(w1559) );
	vdp_slatch g127 (.nQ(w214), .D(w213), .C(w378), .nC(w379) );
	vdp_slatch g128 (.nQ(w216), .D(w259), .C(w380), .nC(w381) );
	vdp_slatch g129 (.nQ(w217), .D(w213), .C(w429), .nC(w1463) );
	vdp_slatch g130 (.nQ(w219), .D(w259), .C(w1462), .nC(w386) );
	vdp_slatch g131 (.nQ(w220), .D(w213), .C(w384), .nC(w383) );
	vdp_slatch g132 (.nQ(w261), .D(w259), .C(w382), .nC(w1461) );
	vdp_slatch g133 (.Q(w259), .D(DB[4]), .C(w368), .nC(w367) );
	vdp_slatch g134 (.Q(w213), .D(w262), .C(w371), .nC(w370) );
	vdp_sr_bit g135 (.D(w256), .Q(FIFOo[4]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g136 (.A(1'b1), .nZ(DB[4]), .nE(w1460) );
	vdp_notif0 g137 (.A(w261), .nZ(w256), .nE(w2019) );
	vdp_notif0 g138 (.A(w220), .nZ(RD_DATA[4]), .nE(w385) );
	vdp_notif0 g139 (.A(w260), .nZ(AD_DATA[4]), .nE(w1605) );
	vdp_notif0 g140 (.A(w219), .nZ(w256), .nE(w1557) );
	vdp_notif0 g141 (.A(w217), .nZ(RD_DATA[4]), .nE(w1604) );
	vdp_notif0 g142 (.A(w218), .nZ(AD_DATA[4]), .nE(w403) );
	vdp_notif0 g143 (.A(w216), .nZ(w256), .nE(w402) );
	vdp_notif0 g144 (.A(w214), .nZ(RD_DATA[4]), .nE(w1464) );
	vdp_notif0 g145 (.A(w215), .nZ(AD_DATA[4]), .nE(w417) );
	vdp_notif0 g146 (.A(w258), .nZ(w256), .nE(w395) );
	vdp_notif0 g147 (.A(w257), .nZ(AD_DATA[4]), .nE(w415) );
	vdp_notif0 g148 (.A(w1568), .nZ(DB[4]), .nE(w1602) );
	vdp_notif0 g149 (.nZ(DB[12]), .nE(w396), .A(w6812) );
	vdp_notif0 g150 (.A(w212), .nZ(RD_DATA[4]), .nE(w1603) );
	vdp_notif0 g151 (.A(w208), .nZ(DB[12]), .nE(w1601) );
	vdp_notif0 g152 (.A(w211), .nZ(DB[4]), .nE(w397) );
	vdp_aon22 g153 (.A2(w1566), .B1(w401), .B2(w208), .A1(w210), .Z(w211) );
	vdp_aon22 g154 (.Z(w255), .A2(w399), .B1(w400), .B2(AD_DATA[4]), .A1(RD_DATA[4]) );
	vdp_aon22 g155 (.Z(w1531), .A2(w6716), .B1(w6717), .B2(RD_DATA[4]), .A1(AD_DATA[4]) );
	vdp_aon22 g156 (.Z(w257), .A2(w398), .B1(w1567), .B2(w258), .A1(w212) );
	vdp_aon22 g157 (.Z(w215), .A2(w422), .B1(w421), .B2(w216), .A1(w214) );
	vdp_aon22 g158 (.Z(w218), .A2(w430), .B1(w431), .B2(w219), .A1(w217) );
	vdp_aon22 g159 (.Z(w260), .A2(w6712), .B1(w6713), .B2(w261), .A1(w220) );
	vdp_aon22 g160 (.Z(w262), .A1(DB[12]), .A2(w369), .B1(w373), .B2(DB[4]) );
	vdp_slatch g161 (.nQ(w322), .D(VPOS[3]), .C(w1564), .nC(w1565) );
	vdp_slatch g162 (.nQ(w1529), .D(HPOS[4]), .C(w375), .nC(w376) );
	vdp_slatch g163 (.nQ(w327), .D(w282), .C(w1466), .nC(w377) );
	vdp_slatch g164 (.D(w283), .C(w1562), .nC(w1563), .nQ(w6813) );
	vdp_slatch g165 (.nQ(w328), .D(w331), .C(w1560), .nC(w1561) );
	vdp_slatch g166 (.nQ(w285), .D(w286), .C(w1558), .nC(w1559) );
	vdp_slatch g167 (.nQ(w329), .D(w331), .C(w378), .nC(w379) );
	vdp_slatch g168 (.nQ(w330), .D(w286), .C(w380), .nC(w381) );
	vdp_slatch g169 (.nQ(w333), .D(w331), .C(w429), .nC(w1463) );
	vdp_slatch g170 (.nQ(w335), .D(w286), .C(w1462), .nC(w386) );
	vdp_slatch g171 (.nQ(w336), .D(w331), .C(w384), .nC(w383) );
	vdp_slatch g172 (.nQ(w288), .D(w286), .C(w382), .nC(w1461) );
	vdp_slatch g173 (.Q(w286), .D(DB[3]), .C(w368), .nC(w367) );
	vdp_slatch g174 (.Q(w331), .D(w289), .C(w371), .nC(w370) );
	vdp_sr_bit g175 (.D(w290), .Q(FIFOo[3]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g176 (.A(1'b1), .nZ(DB[3]), .nE(w1460) );
	vdp_notif0 g177 (.A(w288), .nZ(w290), .nE(w2019) );
	vdp_notif0 g178 (.A(w336), .nZ(w324), .nE(w385) );
	vdp_notif0 g179 (.A(w287), .nZ(AD_DATA[3]), .nE(w1605) );
	vdp_notif0 g180 (.A(w335), .nZ(w290), .nE(w1557) );
	vdp_notif0 g181 (.A(w333), .nZ(w324), .nE(w1604) );
	vdp_notif0 g182 (.A(w334), .nZ(AD_DATA[3]), .nE(w403) );
	vdp_notif0 g183 (.A(w330), .nZ(w290), .nE(w402) );
	vdp_notif0 g184 (.A(w329), .nZ(w324), .nE(w1464) );
	vdp_notif0 g185 (.A(w332), .nZ(AD_DATA[3]), .nE(w417) );
	vdp_notif0 g186 (.A(w285), .nZ(w290), .nE(w395) );
	vdp_notif0 g187 (.A(w284), .nZ(AD_DATA[3]), .nE(w415) );
	vdp_notif0 g188 (.A(w327), .nZ(DB[3]), .nE(w1602) );
	vdp_notif0 g189 (.nZ(DB[11]), .nE(w396), .A(w6813) );
	vdp_notif0 g190 (.A(w328), .nZ(w324), .nE(w1603) );
	vdp_notif0 g191 (.A(w322), .nZ(DB[11]), .nE(w1601) );
	vdp_notif0 g192 (.A(w326), .nZ(DB[3]), .nE(w397) );
	vdp_aon22 g193 (.Z(w326), .A1(w1529), .A2(w1566), .B1(w401), .B2(w322) );
	vdp_aon22 g194 (.A2(w399), .B1(w400), .B2(AD_DATA[3]), .A1(w324), .Z(w282) );
	vdp_aon22 g195 (.A2(w6716), .B1(w6717), .B2(w324), .A1(AD_DATA[3]), .Z(w283) );
	vdp_aon22 g196 (.Z(w284), .A2(w398), .B1(w1567), .B2(w285), .A1(w328) );
	vdp_aon22 g197 (.Z(w332), .A2(w422), .B1(w421), .B2(w329), .A1(w330) );
	vdp_aon22 g198 (.Z(w334), .A2(w430), .B1(w431), .B2(w333), .A1(w335) );
	vdp_aon22 g199 (.Z(w287), .A2(w6712), .B1(w6713), .B2(w288), .A1(w336) );
	vdp_aon22 g200 (.Z(w289), .A1(DB[11]), .A2(w369), .B1(w373), .B2(DB[3]) );
	vdp_slatch g201 (.nQ(w193), .D(VPOS[2]), .C(w1564), .nC(w1565) );
	vdp_slatch g202 (.nQ(w1569), .D(HPOS[3]), .C(w375), .nC(w376) );
	vdp_slatch g203 (.nQ(w195), .D(w246), .C(w1466), .nC(w377) );
	vdp_slatch g204 (.D(w1467), .C(w1562), .nC(w1563), .nQ(w6814) );
	vdp_slatch g205 (.nQ(w196), .D(w199), .C(w1560), .nC(w1561) );
	vdp_slatch g206 (.nQ(w249), .D(w250), .C(w1558), .nC(w1559) );
	vdp_slatch g207 (.nQ(w197), .D(w199), .C(w378), .nC(w379) );
	vdp_slatch g208 (.nQ(w200), .D(w250), .C(w380), .nC(w381) );
	vdp_slatch g209 (.nQ(w201), .D(w199), .C(w429), .nC(w1463) );
	vdp_slatch g210 (.nQ(w203), .D(w250), .C(w1462), .nC(w386) );
	vdp_slatch g211 (.nQ(w204), .D(w199), .C(w384), .nC(w383) );
	vdp_slatch g212 (.nQ(w252), .D(w250), .C(w382), .nC(w1461) );
	vdp_slatch g213 (.Q(w250), .D(DB[2]), .C(w368), .nC(w367) );
	vdp_slatch g214 (.Q(w199), .D(w253), .C(w371), .nC(w370) );
	vdp_sr_bit g215 (.D(w247), .Q(FIFOo[2]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g216 (.A(w205), .nZ(DB[2]), .nE(w1460) );
	vdp_notif0 g217 (.A(w252), .nZ(w247), .nE(w2019) );
	vdp_notif0 g218 (.A(w204), .nZ(RD_DATA[2]), .nE(w385) );
	vdp_notif0 g219 (.A(w251), .nZ(AD_DATA[2]), .nE(w1605) );
	vdp_notif0 g220 (.A(w203), .nZ(w247), .nE(w1557) );
	vdp_notif0 g221 (.A(w201), .nZ(RD_DATA[2]), .nE(w1604) );
	vdp_notif0 g222 (.A(w202), .nZ(AD_DATA[2]), .nE(w403) );
	vdp_notif0 g223 (.A(w200), .nZ(w247), .nE(w402) );
	vdp_notif0 g224 (.A(w197), .nZ(RD_DATA[2]), .nE(w1464) );
	vdp_notif0 g225 (.A(w198), .nZ(AD_DATA[2]), .nE(w417) );
	vdp_notif0 g226 (.A(w249), .nZ(w247), .nE(w395) );
	vdp_notif0 g227 (.A(w248), .nZ(AD_DATA[2]), .nE(w415) );
	vdp_notif0 g228 (.A(w195), .nZ(DB[2]), .nE(w1602) );
	vdp_notif0 g229 (.nZ(DB[10]), .nE(w396), .A(w6814) );
	vdp_notif0 g230 (.A(w196), .nZ(RD_DATA[2]), .nE(w1603) );
	vdp_notif0 g231 (.A(w193), .nZ(DB[10]), .nE(w1601) );
	vdp_notif0 g232 (.A(w194), .nZ(DB[2]), .nE(w397) );
	vdp_aon22 g233 (.A2(w1566), .B1(w401), .B2(w193), .A1(w1569), .Z(w194) );
	vdp_aon22 g234 (.Z(w246), .A2(w399), .B1(w400), .B2(AD_DATA[2]), .A1(RD_DATA[2]) );
	vdp_aon22 g235 (.Z(w1467), .A2(w6716), .B1(w6717), .B2(RD_DATA[2]), .A1(AD_DATA[2]) );
	vdp_aon22 g236 (.Z(w248), .A2(w398), .B1(w1567), .B2(w249), .A1(w196) );
	vdp_aon22 g237 (.Z(w198), .A2(w422), .B1(w421), .B2(w200), .A1(w197) );
	vdp_aon22 g238 (.Z(w202), .A2(w430), .B1(w431), .B2(w203), .A1(w201) );
	vdp_aon22 g239 (.Z(w251), .A2(w6712), .B1(w6713), .B2(w252), .A1(w204) );
	vdp_aon22 g240 (.Z(w253), .A1(DB[10]), .A2(w369), .B1(w373), .B2(DB[2]) );
	vdp_slatch g241 (.nQ(w309), .D(VPOS[1]), .C(w1564), .nC(w1565) );
	vdp_slatch g242 (.nQ(w1530), .D(HPOS[2]), .C(w375), .nC(w376) );
	vdp_slatch g243 (.nQ(w312), .D(w272), .C(w1466), .nC(w377) );
	vdp_slatch g244 (.D(w273), .C(w1562), .nC(w1563), .nQ(w6815) );
	vdp_slatch g245 (.nQ(w313), .D(w316), .C(w1560), .nC(w1561) );
	vdp_slatch g246 (.nQ(w275), .D(w276), .C(w1558), .nC(w1559) );
	vdp_slatch g247 (.nQ(w315), .D(w316), .C(w378), .nC(w379) );
	vdp_slatch g248 (.nQ(w314), .D(w276), .C(w380), .nC(w381) );
	vdp_slatch g249 (.nQ(w318), .D(w316), .C(w429), .nC(w1463) );
	vdp_slatch g250 (.nQ(w320), .D(w276), .C(w1462), .nC(w386) );
	vdp_slatch g251 (.nQ(w321), .D(w316), .C(w384), .nC(w383) );
	vdp_slatch g252 (.nQ(w278), .D(w276), .C(w382), .nC(w1461) );
	vdp_slatch g253 (.Q(w276), .D(DB[1]), .C(w368), .nC(w367) );
	vdp_slatch g254 (.Q(w316), .D(w280), .C(w371), .nC(w370) );
	vdp_sr_bit g255 (.D(w281), .Q(FIFOo[1]), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g256 (.A(w1606), .nZ(DB[1]), .nE(w1460) );
	vdp_notif0 g257 (.A(w278), .nZ(w281), .nE(w2019) );
	vdp_notif0 g258 (.A(w321), .nZ(RD_DATA[1]), .nE(w385) );
	vdp_notif0 g259 (.A(w277), .nZ(AD_DATA[1]), .nE(w1605) );
	vdp_notif0 g260 (.A(w320), .nZ(w281), .nE(w1557) );
	vdp_notif0 g261 (.A(w318), .nZ(RD_DATA[1]), .nE(w1604) );
	vdp_notif0 g262 (.A(w319), .nZ(AD_DATA[1]), .nE(w403) );
	vdp_notif0 g263 (.A(w314), .nZ(w281), .nE(w402) );
	vdp_notif0 g264 (.A(w315), .nZ(RD_DATA[1]), .nE(w1464) );
	vdp_notif0 g265 (.A(w317), .nZ(AD_DATA[1]), .nE(w417) );
	vdp_notif0 g266 (.A(w275), .nZ(w281), .nE(w395) );
	vdp_notif0 g267 (.A(w274), .nZ(AD_DATA[1]), .nE(w415) );
	vdp_notif0 g268 (.A(w312), .nZ(DB[1]), .nE(w1602) );
	vdp_notif0 g269 (.nZ(DB[9]), .nE(w396), .A(w6815) );
	vdp_notif0 g270 (.A(w313), .nZ(RD_DATA[1]), .nE(w1603) );
	vdp_notif0 g271 (.A(w309), .nZ(DB[9]), .nE(w1601) );
	vdp_notif0 g272 (.A(w1465), .nZ(DB[1]), .nE(w397) );
	vdp_aon22 g273 (.Z(w1465), .A1(w1530), .A2(w1566), .B1(w401), .B2(w309) );
	vdp_aon22 g274 (.A2(w399), .B1(w400), .B2(AD_DATA[1]), .A1(RD_DATA[1]), .Z(w272) );
	vdp_aon22 g275 (.A2(w6716), .B1(w6717), .B2(RD_DATA[1]), .A1(AD_DATA[1]), .Z(w273) );
	vdp_aon22 g276 (.Z(w274), .A2(w398), .B1(w1567), .B2(w275), .A1(w313) );
	vdp_aon22 g277 (.Z(w317), .A2(w422), .B1(w421), .B2(w315), .A1(w314) );
	vdp_aon22 g278 (.Z(w319), .A2(w430), .B1(w431), .B2(w318), .A1(w320) );
	vdp_aon22 g279 (.Z(w277), .A2(w6712), .B1(w6713), .B2(w278), .A1(w321) );
	vdp_aon22 g280 (.Z(w280), .A1(DB[9]), .A2(w369), .B1(w373), .B2(DB[1]) );
	vdp_slatch g281 (.nQ(w178), .D(w176), .C(w1564), .nC(w1565) );
	vdp_slatch g282 (.D(HPOS[1]), .nQ(w1459), .C(w375), .nC(w376) );
	vdp_slatch g283 (.nQ(w180), .D(w238), .C(w1466), .nC(w377) );
	vdp_slatch g284 (.D(w1434), .C(w1562), .nC(w1563), .nQ(w6816) );
	vdp_slatch g285 (.nQ(w181), .D(w185), .C(w1560), .nC(w1561) );
	vdp_slatch g286 (.nQ(w241), .D(w242), .C(w1558), .nC(w1559) );
	vdp_slatch g287 (.nQ(w182), .D(w185), .C(w378), .nC(w379) );
	vdp_slatch g288 (.nQ(w184), .D(w242), .C(w380), .nC(w381) );
	vdp_slatch g289 (.nQ(w186), .D(w185), .C(w429), .nC(w1463) );
	vdp_slatch g290 (.nQ(w188), .D(w242), .C(w1462), .nC(w386) );
	vdp_slatch g291 (.nQ(w189), .D(w185), .C(w384), .nC(w383) );
	vdp_slatch g292 (.nQ(w244), .D(w242), .C(w382), .nC(w1461) );
	vdp_slatch g293 (.Q(w242), .D(DB[0]), .C(w368), .nC(w367) );
	vdp_slatch g294 (.D(w245), .Q(w185), .C(w371), .nC(w370) );
	vdp_sr_bit g295 (.D(w239), .C2(HCLK2), .C1(HCLK1), .Q(FIFOo[0]), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_notif0 g296 (.A(1'b1), .nZ(DB[0]), .nE(w1460) );
	vdp_notif0 g297 (.A(w244), .nZ(w239), .nE(w2019) );
	vdp_notif0 g298 (.A(w189), .nZ(RD_DATA[0]), .nE(w385) );
	vdp_notif0 g299 (.A(w243), .nZ(AD_DATA[0]), .nE(w1605) );
	vdp_notif0 g300 (.A(w188), .nZ(w239), .nE(w1557) );
	vdp_notif0 g301 (.A(w186), .nZ(RD_DATA[0]), .nE(w1604) );
	vdp_notif0 g302 (.A(w187), .nZ(AD_DATA[0]), .nE(w403) );
	vdp_notif0 g303 (.A(w184), .nZ(w239), .nE(w402) );
	vdp_notif0 g304 (.A(w182), .nZ(RD_DATA[0]), .nE(w1464) );
	vdp_notif0 g305 (.A(w183), .nZ(AD_DATA[0]), .nE(w417) );
	vdp_notif0 g306 (.A(w241), .nZ(w239), .nE(w395) );
	vdp_notif0 g307 (.A(w240), .nZ(AD_DATA[0]), .nE(w415) );
	vdp_notif0 g308 (.A(w180), .nZ(DB[0]), .nE(w1602) );
	vdp_notif0 g309 (.nZ(DB[8]), .nE(w396), .A(w6816) );
	vdp_notif0 g310 (.A(w181), .nZ(RD_DATA[0]), .nE(w1603) );
	vdp_notif0 g311 (.A(w178), .nZ(DB[8]), .nE(w1601) );
	vdp_notif0 g312 (.A(w179), .nZ(DB[0]), .nE(w397) );
	vdp_aon22 g313 (.A2(w1566), .B1(w401), .B2(w178), .A1(w1459), .Z(w179) );
	vdp_aon22 g314 (.Z(w238), .A2(w399), .B1(w400), .B2(AD_DATA[0]), .A1(RD_DATA[0]) );
	vdp_aon22 g315 (.Z(w1434), .A2(w6716), .B1(w6717), .B2(RD_DATA[0]), .A1(AD_DATA[0]) );
	vdp_aon22 g316 (.Z(w240), .A2(w398), .B1(w1567), .B2(w241), .A1(w181) );
	vdp_aon22 g317 (.Z(w183), .A2(w422), .B1(w421), .B2(w184), .A1(w182) );
	vdp_aon22 g318 (.Z(w187), .A2(w430), .B1(w431), .B2(w188), .A1(w186) );
	vdp_aon22 g319 (.Z(w243), .A2(w6712), .B1(w6713), .B2(w244), .A1(w189) );
	vdp_aon22 g320 (.Z(w245), .A1(DB[8]), .A2(w369), .B1(w373), .B2(DB[0]) );
	vdp_not g321 (.A(w279), .nZ(w1606) );
	vdp_not g322 (.A(w254), .nZ(w205) );
	vdp_not g323 (.A(w405), .nZ(w1601) );
	vdp_not g324 (.A(w409), .nZ(w397) );
	vdp_not g325 (.A(w414), .nZ(w1602) );
	vdp_not g326 (.A(w414), .nZ(w396) );
	vdp_sr_bit g327 (.D(w413), .C2(HCLK2), .C1(HCLK1), .Q(w947), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g328 (.D(w459), .Q(w428), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g329 (.D(w428), .Q(w425), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g330 (.D(w425), .Q(w419), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g331 (.D(w423), .Q(w465), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g332 (.D(w465), .Q(w420), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g333 (.D(w466), .Q(w413), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g334 (.D(w416), .Q(w410), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g335 (.A(w448), .nZ(w1603) );
	vdp_not g336 (.A(w448), .nZ(w415) );
	vdp_not g337 (.A(w448), .nZ(w395) );
	vdp_not g338 (.A(w450), .nZ(w1464) );
	vdp_not g339 (.A(w450), .nZ(w417) );
	vdp_not g340 (.A(w450), .nZ(w402) );
	vdp_not g341 (.A(w462), .nZ(w1604) );
	vdp_not g342 (.A(w462), .nZ(w403) );
	vdp_not g343 (.A(w462), .nZ(w1557) );
	vdp_not g344 (.A(w451), .nZ(w385) );
	vdp_not g345 (.A(w451), .nZ(w1605) );
	vdp_not g346 (.A(w451), .nZ(w2019) );
	vdp_not g347 (.A(w427), .nZ(w1460) );
	vdp_not g348 (.A(w425), .nZ(w404) );
	vdp_not g349 (.A(w406), .nZ(w407) );
	vdp_comp_str g350 (.A(w441), .Z(w1564), .nZ(w1565) );
	vdp_comp_str g351 (.A(w442), .Z(w375), .nZ(w376) );
	vdp_comp_str g352 (.A(w411), .Z(w1466), .nZ(w377) );
	vdp_comp_str g353 (.A(w412), .Z(w1562), .nZ(w1563) );
	vdp_comp_str g354 (.A(w467), .Z(w1560), .nZ(w1561) );
	vdp_comp_str g355 (.A(w467), .Z(w1558), .nZ(w1559) );
	vdp_comp_str g356 (.A(w464), .Z(w378), .nZ(w379) );
	vdp_comp_str g357 (.A(w464), .Z(w380), .nZ(w381) );
	vdp_comp_str g358 (.A(w508), .Z(w429), .nZ(w1463) );
	vdp_comp_str g359 (.A(w508), .Z(w1462), .nZ(w386) );
	vdp_comp_str g360 (.A(w458), .Z(w384), .nZ(w383) );
	vdp_comp_str g361 (.A(w458), .Z(w382), .nZ(w1461) );
	vdp_comp_str g362 (.A(w469), .Z(w368), .nZ(w367) );
	vdp_comp_str g363 (.A(w469), .Z(w371), .nZ(w370) );
	vdp_comp_we g364 (.A(w406), .Z(w369), .nZ(w373) );
	vdp_comp_we g365 (.A(w447), .Z(w6712), .nZ(w6713) );
	vdp_comp_we g366 (.A(w447), .Z(w430), .nZ(w431) );
	vdp_comp_we g367 (.A(w447), .Z(w422), .nZ(w421) );
	vdp_comp_we g368 (.A(w447), .Z(w398), .nZ(w1567) );
	vdp_comp_we g369 (.A(w452), .Z(w6716), .nZ(w6717) );
	vdp_comp_we g370 (.A(w408), .Z(w399), .nZ(w400) );
	vdp_comp_we g371 (.A(w445), .Z(w1566), .nZ(w401) );
	vdp_and g372 (.Z(w411), .B(HCLK1), .A(w410) );
	vdp_and g373 (.Z(w412), .B(HCLK1), .A(w413) );
	vdp_and g374 (.Z(w416), .B(w420), .A(w418) );
	vdp_and g375 (.Z(w466), .B(w420), .A(w424) );
	vdp_nand g376 (.Z(w424), .B(w452), .A(w404) );
	vdp_nand g377 (.Z(w418), .B(w452), .A(w425) );
	vdp_and3 g378 (.Z(w452), .B(w438), .A(w406), .C(w439) );
	vdp_and3 g379 (.Z(w408), .B(w407), .A(w419), .C(128k) );
	vdp_not g380 (.A(128k), .nZ(w439) );
	vdp_sr_bit g381 (.D(w436), .C2(HCLK2), .C1(HCLK1), .Q(w435), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g382 (.D(w1443), .Q(w473), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g383 (.D(w1522), .C2(HCLK2), .C1(HCLK1), .Q(w499), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g384 (.A(w500), .nZ(w426) );
	vdp_fa g385 (.SUM(w460), .A(w499), .B(1'b0), .CI(w501) );
	vdp_not g386 (.A(w436), .nZ(w434) );
	vdp_not g387 (.A(M5), .nZ(w472) );
	vdp_not g388 (.A(w444), .nZ(w442) );
	vdp_not g389 (.A(w454), .nZ(w455) );
	vdp_not g390 (.A(w506), .nZ(w457) );
	vdp_not g391 (.A(w499), .nZ(w456) );
	vdp_slatch g392 (.Q(w493), .D(w497), .C(w479), .nC(w433) );
	vdp_slatch g393 (.Q(w1510), .D(w497), .C(w491), .nC(w463) );
	vdp_slatch g394 (.Q(w494), .D(w497), .C(w477), .nC(w449) );
	vdp_slatch g395 (.Q(w495), .D(w497), .C(w475), .nC(w446) );
	vdp_slatch g396 (.Q(w496), .D(w470), .C(w479), .nC(w433) );
	vdp_slatch g397 (.Q(w498), .D(w470), .C(w491), .nC(w463) );
	vdp_slatch g398 (.Q(w1509), .D(w470), .E(w477), .nE(w449) );
	vdp_slatch g399 (.Q(w492), .D(w470), .C(w475), .nC(w446) );
	vdp_slatch g400 (.Q(w484), .D(w471), .C(w479), .nC(w433) );
	vdp_slatch g401 (.Q(w478), .D(w471), .C(w491), .nC(w463) );
	vdp_slatch g402 (.Q(w482), .D(w471), .C(w477), .nC(w449) );
	vdp_slatch g403 (.Q(w485), .D(w471), .C(w475), .nC(w446) );
	vdp_comp_dff g404 (.D(w440), .C2(HCLK2), .C1(HCLK1), .Q(w436), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and g405 (.Z(w1443), .B(w434), .A(w435) );
	vdp_or g406 (.Z(w441), .B(w472), .A(w442) );
	vdp_or g407 (.Z(w445), .B(CA[0]), .A(w406) );
	vdp_and3 g408 (.Z(w448), .B(w500), .A(w456), .C(w506) );
	vdp_and3 g409 (.Z(w450), .B(w500), .A(w457), .C(w499) );
	vdp_and3 g410 (.Z(w451), .B(w456), .A(w457), .C(w500) );
	vdp_xor g411 (.Z(w453), .B(w504), .A(w503) );
	vdp_aon22 g412 (.Z(w447), .A1(w455), .A2(w504), .B1(w523), .B2(w454) );
	vdp_and3 g413 (.Z(w462), .B(w499), .A(w506), .C(w500) );
	vdp_comp_str g414 (.A(w508), .Z(w479), .nZ(w433) );
	vdp_comp_str g415 (.A(w458), .Z(w475), .nZ(w446) );
	vdp_comp_str g416 (.A(w467), .Z(w477), .nZ(w449) );
	vdp_comp_str g417 (.A(w464), .Z(w491), .nZ(w463) );
	vdp_nand g418 (.Z(w454), .B(w505), .A(w453) );
	vdp_and g419 (.Z(w1522), .B(w502), .A(w460) );
	vdp_aoi21 g420 (.Z(w444), .B(w443), .A1(HCLK1), .A2(w473) );
	vdp_nor g421 (.Z(w443), .B(w476), .A(w472) );
	vdp_nor g422 (.Z(w438), .B(w470), .A(w471) );
	vdp_not g423 (.A(w487), .nZ(w549) );
	vdp_not g424 (.A(w486), .nZ(w553) );
	vdp_nor g425 (.Z(w613), .A(w534), .B(w487) );
	vdp_or g426 (.A(w1442), .Z(w488), .B(w489) );
	vdp_comp_we g427 (.A(w587), .nZ(w480), .Z(w528) );
	vdp_aon22 g428 (.Z(w486), .A1(w528), .A2(w471), .B1(w480), .B2(w490) );
	vdp_aon22 g429 (.Z(w552), .A1(w528), .A2(w513), .B1(w480), .B2(w488) );
	vdp_aon22 g430 (.Z(w543), .A1(w528), .A2(w539), .B1(w480), .B2(w503) );
	vdp_aon22 g431 (.Z(w487), .A1(w528), .A2(w470), .B1(w480), .B2(w535) );
	vdp_aon22 g432 (.Z(w548), .A1(w528), .A2(w533), .B1(w480), .B2(w504) );
	vdp_aon22 g433 (.Z(w534), .A1(w528), .A2(w497), .B1(w480), .B2(w527) );
	vdp_and g434 (.Z(w547), .A(w526), .B(w525) );
	vdp_and g435 (.Z(w483), .A(w526), .B(w506) );
	vdp_and g436 (.Z(w1511), .A(w499), .B(w525) );
	vdp_and g437 (.Z(w481), .A(w499), .B(w506) );
	vdp_and g438 (.Z(w1444), .A(w502), .B(w521) );
	vdp_fa g439 (.SUM(w521), .A(w506), .B(w507), .CO(w501), .CI(w522) );
	vdp_sr_bit g440 (.D(w1444), .C2(HCLK2), .C1(HCLK1), .Q(w506), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g441 (.A(w524), .nZ(w1446) );
	vdp_not g442 (.A(w514), .nZ(w517) );
	vdp_and g443 (.Z(w507), .A(w582), .B(w1446) );
	vdp_and3 g444 (.Z(w464), .B(w515), .A(w514), .C(w518) );
	vdp_and3 g445 (.Z(w508), .B(w515), .A(w514), .C(w516) );
	vdp_xor g446 (.Z(w520), .A(w499), .B(w514) );
	vdp_not g447 (.A(w506), .nZ(w525) );
	vdp_not g448 (.A(w499), .nZ(w526) );
	vdp_not g449 (.A(w505), .nZ(w1445) );
	vdp_and5 g450 (.Z(w38), .A(w550), .B(w543), .C(w554), .D(w553), .E(w487) );
	vdp_and5 g451 (.Z(w37), .A(w550), .B(w548), .C(w554), .D(w553), .E(w487) );
	vdp_aon2222 g452 (.C2(w544), .B2(w542), .A2(w541), .C1(w1511), .B1(w483), .A1(w547), .Z(w489), .D2(w545), .D1(w481) );
	vdp_aon2222 g453 (.C2(w478), .B2(w482), .A2(w485), .C1(w1511), .B1(w483), .A1(w547), .Z(w490), .D2(w484), .D1(w481) );
	vdp_aon2222 g454 (.C2(w1457), .B2(w538), .A2(w1458), .C1(w1511), .B1(w483), .A1(w547), .Z(w503), .D2(w536), .D1(w481) );
	vdp_aon2222 g455 (.C2(w498), .B2(w1509), .A2(w492), .C1(w1511), .B1(w483), .A1(w547), .Z(w535), .D2(w496), .D1(w481) );
	vdp_aon2222 g456 (.C2(w1512), .B2(w532), .A2(w529), .C1(w1511), .B1(w483), .A1(w547), .Z(w504), .D2(w546), .D1(w481) );
	vdp_aon2222 g457 (.C2(w1510), .B2(w494), .A2(w495), .C1(w1511), .B1(w483), .A1(w547), .Z(w527), .D2(w493), .D1(w481) );
	vdp_nor g458 (.Z(w524), .A(w1445), .B(w453) );
	vdp_or g459 (.Z(w469), .B(w511), .A(w975) );
	vdp_cnt_bit g460 (.R(SYSRES), .Q(w514), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2), .CI(w512) );
	vdp_cnt_bit g461 (.R(SYSRES), .Q(w516), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2), .CI(w575), .CO(w512) );
	vdp_not g462 (.A(w516), .nZ(w518) );
	vdp_not g463 (.A(w1447), .nZ(w515) );
	vdp_and3 g464 (.Z(w458), .B(w515), .A(w517), .C(w518) );
	vdp_and3 g465 (.Z(w467), .B(w515), .A(w517), .C(w516) );
	vdp_xor g466 (.Z(w519), .A(w506), .B(w516) );
	vdp_fa g467 (.SUM(w1571), .A(w583), .B(w523), .CO(w522), .CI(1'b0) );
	vdp_and g468 (.Z(w583), .A(w524), .B(w582) );
	vdp_and g469 (.Z(w1456), .A(w502), .B(w1571) );
	vdp_sr_bit g470 (.D(w1456), .C2(HCLK2), .C1(HCLK1), .Q(w523), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g471 (.A(w1454), .nZ(w568) );
	vdp_comp_str g472 (.A(w458), .Z(w562), .nZ(w540) );
	vdp_comp_str g473 (.A(w467), .Z(w570), .nZ(w530) );
	vdp_comp_str g474 (.A(w464), .Z(w569), .nZ(w537) );
	vdp_comp_str g475 (.A(w508), .Z(w571), .nZ(w531) );
	vdp_slatch g476 (.Q(w546), .D(w533), .C(w571), .nC(w531) );
	vdp_slatch g477 (.Q(w1512), .D(w533), .C(w569), .nC(w537) );
	vdp_slatch g478 (.Q(w532), .D(w533), .C(w570), .nC(w530) );
	vdp_slatch g479 (.Q(w529), .D(w533), .C(w562), .nC(w540) );
	vdp_slatch g480 (.Q(w536), .D(w539), .C(w571), .nC(w531) );
	vdp_slatch g481 (.Q(w1457), .D(w539), .C(w569), .nC(w537) );
	vdp_slatch g482 (.Q(w538), .D(w539), .C(w570), .nC(w530) );
	vdp_slatch g483 (.Q(w1458), .D(w539), .C(w562), .nC(w540) );
	vdp_slatch g484 (.Q(w545), .D(w513), .C(w571), .nC(w531) );
	vdp_slatch g485 (.Q(w544), .D(w513), .C(w569), .nC(w537) );
	vdp_slatch g486 (.Q(w542), .D(w513), .C(w570), .nC(w530) );
	vdp_slatch g487 (.Q(w541), .D(w513), .C(w562), .nC(w540) );
	vdp_and5 g488 (.Z(w175), .A(w550), .B(w543), .C(w553), .D(w534), .E(w549) );
	vdp_and5 g489 (.Z(w174), .A(w550), .B(w548), .C(w553), .D(w534), .E(w549) );
	vdp_not g490 (.A(M5), .nZ(w1442) );
	vdp_not g491 (.A(w534), .nZ(w554) );
	vdp_not g492 (.A(w551), .nZ(w550) );
	vdp_oai21 g493 (.A1(w587), .Z(w551), .A2(w582), .B(w552) );
	vdp_and3 g494 (.Z(w573), .B(w582), .A(w505), .C(w523) );
	vdp_nor g495 (.Z(w1455), .A(w572), .B(w523) );
	vdp_nor g496 (.Z(w580), .A(w520), .B(w519) );
	vdp_aoi21 g497 (.A1(DCLK1), .Z(w1447), .A2(w511), .B(w574) );
	vdp_comb1 g498 (.Z(w1454), .A1(w582), .B(w584), .A2(w1455), .C(HCLK1) );
	vdp_not g499 (.A(w560), .nZ(w35) );
	vdp_not g500 (.A(w1514), .nZ(w555) );
	vdp_not g501 (.A(128k), .nZ(w558) );
	vdp_not g502 (.A(w557), .nZ(w133) );
	vdp_not g503 (.A(w1515), .nZ(w134) );
	vdp_not g504 (.A(w1516), .nZ(w556) );
	vdp_not g505 (.A(VRAMA[0]), .nZ(w1517) );
	vdp_not g506 (.A(w564), .nZ(w563) );
	vdp_not g507 (.A(w499), .nZ(w609) );
	vdp_not g508 (.A(w506), .nZ(w611) );
	vdp_not g509 (.A(w585), .nZ(w608) );
	vdp_not g510 (.A(w406), .nZ(w607) );
	vdp_not g511 (.A(128k), .nZ(w1521) );
	vdp_not g512 (.A(w523), .nZ(w603) );
	vdp_not g513 (.A(SYSRES), .nZ(w502) );
	vdp_not g514 (.A(w591), .nZ(w1449) );
	vdp_not g515 (.A(w34), .nZ(w1448) );
	vdp_not g516 (.A(w581), .nZ(w599) );
	vdp_not g517 (.A(w574), .nZ(w578) );
	vdp_not g518 (.A(w578), .nZ(w579) );
	vdp_sr_bit g519 (.D(w1450), .C2(HCLK2), .C1(HCLK1), .Q(w582), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g520 (.D(w1453), .Q(w587), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_slatch g521 (.Q(w459), .D(VRAMA[0]), .C(w599), .nC(w581) );
	vdp_and g522 (.A(w32), .Z(w1450), .B(w1449) );
	vdp_and g523 (.A(w1448), .Z(w500), .B(w3) );
	vdp_and g524 (.A(w3), .Z(w581), .B(HCLK1) );
	vdp_and g525 (.A(w591), .Z(w34), .B(w589) );
	vdp_and g526 (.A(w590), .Z(w36), .B(w591) );
	vdp_and g527 (.A(w590), .B(w573) );
	vdp_or g528 (.A(w577), .Z(w575), .B(w511) );
	vdp_or g529 (.A(w579), .Z(w946), .B(1'b0) );
	vdp_or g530 (.A(SYSRES), .Z(w601), .B(w594) );
	vdp_and g531 (.A(w582), .Z(w1451), .B(DMA_BUSY) );
	vdp_and g532 (.A(w613), .Z(w505), .B(w1520) );
	vdp_and g533 (.A(w1521), .Z(w1520), .B(w406) );
	vdp_or g534 (.A(w573), .Z(w606), .B(w572) );
	vdp_or g535 (.A(DMA_BUSY), .Z(w1518), .B(w567) );
	vdp_or g536 (.A(DMA_BUSY), .Z(w1519), .B(w566) );
	vdp_and g537 (.A(M5), .Z(w585), .B(REG_BUS[0]) );
	vdp_or g538 (.A(w543), .Z(w559), .B(w558) );
	vdp_and g539 (.A(w548), .Z(w1513), .B(128k) );
	vdp_aon22 g540 (.Z(w533), .A2(w1518), .B1(w607), .B2(w585), .A1(w406) );
	vdp_aon22 g541 (.Z(w539), .A2(w1519), .B1(w608), .B2(w607), .A1(w406) );
	vdp_and3 g542 (.A(w32), .Z(w1453), .B(w36), .C(w1452) );
	vdp_rs_ff g543 (.Q(w1452), .R(w601), .S(w1451) );
	vdp_oai21 g544 (.A1(VRAMA[0]), .Z(w564), .A2(128k), .B(w593) );
	vdp_oai21 g545 (.A1(128k), .Z(w1516), .A2(w1517), .B(w593) );
	vdp_aoi21 g546 (.A1(w548), .Z(w1515), .A2(w561), .B(w563) );
	vdp_aoi21 g547 (.A1(w543), .Z(w557), .A2(w561), .B(w556) );
	vdp_aoi21 g548 (.A1(w561), .Z(w1514), .A2(w559), .B(w593) );
	vdp_aoi21 g549 (.A1(w561), .Z(w560), .A2(w1513), .B(w593) );
	vdp_and4 g550 (.A(w550), .Z(w561), .B(w554), .C(w549), .D(w553) );
	vdp_not g551 (.A(w637), .nZ(w1441) );
	vdp_not g552 (.A(w649), .nZ(w648) );
	vdp_and3 g553 (.A(w603), .Z(w604), .B(w639), .C(w648) );
	vdp_and3 g554 (.A(w611), .Z(w626), .B(w614), .C(w609) );
	vdp_and3 g555 (.A(w506), .Z(w630), .B(w614), .C(w609) );
	vdp_and3 g556 (.A(w611), .Z(w619), .B(w614), .C(w499) );
	vdp_and3 g557 (.A(w506), .Z(w623), .B(w614), .C(w499) );
	vdp_or g558 (.A(w605), .Z(w636), .B(w638) );
	vdp_or g559 (.A(w605), .Z(w642), .B(w646) );
	vdp_or g560 (.A(w672), .Z(w592), .B(w645) );
	vdp_and3 g561 (.Z(w590), .B(DMA_BUSY), .A(w671), .C(w644) );
	vdp_or3 g562 (.Z(w596), .B(w587), .A(w593), .C(w643) );
	vdp_and g563 (.A(w597), .Z(w511), .B(w598) );
	vdp_and g564 (.A(w582), .Z(w614), .B(w603) );
	vdp_bufif0 g565 (.A(w595), .Z(VRAMA[8]), .nE(w650) );
	vdp_aoi221 g566 (.Z(w637), .A2(w604), .B1(w591), .B2(w580), .A1(w580), .C(SYSRES) );
	vdp_aon33 g567 (.Z(w1038), .A2(w580), .B1(w1551), .B2(w580), .A1(w647), .A3(w1551), .B3(w600) );
	vdp_not g568 (.A(w606), .nZ(w1469) );
	vdp_comp_str g569 (.A(w568), .Z(w1470), .nZ(w633) );
	vdp_not g570 (.A(w630), .nZ(w632) );
	vdp_comp_str g571 (.A(w467), .Z(w1472), .nZ(w1471) );
	vdp_not g572 (.A(w606), .nZ(w851) );
	vdp_comp_str g573 (.A(w568), .Z(w634), .nZ(w635) );
	vdp_not g574 (.A(w584), .nZ(w650) );
	vdp_not g575 (.A(w630), .nZ(w1552) );
	vdp_comp_str g576 (.A(w467), .Z(w1473), .nZ(w631) );
	vdp_not g577 (.A(w626), .nZ(w625) );
	vdp_comp_str g578 (.A(w458), .Z(w1474), .nZ(w1556) );
	vdp_not g579 (.A(w626), .nZ(w627) );
	vdp_comp_str g580 (.A(w508), .Z(w1475), .nZ(w624) );
	vdp_comp_str g581 (.A(w458), .Z(w628), .nZ(w629) );
	vdp_not g582 (.A(w619), .nZ(w616) );
	vdp_comp_str g583 (.A(w464), .Z(w617), .nZ(w618) );
	vdp_not g584 (.A(w619), .nZ(w850) );
	vdp_comp_str g585 (.A(w464), .Z(w1554), .nZ(w1555) );
	vdp_not g586 (.A(w623), .nZ(w620) );
	vdp_comp_str g587 (.A(w508), .Z(w621), .nZ(w622) );
	vdp_not g588 (.A(w623), .nZ(w1553) );
	vdp_sr_bit g589 (.D(w1441), .Q(w591), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g590 (.D(w639), .Q(w649), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g591 (.D(w582), .Q(w639), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g592 (.D(w1038), .Q(w647), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g593 (.D(w575), .Q(w600), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_not g594 (.A(SYSRES), .nZ(w1551) );
	vdp_not g595 (.A(w1523), .nZ(w643) );
	vdp_sr_bit g596 (.D(w597), .Q(w598), .C2(DCLK2), .C1(DCLK1), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_sr_bit g597 (.D(w588), .C2(HCLK2), .C1(HCLK1), .Q(w594), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_dlatch_inv g598 (.D(w597), .C(HCLK2), .Q(w1523), .nC(nHCLK2) );
	vdp_slatch g599 (.D(w661), .C(w617), .nC(w618), .nQ(w6732) );
	vdp_slatch g600 (.D(REG_BUS[7]), .C(w1554), .nC(w1555), .nQ(w6733) );
	vdp_slatch g601 (.D(w661), .C(w621), .nC(w622), .nQ(w6752) );
	vdp_slatch g602 (.D(REG_BUS[7]), .C(w1475), .nC(w624), .nQ(w6750) );
	vdp_slatch g603 (.D(w661), .C(w1474), .nC(w1556), .nQ(w6766) );
	vdp_slatch g604 (.D(REG_BUS[7]), .C(w628), .nC(w629), .nQ(w6768) );
	vdp_slatch g605 (.D(w661), .C(w1473), .nC(w631), .nQ(w6786) );
	vdp_slatch g606 (.D(REG_BUS[7]), .C(w1472), .nC(w1471), .nQ(w6784) );
	vdp_slatch g607 (.D(VRAMA[9]), .C(w1470), .nC(w633), .nQ(w6800) );
	vdp_slatch g608 (.D(VRAMA[7]), .C(w634), .nC(w635), .nQ(w6801) );
	vdp_notif0 g609 (.nZ(VRAMA[7]), .nE(w851), .A(w6801) );
	vdp_notif0 g610 (.nZ(VRAMA[9]), .nE(w1469), .A(w6800) );
	vdp_notif0 g611 (.nZ(VRAMA[7]), .nE(w632), .A(w6784) );
	vdp_notif0 g612 (.nZ(VRAMA[9]), .nE(w1552), .A(w6786) );
	vdp_notif0 g613 (.nZ(VRAMA[7]), .nE(w627), .A(w6768) );
	vdp_notif0 g614 (.nZ(VRAMA[9]), .nE(w620), .A(w6752) );
	vdp_notif0 g615 (.nZ(VRAMA[7]), .nE(w1553), .A(w6750) );
	vdp_notif0 g616 (.nZ(VRAMA[9]), .nE(w625), .A(w6766) );
	vdp_notif0 g617 (.nZ(VRAMA[9]), .nE(w616), .A(w6732) );
	vdp_notif0 g618 (.nZ(VRAMA[7]), .nE(w850), .A(w6733) );
	vdp_bufif0 g619 (.A(w661), .Z(VRAMA[9]), .nE(w650) );
	vdp_bufif0 g620 (.A(REG_BUS[7]), .Z(VRAMA[7]), .nE(w650) );
	vdp_bufif0 g621 (.A(w654), .Z(VRAMA[8]), .nE(w1505) );
	vdp_bufif0 g622 (.A(w654), .Z(CA[8]), .nE(w853) );
	vdp_bufif0 g623 (.A(w653), .Z(VRAMA[7]), .nE(w1503) );
	vdp_bufif0 g624 (.A(w653), .Z(CA[7]), .nE(w852) );
	vdp_slatch g625 (.Q(w671), .D(REG_BUS[7]), .nQ(w668), .C(w1596), .nC(w1597) );
	vdp_not g626 (.A(REG_BUS[0]), .nZ(w666) );
	vdp_not g627 (.A(REG_BUS[7]), .nZ(w673) );
	vdp_and3 g628 (.Z(w672), .B(w644), .A(w668), .C(DMA_BUSY) );
	vdp_nand g629 (.A(w664), .Z(w693), .B(w665) );
	vdp_cnt_bit_load g630 (.D(REG_BUS[0]), .nL(w1599), .L(w1608), .R(1'b0), .Q(w654), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w636), .CO(w658) );
	vdp_cnt_bit_load g631 (.D(REG_BUS[7]), .nL(w1440), .L(w807), .R(1'b0), .Q(w653), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w656), .CO(w638) );
	vdp_cnt_bit_load g632 (.D(w666), .nL(w1598), .L(w815), .R(1'b0), .Q(w664), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w642), .CO(w663) );
	vdp_cnt_bit_load g633 (.D(w673), .nL(w796), .L(w797), .R(1'b0), .Q(w667), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w669), .CO(w646) );
	vdp_slatch g634 (.D(w681), .C(w617), .nC(w618), .nQ(w6731) );
	vdp_slatch g635 (.D(REG_BUS[6]), .C(w1554), .nC(w1555), .nQ(w6734) );
	vdp_slatch g636 (.D(w681), .C(w621), .nC(w622), .nQ(w6751) );
	vdp_slatch g637 (.D(REG_BUS[6]), .C(w1475), .nC(w624), .nQ(w6749) );
	vdp_slatch g638 (.D(w681), .C(w1474), .nC(w1556), .nQ(w6765) );
	vdp_slatch g639 (.D(REG_BUS[6]), .C(w628), .nC(w629), .nQ(w6767) );
	vdp_slatch g640 (.D(w681), .C(w1473), .nC(w631), .nQ(w6785) );
	vdp_slatch g641 (.D(REG_BUS[6]), .C(w1472), .nC(w1471), .nQ(w6783) );
	vdp_slatch g642 (.D(VRAMA[10]), .C(w1470), .nC(w633), .nQ(w6799) );
	vdp_slatch g643 (.D(VRAMA[6]), .C(w634), .nC(w635), .nQ(w6802) );
	vdp_notif0 g644 (.nZ(VRAMA[6]), .nE(w851), .A(w6802) );
	vdp_notif0 g645 (.nZ(VRAMA[10]), .nE(w1469), .A(w6799) );
	vdp_notif0 g646 (.nZ(VRAMA[6]), .nE(w632), .A(w6783) );
	vdp_notif0 g647 (.nZ(VRAMA[10]), .nE(w1552), .A(w6785) );
	vdp_notif0 g648 (.nZ(VRAMA[6]), .nE(w627), .A(w6767) );
	vdp_notif0 g649 (.nZ(VRAMA[10]), .nE(w620), .A(w6751) );
	vdp_notif0 g650 (.nZ(VRAMA[6]), .nE(w1553), .A(w6749) );
	vdp_notif0 g651 (.nZ(VRAMA[10]), .nE(w625), .A(w6765) );
	vdp_notif0 g652 (.nZ(VRAMA[10]), .nE(w616), .A(w6731) );
	vdp_notif0 g653 (.nZ(VRAMA[6]), .nE(w850), .A(w6734) );
	vdp_bufif0 g654 (.A(w681), .Z(VRAMA[10]), .nE(w650) );
	vdp_bufif0 g655 (.A(REG_BUS[6]), .Z(VRAMA[6]), .nE(w1506) );
	vdp_bufif0 g656 (.A(w652), .Z(VRAMA[9]), .nE(w1505) );
	vdp_bufif0 g657 (.A(w652), .Z(CA[9]), .nE(w853) );
	vdp_bufif0 g658 (.A(w675), .Z(VRAMA[6]), .nE(w1503) );
	vdp_bufif0 g659 (.A(w675), .Z(CA[6]), .nE(w852) );
	vdp_slatch g660 (.Q(w688), .D(REG_BUS[6]), .nQ(w644), .C(w1596), .nC(w1597) );
	vdp_not g661 (.A(REG_BUS[1]), .nZ(w684) );
	vdp_not g662 (.A(REG_BUS[6]), .nZ(w686) );
	vdp_and3 g663 (.Z(w645), .B(DMA_BUSY), .A(w688), .C(w668) );
	vdp_cnt_bit_load g664 (.D(REG_BUS[1]), .nL(w1599), .L(w1608), .R(1'b0), .Q(w652), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w658), .CO(w677) );
	vdp_cnt_bit_load g665 (.D(REG_BUS[6]), .nL(w1440), .L(w807), .R(1'b0), .Q(w675), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w676), .CO(w656) );
	vdp_cnt_bit_load g666 (.D(w684), .nL(w1598), .L(w815), .R(1'b0), .Q(w665), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w663), .CO(w683) );
	vdp_cnt_bit_load g667 (.D(w686), .nL(w796), .L(w797), .R(1'b0), .Q(w685), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w689), .CO(w669) );
	vdp_nand3 g668 (.Z(w692), .B(w685), .A(w691), .C(w667) );
	vdp_slatch g669 (.D(w705), .C(w617), .nC(w618), .nQ(w6730) );
	vdp_slatch g670 (.D(REG_BUS[5]), .C(w1554), .nC(w1555), .nQ(w6735) );
	vdp_slatch g671 (.D(w705), .C(w621), .nC(w622), .nQ(w6753) );
	vdp_slatch g672 (.D(REG_BUS[5]), .C(w1475), .nC(w624), .nQ(w6748) );
	vdp_slatch g673 (.D(w705), .C(w1474), .nC(w1556), .nQ(w6764) );
	vdp_slatch g674 (.D(w705), .C(w1473), .nC(w631), .nQ(w6787) );
	vdp_slatch g675 (.D(REG_BUS[5]), .C(w1472), .nC(w1471), .nQ(w6782) );
	vdp_slatch g676 (.D(VRAMA[11]), .C(w1470), .nC(w633), .nQ(w6798) );
	vdp_slatch g677 (.D(VRAMA[5]), .C(w634), .nC(w635), .nQ(w6803) );
	vdp_notif0 g678 (.nZ(VRAMA[5]), .nE(w851), .A(w6803) );
	vdp_notif0 g679 (.nZ(VRAMA[11]), .nE(w1469), .A(w6798) );
	vdp_notif0 g680 (.nZ(VRAMA[5]), .nE(w632), .A(w6782) );
	vdp_notif0 g681 (.nZ(VRAMA[11]), .nE(w1552), .A(w6787) );
	vdp_notif0 g682 (.nZ(VRAMA[5]), .nE(w627), .A(w6769) );
	vdp_notif0 g683 (.nZ(VRAMA[11]), .nE(w620), .A(w6753) );
	vdp_notif0 g684 (.nZ(VRAMA[5]), .nE(w1553), .A(w6748) );
	vdp_notif0 g685 (.nZ(VRAMA[11]), .nE(w625), .A(w6764) );
	vdp_notif0 g686 (.nZ(VRAMA[11]), .nE(w616), .A(w6730) );
	vdp_notif0 g687 (.nZ(VRAMA[5]), .nE(w850), .A(w6735) );
	vdp_bufif0 g688 (.A(w705), .Z(VRAMA[11]), .nE(w650) );
	vdp_bufif0 g689 (.A(REG_BUS[5]), .Z(VRAMA[5]), .nE(w1506) );
	vdp_bufif0 g690 (.A(w674), .Z(VRAMA[10]), .nE(w1505) );
	vdp_bufif0 g691 (.A(w674), .Z(CA[10]), .nE(w853) );
	vdp_bufif0 g692 (.A(w707), .Z(VRAMA[5]), .nE(w1503) );
	vdp_bufif0 g693 (.A(w707), .Z(CA[5]), .nE(w852) );
	vdp_slatch g694 (.Q(CA[18]), .D(REG_BUS[2]), .C(w1596), .nC(w1597) );
	vdp_not g695 (.A(REG_BUS[2]), .nZ(w700) );
	vdp_not g696 (.A(REG_BUS[5]), .nZ(w699) );
	vdp_and3 g697 (.Z(w589), .B(DMA_BUSY), .A(w688), .C(w671) );
	vdp_cnt_bit_load g698 (.D(REG_BUS[2]), .nL(w1599), .L(w1608), .R(1'b0), .Q(w674), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w677), .CO(w710) );
	vdp_cnt_bit_load g699 (.D(REG_BUS[5]), .nL(w1440), .L(w807), .R(1'b0), .Q(w707), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w706), .CO(w676) );
	vdp_cnt_bit_load g700 (.D(w700), .nL(w1598), .L(w815), .R(1'b0), .Q(w690), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w683), .CO(w701) );
	vdp_cnt_bit_load g701 (.D(w699), .nL(w796), .L(w797), .R(1'b0), .Q(w691), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w696), .CO(w689) );
	vdp_nand3 g702 (.Z(w704), .B(w702), .A(w703), .C(w690) );
	vdp_slatch g703 (.D(w719), .C(w617), .nC(w618), .nQ(w6729) );
	vdp_slatch g704 (.D(REG_BUS[4]), .C(w1554), .nC(w1555), .nQ(w6736) );
	vdp_slatch g705 (.D(w719), .C(w621), .nC(w622), .nQ(w6754) );
	vdp_slatch g706 (.D(REG_BUS[4]), .C(w1475), .nC(w624), .nQ(w6747) );
	vdp_slatch g707 (.D(w719), .C(w1474), .nC(w1556), .nQ(w6763) );
	vdp_slatch g708 (.D(w719), .C(w1473), .nC(w631), .nQ(w6788) );
	vdp_slatch g709 (.D(REG_BUS[4]), .C(w1472), .nC(w1471), .nQ(w6781) );
	vdp_slatch g710 (.D(VRAMA[12]), .C(w1470), .nC(w633), .nQ(w6797) );
	vdp_slatch g711 (.D(VRAMA[4]), .C(w634), .nC(w635), .nQ(w6804) );
	vdp_notif0 g712 (.nZ(VRAMA[4]), .nE(w851), .A(w6804) );
	vdp_notif0 g713 (.nZ(VRAMA[12]), .nE(w1469), .A(w6797) );
	vdp_notif0 g714 (.nZ(VRAMA[4]), .nE(w632), .A(w6781) );
	vdp_notif0 g715 (.nZ(VRAMA[12]), .nE(w1552), .A(w6788) );
	vdp_notif0 g716 (.nZ(VRAMA[4]), .nE(w627), .A(w6770) );
	vdp_notif0 g717 (.nZ(VRAMA[12]), .nE(w620), .A(w6754) );
	vdp_notif0 g718 (.nZ(VRAMA[4]), .nE(w1553), .A(w6747) );
	vdp_notif0 g719 (.nZ(VRAMA[12]), .nE(w625), .A(w6763) );
	vdp_notif0 g720 (.nZ(VRAMA[12]), .nE(w616), .A(w6729) );
	vdp_notif0 g721 (.nZ(VRAMA[4]), .nE(w850), .A(w6736) );
	vdp_bufif0 g722 (.A(w719), .Z(VRAMA[12]), .nE(w650) );
	vdp_bufif0 g723 (.A(REG_BUS[4]), .Z(VRAMA[4]), .nE(w1506) );
	vdp_bufif0 g724 (.A(w709), .Z(VRAMA[11]), .nE(w1505) );
	vdp_bufif0 g725 (.A(w709), .Z(CA[11]), .nE(w853) );
	vdp_bufif0 g726 (.A(w720), .Z(VRAMA[4]), .nE(w1503) );
	vdp_bufif0 g727 (.A(w720), .Z(CA[4]), .nE(w852) );
	vdp_slatch g728 (.Q(CA[19]), .D(REG_BUS[3]), .C(w1596), .nC(w1597) );
	vdp_not g729 (.A(REG_BUS[3]), .nZ(w721) );
	vdp_not g730 (.A(REG_BUS[4]), .nZ(w723) );
	vdp_and g731 (.Z(w588), .B(w698), .A(w731) );
	vdp_cnt_bit_load g732 (.D(REG_BUS[3]), .nL(w1599), .L(w1608), .R(1'b0), .Q(w709), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w710), .CO(w715) );
	vdp_cnt_bit_load g733 (.D(REG_BUS[4]), .nL(w1440), .L(w807), .R(1'b0), .Q(w720), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w725), .CO(w706) );
	vdp_cnt_bit_load g734 (.D(w721), .nL(w1598), .L(w815), .R(1'b0), .Q(w702), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w701), .CO(w726) );
	vdp_cnt_bit_load g735 (.D(w723), .nL(w796), .L(w797), .R(1'b0), .Q(w729), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w730), .CO(w696) );
	vdp_nor3 g736 (.Z(w698), .B(w704), .A(w728), .C(w693) );
	vdp_slatch g737 (.D(w737), .C(w617), .nC(w618), .nQ(w6728) );
	vdp_slatch g738 (.D(REG_BUS[3]), .C(w1554), .nC(w1555), .nQ(w6737) );
	vdp_slatch g739 (.D(w737), .C(w621), .nC(w622), .nQ(w6755) );
	vdp_slatch g740 (.D(REG_BUS[3]), .C(w1475), .nC(w624), .nQ(w6746) );
	vdp_slatch g741 (.D(w737), .C(w1474), .nC(w1556), .nQ(w6762) );
	vdp_slatch g742 (.D(REG_BUS[3]), .C(w628), .nC(w629), .nQ(w6772) );
	vdp_slatch g743 (.D(w737), .C(w1473), .nC(w631), .nQ(w6790) );
	vdp_slatch g744 (.D(REG_BUS[3]), .C(w1472), .nC(w1471), .nQ(w6780) );
	vdp_slatch g745 (.D(VRAMA[13]), .C(w1470), .nC(w633), .nQ(w6796) );
	vdp_slatch g746 (.D(VRAMA[3]), .C(w634), .nC(w635), .nQ(w6805) );
	vdp_notif0 g747 (.nZ(VRAMA[3]), .nE(w851), .A(w6805) );
	vdp_notif0 g748 (.nZ(VRAMA[13]), .nE(w1469), .A(w6796) );
	vdp_notif0 g749 (.nZ(VRAMA[3]), .nE(w632), .A(w6780) );
	vdp_notif0 g750 (.nZ(VRAMA[13]), .nE(w1552), .A(w6790) );
	vdp_notif0 g751 (.nZ(VRAMA[3]), .nE(w627), .A(w6772) );
	vdp_notif0 g752 (.nZ(VRAMA[13]), .nE(w620), .A(w6755) );
	vdp_notif0 g753 (.nZ(VRAMA[3]), .nE(w1553), .A(w6746) );
	vdp_notif0 g754 (.nZ(VRAMA[13]), .nE(w625), .A(w6762) );
	vdp_notif0 g755 (.nZ(VRAMA[13]), .nE(w616), .A(w6728) );
	vdp_notif0 g756 (.nZ(VRAMA[3]), .nE(w850), .A(w6737) );
	vdp_bufif0 g757 (.A(w737), .Z(VRAMA[13]), .nE(w650) );
	vdp_bufif0 g758 (.A(REG_BUS[3]), .Z(VRAMA[3]), .nE(w1506) );
	vdp_bufif0 g759 (.A(w714), .Z(VRAMA[12]), .nE(w1505) );
	vdp_bufif0 g760 (.A(w714), .Z(CA[12]), .nE(w853) );
	vdp_bufif0 g761 (.A(w745), .Z(VRAMA[3]), .nE(w1503) );
	vdp_bufif0 g762 (.A(w745), .Z(CA[3]), .nE(w852) );
	vdp_slatch g763 (.Q(w752), .D(REG_BUS[4]), .C(w1596), .nC(w1597) );
	vdp_not g764 (.A(REG_BUS[4]), .nZ(w739) );
	vdp_not g765 (.A(REG_BUS[3]), .nZ(w740) );
	vdp_cnt_bit_load g766 (.D(REG_BUS[4]), .nL(w1599), .L(w1608), .R(1'b0), .Q(w714), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w715), .CO(w736) );
	vdp_cnt_bit_load g767 (.D(REG_BUS[3]), .nL(w1440), .L(w807), .R(1'b0), .Q(w745), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w734), .CO(w725) );
	vdp_cnt_bit_load g768 (.D(w739), .nL(w1598), .L(w815), .R(1'b0), .Q(w703), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w726), .CO(w744) );
	vdp_cnt_bit_load g769 (.D(w740), .nL(w796), .L(w797), .R(1'b0), .Q(w749), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w741), .CO(w730) );
	vdp_nor3 g770 (.Z(w731), .B(w750), .A(w748), .C(w692) );
	vdp_bufif0 g771 (.A(w752), .Z(CA[20]), .nE(w794) );
	vdp_slatch g772 (.D(w756), .C(w617), .nC(w618), .nQ(w6727) );
	vdp_slatch g773 (.D(REG_BUS[2]), .C(w1554), .nC(w1555), .nQ(w6738) );
	vdp_slatch g774 (.D(w756), .C(w621), .nC(w622), .nQ(w6756) );
	vdp_slatch g775 (.D(REG_BUS[2]), .C(w1475), .nC(w624), .nQ(w6745) );
	vdp_slatch g776 (.D(w756), .C(w1474), .nC(w1556), .nQ(w6761) );
	vdp_slatch g777 (.D(REG_BUS[2]), .C(w628), .nC(w629), .nQ(w6771) );
	vdp_slatch g778 (.D(w756), .C(w1473), .nC(w631), .nQ(w6789) );
	vdp_slatch g779 (.D(REG_BUS[2]), .C(w1472), .nC(w1471), .nQ(w6779) );
	vdp_slatch g780 (.D(VRAMA[14]), .C(w1470), .nC(w633), .nQ(w6795) );
	vdp_slatch g781 (.D(VRAMA[2]), .nC(w635), .C(w634), .nQ(w6806) );
	vdp_notif0 g782 (.nZ(VRAMA[2]), .nE(w851), .A(w6806) );
	vdp_notif0 g783 (.nZ(VRAMA[14]), .nE(w1469), .A(w6795) );
	vdp_notif0 g784 (.nZ(VRAMA[2]), .nE(w632), .A(w6779) );
	vdp_notif0 g785 (.nZ(VRAMA[14]), .nE(w1552), .A(w6789) );
	vdp_notif0 g786 (.nZ(VRAMA[2]), .nE(w627), .A(w6771) );
	vdp_notif0 g787 (.nZ(VRAMA[14]), .nE(w620), .A(w6756) );
	vdp_notif0 g788 (.nZ(VRAMA[2]), .nE(w1553), .A(w6745) );
	vdp_notif0 g789 (.nZ(VRAMA[14]), .nE(w625), .A(w6761) );
	vdp_notif0 g790 (.nZ(VRAMA[14]), .nE(w616), .A(w6727) );
	vdp_notif0 g791 (.nZ(VRAMA[2]), .nE(w850), .A(w6738) );
	vdp_bufif0 g792 (.A(w756), .Z(VRAMA[14]), .nE(w1504) );
	vdp_bufif0 g793 (.A(REG_BUS[2]), .Z(VRAMA[2]), .nE(w1506) );
	vdp_bufif0 g794 (.A(w735), .Z(VRAMA[13]), .nE(w1505) );
	vdp_bufif0 g795 (.A(w735), .Z(CA[13]), .nE(w853) );
	vdp_bufif0 g796 (.A(w757), .Z(VRAMA[2]), .nE(w1503) );
	vdp_bufif0 g797 (.A(w757), .Z(CA[2]), .nE(w852) );
	vdp_slatch g798 (.Q(w764), .D(REG_BUS[5]), .C(w1596), .nC(w1597) );
	vdp_not g799 (.A(REG_BUS[5]), .nZ(w758) );
	vdp_not g800 (.A(REG_BUS[2]), .nZ(w759) );
	vdp_cnt_bit_load g801 (.D(REG_BUS[5]), .nL(w1599), .L(w1608), .R(1'b0), .Q(w735), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w736), .CO(w770) );
	vdp_cnt_bit_load g802 (.D(REG_BUS[2]), .nL(w1440), .L(w807), .R(1'b0), .Q(w757), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w769), .CO(w734) );
	vdp_cnt_bit_load g803 (.D(w758), .nL(w1598), .L(w815), .R(1'b0), .Q(w768), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w744), .CO(w760) );
	vdp_cnt_bit_load g804 (.D(w759), .nL(w796), .L(w797), .R(1'b0), .Q(w766), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w772), .CO(w741) );
	vdp_nand3 g805 (.Z(w750), .B(w749), .A(w766), .C(w729) );
	vdp_bufif0 g806 (.A(w764), .Z(CA[21]), .nE(w794) );
	vdp_slatch g807 (.D(w777), .C(w617), .nC(w618), .nQ(w6726) );
	vdp_slatch g808 (.D(REG_BUS[1]), .C(w1554), .nC(w1555), .nQ(w6739) );
	vdp_slatch g809 (.D(w777), .C(w621), .nC(w622), .nQ(w6758) );
	vdp_slatch g810 (.D(REG_BUS[1]), .C(w1475), .nC(w624), .nQ(w6744) );
	vdp_slatch g811 (.D(w777), .C(w1474), .nC(w1556), .nQ(w6760) );
	vdp_slatch g812 (.D(REG_BUS[1]), .C(w628), .nC(w629), .nQ(w6774) );
	vdp_slatch g813 (.D(w777), .C(w1473), .nC(w631), .nQ(w6791) );
	vdp_slatch g814 (.D(REG_BUS[1]), .C(w1472), .nC(w1471), .nQ(w6778) );
	vdp_slatch g815 (.D(VRAMA[15]), .C(w1470), .nC(w633), .nQ(w6794) );
	vdp_slatch g816 (.D(VRAMA[1]), .C(w634), .nC(w635), .nQ(w6807) );
	vdp_notif0 g817 (.nZ(VRAMA[1]), .nE(w851), .A(w6807) );
	vdp_notif0 g818 (.nZ(VRAMA[15]), .nE(w1469), .A(w6794) );
	vdp_notif0 g819 (.nZ(VRAMA[1]), .nE(w632), .A(w6778) );
	vdp_notif0 g820 (.nZ(VRAMA[15]), .nE(w1552), .A(w6791) );
	vdp_notif0 g821 (.nZ(VRAMA[1]), .nE(w627), .A(w6774) );
	vdp_notif0 g822 (.nZ(VRAMA[15]), .nE(w620), .A(w6758) );
	vdp_notif0 g823 (.nZ(VRAMA[1]), .nE(w1553), .A(w6744) );
	vdp_notif0 g824 (.nZ(VRAMA[15]), .nE(w625), .A(w6760) );
	vdp_notif0 g825 (.nZ(VRAMA[15]), .nE(w616), .A(w6726) );
	vdp_notif0 g826 (.nZ(VRAMA[1]), .nE(w850), .A(w6739) );
	vdp_bufif0 g827 (.A(w777), .Z(VRAMA[15]), .nE(w1504) );
	vdp_bufif0 g828 (.A(REG_BUS[1]), .Z(VRAMA[1]), .nE(w1506) );
	vdp_bufif0 g829 (.A(w753), .Z(VRAMA[14]), .nE(w1505) );
	vdp_bufif0 g830 (.A(w753), .Z(CA[14]), .nE(w853) );
	vdp_bufif0 g831 (.A(w779), .Z(VRAMA[1]), .nE(w1503) );
	vdp_bufif0 g832 (.A(w779), .Z(CA[1]), .nE(w852) );
	vdp_slatch g833 (.Q(w1507), .D(REG_BUS[1]), .C(w1596), .nC(w1597) );
	vdp_not g834 (.A(REG_BUS[6]), .nZ(w782) );
	vdp_not g835 (.A(REG_BUS[1]), .nZ(w785) );
	vdp_cnt_bit_load g836 (.D(REG_BUS[6]), .nL(w1599), .L(w1608), .R(1'b0), .Q(w753), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w770), .CO(w786) );
	vdp_cnt_bit_load g837 (.D(REG_BUS[1]), .nL(w1440), .L(w807), .R(1'b0), .Q(w779), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w787), .CO(w769) );
	vdp_cnt_bit_load g838 (.D(w782), .nL(w1598), .L(w815), .R(1'b0), .Q(w767), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w760), .CO(w780) );
	vdp_cnt_bit_load g839 (.D(w785), .nL(w796), .L(w797), .R(1'b0), .Q(w784), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w783), .CO(w772) );
	vdp_nand3 g840 (.Z(w728), .B(w767), .A(w768), .C(w781) );
	vdp_bufif0 g841 (.A(w1507), .Z(CA[17]), .nE(w794) );
	vdp_slatch g842 (.nQ(w778), .D(w791), .C(w617), .nC(w618) );
	vdp_slatch g843 (.D(REG_BUS[0]), .C(w1554), .nC(w1555), .nQ(w6740) );
	vdp_slatch g844 (.D(w791), .C(w621), .nC(w622), .nQ(w6757) );
	vdp_slatch g845 (.D(REG_BUS[0]), .C(w1475), .nC(w624), .nQ(w6743) );
	vdp_slatch g846 (.D(w791), .C(w1474), .nC(w1556), .nQ(w6759) );
	vdp_slatch g847 (.D(REG_BUS[0]), .C(w628), .nC(w629), .nQ(w6773) );
	vdp_slatch g848 (.D(w791), .C(w1473), .nC(w631), .nQ(w6792) );
	vdp_slatch g849 (.D(REG_BUS[0]), .C(w1472), .nC(w1471), .nQ(w6777) );
	vdp_slatch g850 (.D(VRAMA[16]), .C(w1470), .nC(w633), .nQ(w6793) );
	vdp_slatch g851 (.Q(w6808), .D(VRAMA[0]), .C(w634), .nC(w635) );
	vdp_notif0 g852 (.nZ(VRAMA[0]), .nE(w851), .A(w6808) );
	vdp_notif0 g853 (.nZ(VRAMA[16]), .nE(w1469), .A(w6793) );
	vdp_notif0 g854 (.nZ(VRAMA[0]), .nE(w632), .A(w6777) );
	vdp_notif0 g855 (.nZ(VRAMA[16]), .nE(w1552), .A(w6792) );
	vdp_notif0 g856 (.nZ(VRAMA[0]), .nE(w627), .A(w6773) );
	vdp_notif0 g857 (.nZ(VRAMA[16]), .nE(w620), .A(w6757) );
	vdp_notif0 g858 (.nZ(VRAMA[0]), .nE(w1553), .A(w6743) );
	vdp_notif0 g859 (.nZ(VRAMA[16]), .nE(w625), .A(w6759) );
	vdp_notif0 g860 (.A(w778), .nZ(VRAMA[16]), .nE(w616) );
	vdp_notif0 g861 (.nZ(VRAMA[0]), .nE(w850), .A(w6740) );
	vdp_bufif0 g862 (.A(w791), .Z(VRAMA[16]), .nE(w1504) );
	vdp_bufif0 g863 (.A(REG_BUS[0]), .Z(VRAMA[0]), .nE(w1506) );
	vdp_bufif0 g864 (.A(w773), .Z(VRAMA[15]), .nE(w1505) );
	vdp_bufif0 g865 (.A(w773), .Z(CA[15]), .nE(w853) );
	vdp_bufif0 g866 (.A(w801), .Z(VRAMA[0]), .nE(w1503) );
	vdp_bufif0 g867 (.A(w801), .Z(CA[0]), .nE(w852) );
	vdp_slatch g868 (.Q(w792), .D(REG_BUS[0]), .C(w1596), .nC(w1597) );
	vdp_not g869 (.A(REG_BUS[7]), .nZ(w1600) );
	vdp_not g870 (.A(REG_BUS[0]), .nZ(w1477) );
	vdp_cnt_bit_load g871 (.D(REG_BUS[7]), .nL(w1599), .L(w1608), .R(1'b0), .Q(w773), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w786) );
	vdp_cnt_bit_load g872 (.D(REG_BUS[0]), .nL(w1440), .L(w807), .R(1'b0), .Q(w801), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w799), .CO(w787) );
	vdp_cnt_bit_load g873 (.D(w1600), .nL(w1598), .L(w815), .R(1'b0), .Q(w781), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w780) );
	vdp_cnt_bit_load g874 (.D(w1477), .nL(w796), .L(w797), .R(1'b0), .Q(w1476), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w799), .CO(w783) );
	vdp_nand3 g875 (.Z(w748), .B(w784), .A(w596), .C(w1435) );
	vdp_bufif0 g876 (.A(w792), .Z(CA[16]), .nE(w794) );
	vdp_slatch g877 (.D(VRAMA[8]), .C(w634), .nC(w635), .nQ(w6809) );
	vdp_slatch g878 (.D(w595), .C(w1472), .nC(w1471), .nQ(w6776) );
	vdp_slatch g879 (.D(w595), .C(w628), .nC(w629), .nQ(w6775) );
	vdp_slatch g880 (.D(w595), .C(w1475), .nC(w624), .nQ(w6742) );
	vdp_slatch g881 (.D(w595), .C(w1554), .nC(w1555), .nQ(w6741) );
	vdp_notif0 g882 (.nZ(VRAMA[8]), .nE(w850), .A(w6741) );
	vdp_notif0 g883 (.nZ(VRAMA[8]), .nE(w1553), .A(w6742) );
	vdp_notif0 g884 (.nZ(VRAMA[8]), .nE(w627), .A(w6775) );
	vdp_notif0 g885 (.nZ(VRAMA[8]), .nE(w632), .A(w6776) );
	vdp_notif0 g886 (.nZ(VRAMA[8]), .nE(w851), .A(w6809) );
	vdp_bufif0 g887 (.A(w792), .Z(VRAMA[16]), .nE(w1505) );
	vdp_not g888 (.A(w1468), .nZ(w1504) );
	vdp_not g889 (.A(w584), .nZ(w1506) );
	vdp_not g890 (.A(w33), .nZ(w1505) );
	vdp_not g891 (.A(w592), .nZ(w853) );
	vdp_not g892 (.A(w33), .nZ(w1503) );
	vdp_not g893 (.A(w592), .nZ(w852) );
	vdp_not g894 (.A(w592), .nZ(w794) );
	vdp_not g895 (.A(w1476), .nZ(w1435) );
	vdp_not g896 (.A(w795), .nZ(w1439) );
	vdp_not g897 (.A(M5), .nZ(w812) );
	vdp_and4 g898 (.Z(w808), .B(w681), .A(w817), .D(w595), .C(w818) );
	vdp_and4 g899 (.Z(w809), .B(w681), .A(w817), .D(w820), .C(w661) );
	vdp_and4 g900 (.B(w821), .A(w802), .D(w820), .C(w818), .Z(w811) );
	vdp_and4 g901 (.B(w821), .A(w802), .D(w595), .C(w818), .Z(w810) );
	vdp_and4 g902 (.Z(w805), .B(w818), .A(w595), .D(w822), .C(w681) );
	vdp_and4 g903 (.Z(w803), .B(w661), .A(w820), .D(w802), .C(w821) );
	vdp_and4 g904 (.Z(w804), .B(w661), .A(w595), .D(w822), .C(w681) );
	vdp_and4 g905 (.B(w825), .A(M5), .D(w705), .C(w826), .Z(w817) );
	vdp_comp_str g906 (.A(w828), .Z(w1596), .nZ(w1597) );
	vdp_comp_we g907 (.A(w1481), .Z(w1608), .nZ(w1599) );
	vdp_comp_we g908 (.A(w806), .Z(w807), .nZ(w1440) );
	vdp_comp_we g909 (.A(w829), .Z(w815), .nZ(w1598) );
	vdp_comp_we g910 (.A(w830), .Z(w797), .nZ(w796) );
	vdp_and g911 (.Z(w605), .B(w596), .A(w795) );
	vdp_and g912 (.Z(w799), .B(w596), .A(w1439) );
	vdp_or g913 (.Z(w828), .B(w804), .A(SYSRES) );
	vdp_or g914 (.Z(w806), .B(w805), .A(SYSRES) );
	vdp_or g915 (.Z(w1468), .B(w812), .A(w584) );
	vdp_or g916 (.B(w810), .A(SYSRES), .Z(w87) );
	vdp_or g917 (.B(w811), .A(SYSRES), .Z(w86) );
	vdp_or g918 (.Z(w85), .B(w809), .A(SYSRES) );
	vdp_or g919 (.Z(w68), .B(w808), .A(SYSRES) );
	vdp_or g920 (.B(w1478), .A(SYSRES), .Z(w72) );
	vdp_and4 g921 (.B(w681), .A(w819), .D(w595), .C(w661), .Z(w837) );
	vdp_or g922 (.B(w837), .A(SYSRES), .Z(w73) );
	vdp_and4 g923 (.B(w821), .A(w822), .D(w820), .C(w661), .Z(w836) );
	vdp_or g924 (.B(w836), .A(SYSRES), .Z(w75) );
	vdp_and4 g925 (.B(w821), .A(w822), .D(w595), .C(w818), .Z(w835) );
	vdp_or g926 (.B(w835), .A(SYSRES), .Z(w74) );
	vdp_and4 g927 (.B(w821), .A(w822), .D(w820), .C(w818), .Z(w1479) );
	vdp_or g928 (.B(w1479), .A(SYSRES), .Z(w69) );
	vdp_and4 g929 (.B(w681), .A(w819), .D(w820), .C(w661), .Z(w834) );
	vdp_or g930 (.B(w834), .A(SYSRES), .Z(w143) );
	vdp_and4 g931 (.B(w681), .A(w819), .D(w595), .C(w818), .Z(w833) );
	vdp_or g932 (.B(w833), .A(SYSRES), .Z(w142) );
	vdp_or g933 (.B(w838), .A(SYSRES), .Z(w71) );
	vdp_and4 g934 (.B(w681), .A(w819), .D(w820), .C(w818), .Z(w1478) );
	vdp_or g935 (.B(w839), .A(SYSRES), .Z(w70) );
	vdp_and4 g936 (.B(w821), .A(w819), .D(w595), .C(w661), .Z(w838) );
	vdp_and4 g937 (.B(w821), .A(w819), .D(w820), .C(w661), .Z(w839) );
	vdp_and4 g938 (.B(w818), .A(w595), .D(w819), .C(w821), .Z(w841) );
	vdp_or g939 (.B(w841), .A(SYSRES), .Z(w1137) );
	vdp_and4 g940 (.B(w818), .A(w820), .D(w819), .C(w821), .Z(w1480) );
	vdp_or g941 (.B(w1480), .A(SYSRES), .Z(w1176) );
	vdp_and4 g942 (.B(w818), .A(w820), .D(w817), .C(w681), .Z(w840) );
	vdp_or g943 (.B(w840), .A(SYSRES), .Z(w1138) );
	vdp_and4 g944 (.B(w661), .A(w820), .D(w822), .C(w681), .Z(w842) );
	vdp_or g945 (.B(w842), .A(SYSRES), .Z(w1481) );
	vdp_and4 g946 (.B(w661), .A(w595), .D(w817), .C(w821), .Z(w1482) );
	vdp_or g947 (.B(w1482), .A(SYSRES), .Z(CA[14]) );
	vdp_and4 g948 (.B(w818), .A(w820), .D(w822), .C(w681), .Z(w843) );
	vdp_or g949 (.B(w843), .A(SYSRES), .Z(w829) );
	vdp_and4 g950 (.B(w661), .A(w595), .D(w822), .C(w821), .Z(w844) );
	vdp_or g951 (.B(w844), .A(SYSRES), .Z(w830) );
	vdp_and4 g952 (.B(w661), .A(w831), .D(w817), .C(w681), .Z(w845) );
	vdp_or g953 (.B(w845), .A(SYSRES), .Z(w846) );
	vdp_and4 g954 (.B(w827), .A(w825), .D(M5), .C(w719), .Z(w822) );
	vdp_and3 g955 (.B(w826), .A(w825), .C(w705), .Z(w802) );
	vdp_and3 g956 (.B(w827), .A(w825), .C(w826), .Z(w819) );
	vdp_or g957 (.Z(w847), .B(w848), .A(w6711) );
	vdp_and g958 (.B(w824), .A(HCLK1), .Z(w825) );
	vdp_dlatch_inv g959 (.D(w823), .C(DCLK2), .nQ(w848), .nC(nDCLK2) );
	vdp_dlatch_inv g960 (.D(w6710), .C(HCLK2), .nQ(w824), .nC(nHCLK2) );
	vdp_not g961 (.A(w719), .nZ(w826) );
	vdp_not g962 (.A(w705), .nZ(w827) );
	vdp_not g963 (.A(w661), .nZ(w818) );
	vdp_not g964 (.A(w681), .nZ(w821) );
	vdp_not g965 (.A(w595), .nZ(w820) );
	vdp_slatch g966 (.D(REG_BUS[5]), .C(w628), .nC(w629), .nQ(w6769) );
	vdp_slatch g967 (.D(REG_BUS[4]), .C(w628), .nC(w629), .nQ(w6770) );
	vdp_sr_bit g968 (.D(w848), .C2(DCLK2), .C1(DCLK1), .Q(w6711), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_dlatch_inv g969 (.D(w847), .C(DCLK1), .nQ(w6710), .nC(nDCLK1) );
	vdp_comp_str g970 (.A(w885), .Z(w855), .nZ(w863) );
	vdp_fa g971 (.SUM(w882), .A(REG_BUS[6]), .B(w1573), .CO(w884), .CI(w880) );
	vdp_fa g972 (.SUM(w878), .A(REG_BUS[5]), .B(w879), .CO(w880), .CI(w877) );
	vdp_fa g973 (.SUM(w875), .A(REG_BUS[4]), .B(w876), .CO(w877), .CI(w872) );
	vdp_fa g974 (.SUM(w871), .A(REG_BUS[3]), .B(w874), .CO(w872), .CI(w869) );
	vdp_fa g975 (.SUM(w867), .A(REG_BUS[2]), .B(w868), .CO(w869), .CI(w866) );
	vdp_fa g976 (.SUM(w6714), .A(REG_BUS[1]), .B(w865), .CO(w866), .CI(w862) );
	vdp_fa g977 (.SUM(w6715), .A(REG_BUS[0]), .B(w859), .CO(w862), .CI(w857) );
	vdp_fa g978 (.SUM(w1483), .A(REG_BUS[7]), .B(w1572), .CO(w886), .CI(w884) );
	vdp_slatch g979 (.Q(w883), .D(DB[7]), .C(w855), .nC(w863) );
	vdp_aon22 g980 (.Z(w1583), .A1(w883), .A2(w854), .B1(w860), .B2(w1483) );
	vdp_slatch g981 (.Q(w881), .D(DB[6]), .C(w855), .nC(w863) );
	vdp_aon22 g982 (.Z(w1584), .A1(w881), .A2(w854), .B1(w860), .B2(w882) );
	vdp_slatch g983 (.Q(w1526), .D(DB[5]), .C(w855), .nC(w863) );
	vdp_aon22 g984 (.Z(w1585), .A1(w1526), .A2(w854), .B1(w860), .B2(w878) );
	vdp_slatch g985 (.Q(w873), .D(DB[4]), .C(w855), .nC(w863) );
	vdp_aon22 g986 (.Z(w1586), .A1(w873), .A2(w854), .B1(w860), .B2(w875) );
	vdp_slatch g987 (.Q(w870), .D(DB[3]), .C(w855), .nC(w863) );
	vdp_aon22 g988 (.Z(w1587), .A1(w870), .A2(w854), .B1(w860), .B2(w871) );
	vdp_slatch g989 (.Q(w864), .D(DB[2]), .C(w855), .nC(w863) );
	vdp_aon22 g990 (.Z(w1588), .A1(w864), .A2(w854), .B1(w860), .B2(w867) );
	vdp_slatch g991 (.Q(w861), .D(DB[1]), .C(w855), .nC(w863) );
	vdp_aon22 g992 (.Z(w1589), .A1(w861), .A2(w854), .B1(w860), .B2(w6714) );
	vdp_slatch g993 (.Q(w856), .D(DB[0]), .C(w855), .nC(w863) );
	vdp_aon22 g994 (.Z(w1590), .A1(w856), .A2(w854), .B1(w860), .B2(w6715) );
	vdp_dff g995 (.Q(REG_BUS[0]), .R(SYSRES), .C(w888), .D(w1590) );
	vdp_slatch g996 (.Q(w859), .D(REG_BUS[0]), .C(w887), .nC(w858) );
	vdp_dff g997 (.Q(REG_BUS[1]), .R(SYSRES), .D(w1589), .C(w888) );
	vdp_slatch g998 (.Q(w865), .D(REG_BUS[1]), .C(w887), .nC(w858) );
	vdp_dff g999 (.Q(REG_BUS[2]), .R(SYSRES), .C(w888), .D(w1588) );
	vdp_slatch g1000 (.Q(w868), .D(REG_BUS[2]), .C(w887), .nC(w858) );
	vdp_dff g1001 (.Q(REG_BUS[3]), .R(SYSRES), .D(w1587), .C(w888) );
	vdp_slatch g1002 (.Q(w874), .D(REG_BUS[3]), .C(w887), .nC(w858) );
	vdp_dff g1003 (.Q(REG_BUS[4]), .R(SYSRES), .C(w888), .D(w1586) );
	vdp_slatch g1004 (.Q(w876), .D(REG_BUS[4]), .C(w887), .nC(w858) );
	vdp_dff g1005 (.Q(REG_BUS[5]), .R(SYSRES), .C(w888), .D(w1585) );
	vdp_slatch g1006 (.Q(w879), .D(REG_BUS[5]), .C(w887), .nC(w858) );
	vdp_dff g1007 (.Q(REG_BUS[6]), .R(SYSRES), .C(w888), .D(w1584) );
	vdp_slatch g1008 (.Q(w1573), .D(REG_BUS[6]), .C(w887), .nC(w858) );
	vdp_dff g1009 (.Q(REG_BUS[7]), .R(SYSRES), .D(w1583), .C(w888) );
	vdp_slatch g1010 (.Q(w1572), .D(REG_BUS[7]), .C(w887), .nC(w858) );
	vdp_comp_str g1011 (.A(w846), .Z(w887), .nZ(w858) );
	vdp_comp_we g1012 (.A(w891), .Z(w854), .nZ(w860) );
	vdp_dff g1013 (.Q(w791), .R(w895), .C(w888), .D(w1574) );
	vdp_dff g1014 (.Q(w777), .R(w895), .C(w888), .D(w1575) );
	vdp_dff g1015 (.Q(w756), .R(w895), .C(w888), .D(w1576) );
	vdp_dff g1016 (.Q(w737), .R(SYSRES), .C(w888), .D(w1577) );
	vdp_dff g1017 (.Q(w719), .R(SYSRES), .C(w888), .D(w1578) );
	vdp_dff g1018 (.Q(w705), .R(SYSRES), .C(w888), .D(w1579) );
	vdp_dff g1019 (.Q(w681), .R(SYSRES), .C(w888), .D(w1580) );
	vdp_dff g1020 (.Q(w661), .R(SYSRES), .C(w888), .D(w1581) );
	vdp_dff g1021 (.Q(w595), .R(SYSRES), .C(w888), .D(w1582) );
	vdp_not g1022 (.A(w917), .nZ(w888) );
	vdp_or g1023 (.Z(w895), .B(SYSRES), .A(w857) );
	vdp_not g1024 (.A(M5), .nZ(w857) );
	vdp_slatch g1025 (.Q(w914), .D(w929), .C(w928), .nC(w905) );
	vdp_aon22 g1026 (.Z(w1582), .A1(w918), .A2(w926), .B1(w892), .B2(w916) );
	vdp_slatch g1027 (.Q(w918), .D(w245), .C(w928), .nC(w905) );
	vdp_comp_str g1028 (.A(w933), .Z(w928), .nZ(w905) );
	vdp_comp_we g1029 (.A(w891), .Z(w926), .nZ(w892) );
	vdp_ha g1030 (.SUM(w916), .A(w595), .B(w886), .CO(w913) );
	vdp_slatch g1031 (.Q(w912), .D(w253), .C(w928), .nC(w905) );
	vdp_aon22 g1032 (.Z(w1581), .A1(w914), .A2(w926), .B1(w892), .B2(w915) );
	vdp_ha g1033 (.SUM(w915), .A(w661), .B(w913), .CO(w1593) );
	vdp_slatch g1034 (.Q(w910), .D(w289), .C(w928), .nC(w905) );
	vdp_aon22 g1035 (.Z(w1580), .A1(w912), .A2(w926), .B1(w892), .B2(w911) );
	vdp_ha g1036 (.SUM(w911), .A(w681), .B(w1593), .CO(w909) );
	vdp_slatch g1037 (.Q(w907), .D(w262), .C(w928), .nC(w905) );
	vdp_aon22 g1038 (.Z(w1579), .A1(w910), .A2(w926), .B1(w892), .B2(w908) );
	vdp_ha g1039 (.SUM(w908), .A(w705), .B(w909), .CO(w1592) );
	vdp_slatch g1040 (.Q(w904), .D(w299), .C(w928), .nC(w905) );
	vdp_aon22 g1041 (.Z(w1578), .A1(w907), .A2(w926), .B1(w892), .B2(w906) );
	vdp_ha g1042 (.SUM(w906), .A(w719), .B(w1592), .CO(w903) );
	vdp_aon22 g1043 (.Z(w1577), .A1(w904), .A2(w926), .B1(w892), .B2(w901) );
	vdp_ha g1044 (.SUM(w901), .A(w737), .B(w903), .CO(w902) );
	vdp_comp_str g1045 (.A(w927), .Z(w925), .nZ(w894) );
	vdp_aon22 g1046 (.Z(w1576), .A1(w900), .A2(w926), .B1(w892), .B2(w1591) );
	vdp_ha g1047 (.SUM(w1591), .A(w756), .B(w902), .CO(w897) );
	vdp_slatch_r g1048 (.Q(w900), .D(DB[0]), .R(w895), .C(w925), .nC(w894) );
	vdp_slatch_r g1049 (.Q(w899), .D(DB[1]), .R(w895), .C(w925), .nC(w894) );
	vdp_aon22 g1050 (.Z(w1575), .A1(w899), .A2(w926), .B1(w892), .B2(w898) );
	vdp_ha g1051 (.SUM(w898), .A(w777), .B(w897), .CO(w896) );
	vdp_slatch_r g1052 (.Q(w893), .D(DB[2]), .R(w895), .C(w925), .nC(w894) );
	vdp_aon22 g1053 (.Z(w1574), .A1(w893), .A2(w926), .B1(w892), .B2(w1525) );
	vdp_ha g1054 (.SUM(w1525), .A(w791), .B(w896) );
	vdp_and3 g1055 (.C(w922), .A(w920), .B(w921), .Z(w924) );
	vdp_sr_bit g1056 (.D(w1489), .C2(HCLK2), .C1(HCLK1), .nQ(w110), .nC1(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1057 (.D(w942), .Q(w1489), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK2), .nC1(nHCLK1) );
	vdp_not g1058 (.A(w969), .nZ(w944) );
	vdp_not g1059 (.A(w470), .nZ(w1490) );
	vdp_not g1060 (.A(w471), .nZ(w955) );
	vdp_not g1061 (.A(w920), .nZ(w956) );
	vdp_not g1062 (.A(w953), .nZ(w961) );
	vdp_not g1063 (.A(w513), .nZ(w938) );
	vdp_not g1064 (.A(w589), .nZ(w950) );
	vdp_not g1065 (.A(w976), .nZ(w964) );
	vdp_not g1066 (.A(w1491), .nZ(w967) );
	vdp_not g1067 (.A(w965), .nZ(w934) );
	vdp_slatch g1068 (.Q(w497), .D(w931), .C(w932), .nC(w945) );
	vdp_slatch g1069 (.Q(w513), .D(w271), .C(w932), .nC(w945) );
	vdp_comp_str g1070 (.A(w933), .Z(w932), .nZ(w945) );
	vdp_dlatch_inv g1071 (.D(w597), .C(DCLK1), .nQ(w965), .nC(nDCLK1) );
	vdp_dlatch_inv g1072 (.D(w964), .C(DCLK1), .nQ(w963), .nC(nDCLK1) );
	vdp_dlatch_inv g1073 (.D(w978), .C(DCLK2), .nQ(w976), .nC(nDCLK2) );
	vdp_dlatch_inv g1074 (.D(w983), .C(DCLK1), .nQ(w978), .nC(nDCLK1) );
	vdp_slatch g1075 (.Q(w983), .D(w940), .C(DCLK2), .nC(nDCLK2) );
	vdp_slatch g1076 (.Q(w940), .D(w977), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g1077 (.D(w584), .C(HCLK1), .nQ(w939), .nC(nHCLK1) );
	vdp_rs_FF g1078 (.nQ(w936), .R(w985), .S(w984), .Q(w948) );
	vdp_rs_FF g1079 (.Q(w960), .R(w958), .S(w937) );
	vdp_and3 g1080 (.C(w423), .A(w471), .B(w1490), .Z(w943) );
	vdp_and3 g1081 (.C(w955), .A(w470), .B(w423), .Z(w109) );
	vdp_comp_dff g1082 (.D(w959), .C2(HCLK2), .C1(HCLK1), .Q(w952), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_comp_dff g1083 (.D(w949), .C2(HCLK2), .C1(HCLK1), .Q(w951), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g1084 (.C(w32), .A(w948), .B(w591), .Z(w949) );
	vdp_and g1085 (.A(DB[7]), .B(w968), .Z(w930) );
	vdp_and g1086 (.A(w939), .B(w983), .Z(w891) );
	vdp_and g1087 (.A(w951), .B(w950), .Z(w572) );
	vdp_and g1088 (.A(w589), .B(w951), .Z(w593) );
	vdp_and g1089 (.A(w952), .B(w950), .Z(w962) );
	vdp_and g1090 (.A(w589), .B(w952), .Z(w33) );
	vdp_or g1091 (.A(w952), .B(w974), .Z(w958) );
	vdp_or g1092 (.A(w952), .B(w572), .Z(w423) );
	vdp_or g1093 (.A(w589), .B(w452), .Z(w982) );
	vdp_aoi21 g1094 (.A1(w963), .B(SYSRES), .Z(w1491), .A2(w964) );
	vdp_or3 g1095 (.C(w935), .A(w957), .B(w924), .Z(w937) );
	vdp_or3 g1096 (.C(w593), .A(w962), .B(w587), .Z(w584) );
	vdp_or5 g1097 (.C(w946), .A(w934), .B(w584), .Z(w917), .D(w933), .E(w927) );
	vdp_nand3 g1098 (.C(w923), .A(w961), .B(w972), .Z(w823) );
	vdp_2a3oi g1099 (.A1(w922), .B(w979), .Z(w973), .A2(w972), .C(w921) );
	vdp_nand g1100 (.A(w497), .B(w938), .Z(w953) );
	vdp_nor g1101 (.A(w940), .B(w978), .Z(w923) );
	vdp_and4 g1102 (.C(w936), .A(w591), .B(w32), .Z(w959), .D(w960) );
	vdp_nor5 g1103 (.C(w513), .A(w987), .B(w973), .Z(w935), .D(w497), .E(w956) );
	vdp_and g1104 (.A(w589), .B(w987), .Z(w957) );
	vdp_not g1105 (.A(w577), .nZ(w1543) );
	vdp_not g1106 (.A(w1543), .nZ(w1021) );
	vdp_not g1107 (.A(w1002), .nZ(w1037) );
	vdp_not g1108 (.A(w978), .nZ(w1496) );
	vdp_not g1109 (.A(w983), .nZ(w1022) );
	vdp_not g1110 (.A(w1025), .nZ(w933) );
	vdp_not g1111 (.A(w406), .nZ(w954) );
	vdp_not g1112 (.A(w1011), .nZ(w1019) );
	vdp_not g1113 (.A(M5), .nZ(w922) );
	vdp_rs_FF g1114 (.Q(w972), .R(w970), .S(w933) );
	vdp_rs_FF g1115 (.Q(w921), .R(w970), .S(w1045) );
	vdp_rs_FF g1116 (.Q(w979), .R(w970), .S(w968) );
	vdp_rs_FF g1117 (.nQ(w981), .R(w980), .S(w947) );
	vdp_rs_FF g1118 (.Q(w1042), .R(w967), .S(w975) );
	vdp_rs_FF g1119 (.Q(w567), .R(w967), .S(w1035) );
	vdp_rs_FF g1120 (.Q(w566), .R(w967), .S(w993) );
	vdp_or g1121 (.A(w993), .B(w1035), .Z(w1044) );
	vdp_and g1122 (.A(w1042), .B(w920), .Z(w574) );
	vdp_and g1123 (.A(w1041), .B(w1042), .Z(w577) );
	vdp_and g1124 (.A(w1022), .B(w1496), .Z(w920) );
	vdp_and g1125 (.A(w1022), .B(w976), .Z(w1041) );
	vdp_and g1126 (.A(w978), .B(w976), .Z(w1009) );
	vdp_and g1127 (.A(w952), .B(w982), .Z(w984) );
	vdp_and g1128 (.A(w1005), .B(w994), .Z(w414) );
	vdp_and g1129 (.A(w954), .B(w885), .Z(w1051) );
	vdp_and g1130 (.A(w1028), .B(w1027), .Z(w975) );
	vdp_or g1131 (.A(w951), .B(w974), .Z(w985) );
	vdp_or g1132 (.A(w427), .B(w1024), .Z(w966) );
	vdp_or g1133 (.A(SYSRES), .B(w920), .Z(w980) );
	vdp_or g1134 (.A(SYSRES), .B(w983), .Z(w1048) );
	vdp_or g1135 (.A(w978), .B(w977), .Z(w1043) );
	vdp_or g1136 (.A(w1005), .B(w1028), .Z(w1049) );
	vdp_or g1137 (.A(w971), .B(SYSRES), .Z(w1015) );
	vdp_or g1138 (.A(SYSRES), .B(w1010), .Z(w1053) );
	vdp_or g1139 (.A(SYSRES), .B(w1009), .Z(w970) );
	vdp_and g1140 (.A(w969), .B(w943), .Z(w131) );
	vdp_and g1141 (.A(w943), .B(w944), .Z(w108) );
	vdp_and g1142 (.A(w920), .B(w1017), .Z(w1052) );
	vdp_nand g1143 (.A(w414), .B(w981), .Z(w1033) );
	vdp_nor g1144 (.A(w1038), .B(w1021), .Z(w1034) );
	vdp_or5 g1145 (.C(w933), .A(w1020), .B(w1032), .Z(w1031), .D(w885), .E(w1036) );
	vdp_or3 g1146 (.C(w1023), .A(w1005), .B(w409), .Z(w1024) );
	vdp_nor g1147 (.A(w109), .B(w943), .Z(w942) );
	vdp_and3 g1148 (.C(w1054), .A(w1050), .B(w1007), .Z(w1026) );
	vdp_or4 g1149 (.C(w975), .A(w968), .B(w1004), .Z(w971), .D(w414) );
	vdp_and4 g1150 (.C(w1050), .A(w1028), .B(w1012), .Z(w885), .D(w1029) );
	vdp_aoi21 g1151 (.A1(w920), .B(SYSRES), .Z(w1011), .A2(w1018) );
	vdp_aoi21 g1152 (.A1(w885), .B(w1026), .Z(w1025), .A2(w406) );
	vdp_or5 g1153 (.C(w414), .A(w1004), .B(w968), .Z(w1010), .D(w975), .E(w933) );
	vdp_and5 g1154 (.C(w1016), .A(M5), .B(w1050), .Z(w968), .D(w1029), .E(w1028) );
	vdp_not g1155 (.A(CA[7]), .nZ(w998) );
	vdp_not g1156 (.A(w1028), .nZ(w1006) );
	vdp_not g1157 (.A(w1006), .nZ(w991) );
	vdp_not g1158 (.A(w1005), .nZ(w990) );
	vdp_not g1159 (.A(w990), .nZ(w989) );
	vdp_slatch g1160 (.Q(w1030), .D(w992), .nC(w989), .C(w990) );
	vdp_slatch g1161 (.Q(w1050), .D(w992), .nC(w991), .C(w1006), .nQ(w1027) );
	vdp_rs_FF g1162 (.Q(w1013), .R(w1009), .S(w1015) );
	vdp_rs_FF g1163 (.Q(w1017), .R(w1053), .S(w1051), .nQ(w1018) );
	vdp_rs_FF g1164 (.Q(w1054), .R(w1019), .S(w1052), .nQ(w1029) );
	vdp_rs_FF g1165 (.Q(w1016), .R(w1014), .S(w1487), .nQ(w1012) );
	vdp_slatch_r g1166 (.Q(w987), .D(DB[6]), .C(w1008), .nC(w988), .R(w895) );
	vdp_slatch_r g1167 (.Q(w471), .D(DB[5]), .R(w895), .C(w1008), .nC(w988) );
	vdp_slatch_r g1168 (.Q(w470), .D(DB[4]), .R(w895), .C(w1008), .nC(w988) );
	vdp_comp_str g1169 (.A(w968), .Z(w1008), .nZ(w988) );
	vdp_not g1170 (.A(w1488), .nZ(w1014) );
	vdp_aoi21 g1171 (.A1(w920), .B(SYSRES), .Z(w1488), .A2(w1013) );
	vdp_and4 g1172 (.C(w953), .A(M5), .B(w972), .Z(w1487), .D(w920) );
	vdp_and g1173 (.A(w1005), .B(w1030), .Z(w1045) );
	vdp_rs_FF g1174 (.nQ(w1047), .R(w1046), .S(w1045) );
	vdp_rs_FF g1175 (.Q(w977), .R(w1048), .S(w1049) );
	vdp_not g1176 (.A(w992), .nZ(w1594) );
	vdp_not g1177 (.A(CA[2]), .nZ(w1078) );
	vdp_not g1178 (.A(CA[3]), .nZ(w1079) );
	vdp_aon22 g1179 (.Z(w992), .A1(CA[0]), .A2(w1106), .B1(w406), .B2(w1081) );
	vdp_and4 g1180 (.C(w997), .A(w998), .B(CA[6]), .Z(w1040), .D(w996) );
	vdp_and4 g1181 (.C(w1001), .A(w1000), .B(CA[7]), .Z(w1007), .D(w996) );
	vdp_and4 g1182 (.C(CA[3]), .A(w1037), .B(w1039), .Z(w1023), .D(CA[9]) );
	vdp_and4 g1183 (.C(CA[2]), .A(w1037), .B(w1039), .Z(w405), .D(w1079) );
	vdp_and4 g1184 (.C(w1002), .A(w1078), .B(CA[3]), .Z(w999), .D(w1039) );
	vdp_or g1185 (.A(w1040), .B(w405), .Z(w409) );
	vdp_and g1186 (.A(w975), .B(w1034), .Z(w1032) );
	vdp_and g1187 (.A(w1024), .B(w1033), .Z(w1036) );
	vdp_and g1188 (.A(w406), .B(w1031), .Z(w1069) );
	vdp_or g1189 (.A(SYSRES), .B(w947), .Z(w1046) );
	vdp_or g1190 (.A(w1007), .B(w995), .Z(w1028) );
	vdp_or g1191 (.A(SYSRES), .B(w594), .Z(w974) );
	vdp_and3 g1192 (.C(w1077), .A(w968), .B(w1047), .Z(w1020) );
	vdp_and3 g1193 (.C(w1080), .A(w1043), .B(w1212), .Z(w1039) );
	vdp_and5 g1194 (.C(CA[2]), .A(w1002), .B(CA[3]), .Z(w1074), .D(w1594), .E(w1039) );
	vdp_and5 g1195 (.C(CA[2]), .A(w1002), .B(w992), .Z(w1073), .D(CA[3]), .E(w1039) );
	vdp_and5 g1196 (.C(w1078), .A(w1044), .B(w1037), .Z(w1003), .D(w1079), .E(w1039) );
	vdp_and5 g1197 (.C(w1079), .A(w1078), .B(w1044), .Z(w995), .D(w1002), .E(w1039) );
	vdp_nor5 g1198 (.C(w1070), .A(w1073), .B(w1074), .Z(w1056), .D(w999), .E(w1069) );
	vdp_aon22 g1199 (.Z(w1067), .A1(w4), .A2(w1076), .B1(w27), .B2(w406) );
	vdp_aon22 g1200 (.Z(w176), .A1(LS0), .A2(VPOS[8]), .B1(w1064), .B2(VPOS[0]) );
	vdp_not g1201 (.A(LS0), .nZ(w1064) );
	vdp_not g1202 (.A(w406), .nZ(w1060) );
	vdp_not g1203 (.A(w406), .nZ(w1076) );
	vdp_not g1204 (.A(w1540), .nZ(w114) );
	vdp_not g1205 (.A(CA[6]), .nZ(w1000) );
	vdp_not g1206 (.A(w1485), .nZ(w1065) );
	vdp_not g1207 (.A(w992), .nZ(w994) );
	vdp_aoi21 g1208 (.A1(w993), .B(w1486), .Z(w1485), .A2(w999) );
	vdp_and4 g1209 (.C(w997), .A(w1000), .B(CA[7]), .Z(w1484), .D(w996) );
	vdp_and4 g1210 (.C(w1001), .A(w998), .B(CA[6]), .Z(w1486), .D(w996) );
	vdp_slatch g1211 (.Q(w116), .D(w997), .C(w1595), .nC(w1541) );
	vdp_comp_we g1212 (.A(w1058), .Z(w1595), .nZ(w1541) );
	vdp_and g1213 (.A(w47), .B(w1071), .Z(w1542) );
	vdp_and g1214 (.A(w992), .B(w1005), .Z(w1004) );
	vdp_or g1215 (.A(w1003), .B(w1484), .Z(w1005) );
	vdp_or g1216 (.A(w1070), .B(w1542), .Z(w1072) );
	vdp_or g1217 (.Z(w1066), .A(w7), .B(SYSRES) );
	vdp_and g1218 (.Z(w112), .A(w58), .B(w1067) );
	vdp_rs_FF g1219 (.Q(w1062), .R(w1066), .S(w112) );
	vdp_aoi221 g1220 (.Z(w1540), .A1(w113), .A2(1'b0), .B1(w1068), .B2(w1072), .C(w115) );
	vdp_aoi22 g1221 (.Z(w1057), .A1(w1063), .A2(w1060), .B1(w406), .B2(w1062) );
	vdp_comp_str g1222 (.Z(w1094), .A(w58), .nZ(w1095) );
	vdp_comp_str g1223 (.Z(w1120), .A(CA[14]), .nZ(w1121) );
	vdp_comp_str g1224 (.Z(w1130), .A(w1138), .nZ(w1131) );
	vdp_comp_str g1225 (.Z(w1127), .A(w1137), .nZ(w1126) );
	vdp_not g1226 (.A(w1136), .nZ(w1139) );
	vdp_not g1227 (.A(w1128), .nZ(w1141) );
	vdp_not g1228 (.A(w1125), .nZ(w1140) );
	vdp_not g1229 (.A(w1140), .nZ(w1105) );
	vdp_not g1230 (.A(w406), .nZ(w1106) );
	vdp_not g1231 (.A(w1141), .nZ(w1124) );
	vdp_not g1232 (.A(w1143), .nZ(w1123) );
	vdp_not g1233 (.A(w1142), .nZ(w1122) );
	vdp_aon222 g1234 (.C2(w1122), .B2(w1123), .A2(w1124), .C1(w1103), .B1(CA[15]), .A1(CA[7]), .Z(w1115) );
	vdp_aon222 g1235 (.C2(w1122), .B2(w1123), .A2(w1124), .C1(w1102), .B1(CA[13]), .A1(CA[6]), .Z(w1114) );
	vdp_aon222 g1236 (.C2(w1122), .B2(w1123), .A2(w1124), .C1(w1101), .B1(CA[12]), .A1(CA[5]), .Z(w1113) );
	vdp_aon222 g1237 (.C2(w1122), .B2(w1123), .A2(w1124), .C1(w1100), .B1(CA[11]), .A1(CA[4]), .Z(w1112) );
	vdp_aon222 g1238 (.C2(w1122), .B2(w1123), .A2(w1124), .C1(w1104), .B1(CA[10]), .A1(CA[3]), .Z(w1111) );
	vdp_aon222 g1239 (.C2(w1122), .B2(w1123), .A2(w1124), .C1(w1524), .B1(CA[9]), .A1(CA[2]), .Z(w1110) );
	vdp_aon222 g1240 (.C2(w1122), .B2(w1123), .A2(w1124), .C1(w1107), .B1(CA[8]), .A1(w1081), .Z(w1109) );
	vdp_aon222 g1241 (.C2(w1122), .B2(w1123), .A2(w1124), .C1(w1097), .B1(CA[14]), .A1(CA[0]), .Z(w1108) );
	vdp_aon222 g1242 (.C2(w1122), .B2(w1123), .A2(w1124), .C1(nHCLK1), .B1(1'b1), .A1(1'b0), .Z(w1125) );
	vdp_slatch g1243 (.Q(LS0), .D(w1117), .C(w1094), .nC(w1095) );
	vdp_slatch g1244 (.Q(w1093), .D(w1129), .C(w1094), .nC(w1095) );
	vdp_aon22 g1245 (.Z(w1096), .A1(COL[6]), .A2(w1132), .B1(w129), .B2(w1494) );
	vdp_not g1246 (.A(w1119), .nZ(w1091) );
	vdp_not g1247 (.A(w1132), .nZ(w1494) );
	vdp_and g1248 (.Z(w1), .A(w1093), .B(LS0) );
	vdp_and g1249 (.Z(w1092), .A(M5), .B(w1091) );
	vdp_and g1250 (.Z(w1495), .A(M5), .B(w1119) );
	vdp_and g1251 (.Z(128k), .A(M5), .B(w1118) );
	vdp_or3 g1252 (.Z(w1136), .A(w1133), .B(w1134), .C(w1401) );
	vdp_and g1253 (.Z(w1135), .A(w1133), .B(w1105) );
	vdp_nand g1254 (.Z(w1143), .A(w1141), .B(w1136) );
	vdp_nand g1255 (.Z(w1142), .A(w1141), .B(w1139) );
	vdp_slatch g1256 (.Q(w91), .D(REG_BUS[0]), .C(w1120), .nC(w1121) );
	vdp_slatch g1257 (.Q(w93), .D(REG_BUS[1]), .C(w1120), .nC(w1121) );
	vdp_slatch g1258 (.Q(w44), .D(REG_BUS[2]), .C(w1120), .nC(w1121) );
	vdp_slatch g1259 (.Q(w1144), .D(REG_BUS[3]), .C(w1120), .nC(w1121) );
	vdp_slatch g1260 (.Q(w111), .D(REG_BUS[4]), .C(w1120), .nC(w1121) );
	vdp_slatch g1261 (.Q(w94), .D(REG_BUS[5]), .C(w1120), .nC(w1121) );
	vdp_slatch g1262 (.Q(w1071), .D(REG_BUS[6]), .C(w1120), .nC(w1121) );
	vdp_slatch g1263 (.Q(w1128), .D(REG_BUS[7]), .C(w1120), .nC(w1121) );
	vdp_slatch g1264 (.Q(w1119), .D(REG_BUS[3]), .C(w1127), .nC(w1126) );
	vdp_slatch g1265 (.Q(w1118), .D(REG_BUS[7]), .C(w1127), .nC(w1126) );
	vdp_slatch g1266 (.Q(w19), .D(REG_BUS[4]), .C(w1130), .nC(w1131) );
	vdp_slatch g1267 (.Q(w89), .D(REG_BUS[3]), .C(w1130), .nC(w1131) );
	vdp_slatch g1268 (.Q(w1129), .D(REG_BUS[2]), .C(w1130), .nC(w1131) );
	vdp_slatch g1269 (.Q(w1117), .D(REG_BUS[1]), .C(w1130), .nC(w1131) );
	vdp_slatch g1270 (.Q(H40), .D(REG_BUS[0]), .C(w1130), .nC(w1131) );
	vdp_slatch g1271 (.Q(w45), .D(REG_BUS[0]), .C(w1127), .nC(w1126) );
	vdp_slatch g1272 (.Q(w132), .D(REG_BUS[1]), .C(w1127), .nC(w1126) );
	vdp_slatch g1273 (.Q(M5), .D(REG_BUS[2]), .C(w1127), .nC(w1126) );
	vdp_slatch g1274 (.Q(w1146), .D(REG_BUS[4]), .C(w1127), .nC(w1126) );
	vdp_slatch g1275 (.Q(w1145), .D(REG_BUS[5]), .C(w1127), .nC(w1126) );
	vdp_slatch g1276 (.Q(w1116), .D(REG_BUS[6]), .C(w1127), .nC(w1126) );
	vdp_and g1277 (.Z(w119), .A(w1073), .B(w1155) );
	vdp_and g1278 (.Z(w123), .A(w1023), .B(w1155) );
	vdp_and g1279 (.Z(w118), .A(w1073), .B(w1156) );
	vdp_and g1280 (.Z(w122), .A(w1023), .B(w1156) );
	vdp_and g1281 (.Z(w120), .A(w1073), .B(w1150) );
	vdp_and g1282 (.Z(w121), .A(w1023), .B(w1150) );
	vdp_and g1283 (.Z(w57), .A(w1073), .B(w1151) );
	vdp_and g1284 (.Z(w48), .A(w1023), .B(w1151) );
	vdp_and g1285 (.Z(w90), .A(w1073), .B(w1153) );
	vdp_and g1286 (.Z(w88), .A(w1023), .B(w1153) );
	vdp_and g1287 (.Z(w92), .A(w1073), .B(w1154) );
	vdp_and g1288 (.Z(PSG_TEST_OE), .A(w1023), .B(w1154) );
	vdp_and g1289 (.Z(w1172), .A(w1073), .B(w1158) );
	vdp_and g1290 (.Z(w1147), .A(w1073), .B(w1159) );
	vdp_and g1291 (.Z(w56), .A(w1073), .B(w1152) );
	vdp_and g1292 (.Z(w54), .A(w1023), .B(w1152) );
	vdp_dslatch g1293 (.D(COL[0]), .C(HCLK1), .Q(w1097), .nC(nHCLK1) );
	vdp_dslatch g1294 (.D(COL[1]), .Q(w1107), .C(HCLK1), .nC(nHCLK1) );
	vdp_dslatch g1295 (.D(COL[2]), .Q(w1524), .C(HCLK1), .nC(nHCLK1) );
	vdp_dslatch g1296 (.D(COL[3]), .Q(w1104), .C(HCLK1), .nC(nHCLK1) );
	vdp_dslatch g1297 (.D(COL[4]), .Q(w1100), .C(HCLK1), .nC(nHCLK1) );
	vdp_dslatch g1298 (.D(COL[5]), .Q(w1101), .C(HCLK1), .nC(nHCLK1) );
	vdp_dslatch g1299 (.D(w1096), .Q(w1102), .C(HCLK1), .nC(nHCLK1) );
	vdp_dslatch g1300 (.D(w130), .Q(w1103), .C(HCLK1), .nC(nHCLK1) );
	vdp_slatch g1301 (.Q(w52), .D(REG_BUS[5]), .C(w1131), .nC(w1130) );
	vdp_slatch g1302 (.Q(w39), .D(REG_BUS[6]), .C(w1131), .nC(w1130) );
	vdp_slatch g1303 (.Q(w1148), .D(REG_BUS[7]), .C(w1131), .nC(w1130) );
	vdp_slatch g1304 (.Q(w23), .D(REG_BUS[3]), .nC(w1180), .C(w1178) );
	vdp_slatch g1305 (.Q(w97), .D(REG_BUS[2]), .nC(w1180), .C(w1178) );
	vdp_slatch g1306 (.Q(w476), .D(REG_BUS[1]), .nC(w1180), .C(w1178) );
	vdp_slatch g1307 (.Q(w53), .D(REG_BUS[0]), .nC(w1180), .C(w1178) );
	vdp_slatch g1308 (.Q(w95), .D(REG_BUS[7]), .nC(w1180), .C(w1178) );
	vdp_slatch g1309 (.Q(w96), .D(REG_BUS[6]), .nC(w1180), .C(w1178) );
	vdp_slatch g1310 (.Q(w59), .D(REG_BUS[5]), .nC(w1180), .C(w1178) );
	vdp_slatch g1311 (.Q(w1177), .D(REG_BUS[4]), .nC(w1180), .C(w1178) );
	vdp_slatch_r g1312 (.Q(w124), .D(DB[14]), .nC(w1171), .R(w1167), .C(w1175) );
	vdp_slatch_r g1313 (.Q(w128), .D(DB[13]), .R(w1167), .nC(w1171), .C(w1175) );
	vdp_slatch_r g1314 (.Q(w125), .D(DB[12]), .R(w1167), .nC(w1171), .C(w1175) );
	vdp_comp_str g1315 (.Z(w1178), .A(w1176), .nZ(w1180) );
	vdp_comp_str g1316 (.Z(w1174), .A(w1147), .nZ(w1173) );
	vdp_not g1317 (.A(REG_BUS[6]), .nZ(w1492) );
	vdp_not g1318 (.A(REG_BUS[7]), .nZ(w1195) );
	vdp_not g1319 (.A(REG_BUS[4]), .nZ(w1181) );
	vdp_not g1320 (.A(REG_BUS[5]), .nZ(w1179) );
	vdp_not g1321 (.A(REG_BUS[2]), .nZ(w1196) );
	vdp_not g1322 (.A(REG_BUS[3]), .nZ(w1182) );
	vdp_not g1323 (.A(REG_BUS[0]), .nZ(w1190) );
	vdp_not g1324 (.A(REG_BUS[1]), .nZ(w1191) );
	vdp_not g1325 (.A(w1165), .nZ(w1184) );
	vdp_not g1326 (.A(w1166), .nZ(w1169) );
	vdp_not g1327 (.A(w1157), .nZ(w1183) );
	vdp_not g1328 (.A(w1170), .nZ(w1185) );
	vdp_comp_str g1329 (.Z(DB[9]), .nZ(w1168), .A(w1074) );
	vdp_slatch_r g1330 (.Q(w1170), .R(w1167), .D(DB[11]), .nC(w1168), .C(DB[9]) );
	vdp_slatch_r g1331 (.Q(w1157), .D(DB[10]), .nC(w1168), .R(w1167), .C(DB[9]) );
	vdp_and4 g1332 (.Z(w1501), .A(w1165), .B(w1166), .C(w1170), .D(w1157) );
	vdp_and4 g1333 (.Z(w1150), .A(w1170), .B(w1183), .C(w1169), .D(w1184) );
	vdp_and4 g1334 (.Z(w1156), .A(w1185), .B(w1157), .C(w1166), .D(w1165) );
	vdp_and4 g1335 (.Z(w1155), .A(w1185), .B(w1157), .C(w1166), .D(w1184) );
	vdp_and4 g1336 (.Z(w1154), .A(w1185), .B(w1157), .C(w1169), .D(w1165) );
	vdp_and4 g1337 (.Z(w1153), .A(w1185), .B(w1157), .C(w1169), .D(w1184) );
	vdp_and4 g1338 (.Z(w1151), .A(w1185), .B(w1183), .C(w1166), .D(w1165) );
	vdp_and4 g1339 (.Z(w1152), .A(w1185), .B(w1183), .C(w1166), .D(w1184) );
	vdp_and4 g1340 (.Z(w1159), .A(w1185), .B(w1183), .C(w1169), .D(w1165) );
	vdp_and4 g1341 (.Z(w1158), .A(w1185), .B(w1183), .C(w1169), .D(w1184) );
	vdp_nand g1342 (.Z(w1438), .A(w1501), .B(w1073) );
	vdp_slatch_r g1343 (.Q(w1165), .D(DB[8]), .R(w1167), .C(DB[9]), .nC(w1168) );
	vdp_slatch_r g1344 (.Q(w1164), .D(DB[11]), .R(w1167), .C(w1175), .nC(w1171) );
	vdp_slatch_r g1345 (.nC(w1187), .Q(w1166), .D(DB[9]), .R(w1167), .C(w1168) );
	vdp_slatch_r g1346 (.Q(w1163), .D(DB[10]), .R(w1167), .C(w1175), .nC(w1171) );
	vdp_slatch_r g1347 (.Q(w99), .D(DB[8]), .R(w1167), .C(w1175), .nC(w1171) );
	vdp_slatch_r g1348 (.Q(w1162), .D(DB[9]), .R(w1167), .C(w1175), .nC(w1171) );
	vdp_slatch_r g1349 (.Q(w98), .D(DB[7]), .R(w1167), .C(w1175), .nC(w1171) );
	vdp_slatch_r g1350 (.Q(w100), .D(DB[5]), .R(w1167), .C(w1175), .nC(w1171) );
	vdp_slatch_r g1351 (.Q(w101), .D(DB[6]), .R(w1167), .C(w1175), .nC(w1171) );
	vdp_slatch_r g1352 (.Q(w969), .D(DB[4]), .R(w1167), .C(w1175), .nC(w1171) );
	vdp_slatch_r g1353 (.Q(w1193), .D(DB[2]), .R(w1167), .C(w1175), .nC(w1171) );
	vdp_slatch_r g1354 (.Q(w1194), .D(DB[3]), .R(w1167), .C(w1175), .nC(w1171) );
	vdp_slatch_r g1355 (.Q(w1132), .D(DB[0]), .R(w1167), .C(w1175), .nC(w1171) );
	vdp_slatch_r g1356 (.Q(w795), .D(DB[1]), .R(w1167), .C(w1175), .nC(w1171) );
	vdp_slatch_r g1357 (.Q(w105), .D(DB[9]), .R(w1167), .C(w1174), .nC(w1173) );
	vdp_slatch_r g1358 (.Q(w106), .D(DB[10]), .R(w1167), .C(w1174), .nC(w1173) );
	vdp_slatch_r g1359 (.Q(w103), .D(DB[7]), .R(w1167), .C(w1174), .nC(w1173) );
	vdp_slatch_r g1360 (.Q(w104), .D(DB[8]), .R(w1167), .C(w1174), .nC(w1173) );
	vdp_slatch_r g1361 (.Q(w51), .D(DB[5]), .R(w1167), .C(w1174), .nC(w1173) );
	vdp_slatch_r g1362 (.Q(w41), .D(DB[6]), .R(w1167), .C(w1174), .nC(w1173) );
	vdp_slatch_r g1363 (.Q(w40), .D(DB[3]), .R(w1167), .C(w1174), .nC(w1173) );
	vdp_slatch_r g1364 (.Q(w42), .D(DB[4]), .R(w1167), .C(w1174), .nC(w1173) );
	vdp_slatch_r g1365 (.Q(w1493), .D(DB[1]), .R(w1167), .C(w1174), .nC(w1173) );
	vdp_slatch_r g1366 (.Q(w55), .D(DB[2]), .R(w1167), .C(w1174), .nC(w1173) );
	vdp_slatch_r g1367 (.Q(w43), .D(DB[0]), .R(w1167), .C(w1174), .nC(w1173) );
	vdp_comp_str g1368 (.Z(w1175), .nZ(w1171), .A(w1172) );
	vdp_notif0 g1369 (.A(VPOS[9]), .nZ(DB[10]), .nE(w1188) );
	vdp_notif0 g1370 (.A(VPOS[8]), .nZ(DB[9]), .nE(w1188) );
	vdp_bufif0 g1371 (.A(w591), .Z(DB[9]), .nE(w1220) );
	vdp_bufif0 g1372 (.A(w1038), .Z(DB[8]), .nE(w1220) );
	vdp_bufif0 g1373 (.A(w1219), .Z(DB[1]), .nE(w1220) );
	vdp_bufif0 g1374 (.A(w1221), .Z(DB[0]), .nE(w1220) );
	vdp_bufif0 g1375 (.A(w1201), .Z(DB[7]), .nE(w1220) );
	vdp_bufif0 g1376 (.A(w1200), .Z(DB[6]), .nE(w1220) );
	vdp_bufif0 g1377 (.A(w1199), .Z(DB[5]), .nE(w1220) );
	vdp_bufif0 g1378 (.A(ODD/EVEN), .Z(DB[4]), .nE(w1220) );
	vdp_bufif0 g1379 (.A(w46), .Z(DB[3]), .nE(w1220) );
	vdp_bufif0 g1380 (.A(w21), .Z(DB[2]), .nE(w1220) );
	vdp_slatch_r g1381 (.Q(w80), .D(DB[4]), .R(w1167), .C(w1168), .nC(w1187) );
	vdp_slatch_r g1382 (.Q(w81), .D(DB[5]), .R(w1167), .C(w1168), .nC(w1187) );
	vdp_slatch_r g1383 (.Q(w83), .D(DB[7]), .R(w1167), .C(w1168), .nC(w1187) );
	vdp_slatch_r g1384 (.Q(w82), .D(DB[6]), .R(w1167), .C(w1168), .nC(w1187) );
	vdp_slatch_r g1385 (.Q(w76), .D(DB[0]), .R(w1167), .C(w1168), .nC(w1187) );
	vdp_slatch_r g1386 (.Q(w77), .D(DB[1]), .R(w1167), .C(w1168), .nC(w1187) );
	vdp_slatch_r g1387 (.Q(w79), .D(DB[3]), .R(w1167), .C(w1168), .nC(w1187) );
	vdp_slatch_r g1388 (.Q(w78), .D(DB[2]), .R(w1167), .C(w1168), .nC(w1187) );
	vdp_notif0 g1389 (.A(HPOS[0]), .nZ(DB[8]), .nE(w1188) );
	vdp_not g1390 (.A(w406), .nZ(w1502) );
	vdp_comp_str g1391 (.Z(w1189), .A(w803), .nZ(w1192) );
	vdp_slatch_r g1392 (.Q(w1205), .D(w1190), .R(w1208), .C(w1189), .nC(w1192) );
	vdp_slatch_r g1393 (.Q(w1216), .D(w1196), .R(w1208), .C(w1189), .nC(w1192) );
	vdp_slatch_r g1394 (.Q(w1222), .D(w1191), .R(w1208), .C(w1189), .nC(w1192) );
	vdp_slatch_r g1395 (.Q(w1210), .D(w1492), .R(w1208), .C(w1189), .nC(w1192) );
	vdp_slatch_r g1396 (.Q(w1217), .D(w1182), .R(w1208), .C(w1189), .nC(w1192) );
	vdp_slatch_r g1397 (.Q(w1209), .D(w1179), .R(w1208), .C(w1189), .nC(w1192) );
	vdp_slatch_r g1398 (.Q(w1218), .D(w1181), .R(w1208), .C(w1189), .nC(w1192) );
	vdp_slatch_r g1399 (.Q(w1211), .D(w1195), .R(w1208), .C(w1189), .nC(w1192) );
	vdp_aon22 g1400 (.Z(w1219), .A1(w591), .A2(w1203), .B1(w1204), .B2(DMA_BUSY) );
	vdp_aon22 g1401 (.Z(w1221), .A1(w1038), .A2(w1203), .B1(w1204), .B2(PAL) );
	vdp_and3 g1402 (.C(w1193), .A(w409), .B(w1502), .Z(w1198) );
	vdp_not g1403 (.A(w1198), .nZ(w1188) );
	vdp_not g1404 (.A(w1004), .nZ(w1220) );
	vdp_cnt_bit_load g1405 (.V(w1211), .nL(w1227), .L(w1206), .R(1'b0), .Q(w1228), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1256) );
	vdp_cnt_bit_load g1406 (.V(w1210), .nL(w1227), .L(w1206), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1534), .CO(w1256) );
	vdp_cnt_bit_load g1407 (.V(w1209), .nL(w1227), .L(w1206), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1255), .CO(w1534) );
	vdp_cnt_bit_load g1408 (.V(w1218), .nL(w1227), .L(w1206), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1254), .CO(w1255) );
	vdp_cnt_bit_load g1409 (.V(w1217), .nL(w1227), .L(w1206), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1253), .CO(w1254) );
	vdp_cnt_bit_load g1410 (.V(w1216), .nL(w1227), .L(w1206), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1544), .CO(w1253) );
	vdp_cnt_bit_load g1411 (.V(w1222), .nL(w1227), .L(w1206), .R(1'b0), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2), .CI(w1252), .CO(w1544) );
	vdp_cnt_bit_load g1412 (.V(w1205), .nL(w1227), .L(w1206), .R(1'b0), .CI(w1224), .CO(w1252), .C1(HCLK1), .C2(HCLK2), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g1413 (.D(w1498), .C2(HCLK2), .C1(HCLK1), .Q(w1229), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_rs_FF g1414 (.Q(w1200), .R(w1245), .S(w1246) );
	vdp_rs_FF g1415 (.Q(w1201), .R(w1244), .S(w112) );
	vdp_rs_FF g1416 (.Q(w1199), .R(w1245), .S(w126) );
	vdp_not g1417 (.A(M5), .nZ(w1243) );
	vdp_not g1418 (.A(w1201), .nZ(w1223) );
	vdp_not g1419 (.A(w1207), .nZ(w1213) );
	vdp_not g1420 (.A(CA[21]), .nZ(w1499) );
	vdp_not g1421 (.A(w406), .nZ(w1214) );
	vdp_not g1422 (.A(w1248), .nZ(w1215) );
	vdp_comp_we g1423 (.Z(w1227), .A(w1497), .nZ(w1206) );
	vdp_or g1424 (.A(w1248), .B(w1229), .Z(w1497) );
	vdp_and g1425 (.A(w1215), .B(w1228), .Z(w1498) );
	vdp_and g1426 (.A(w1223), .B(w127), .Z(w1246) );
	vdp_or g1427 (.A(w1194), .B(w4), .Z(w1224) );
	vdp_not g1428 (.A(w1203), .nZ(w1204) );
	vdp_nor3 g1429 (.A(w406), .B(w1243), .Z(w1203), .C(CA[1]) );
	vdp_nor3 g1430 (.A(w1194), .B(w5), .Z(w1248), .C(w31) );
	vdp_nor g1431 (.A(w1251), .B(w1230), .Z(w1212) );
	vdp_or5 g1432 (.A(w1214), .B(CA[4]), .C(CA[5]), .D(CA[15]), .Z(w1251), .E(CA[6]) );
	vdp_or5 g1433 (.A(CA[16]), .B(CA[17]), .C(CA[20]), .D(w1213), .Z(w1230), .E(w1499) );
	vdp_rs_FF g1434 (.Q(w1236), .R(w1289), .S(w1498) );
	vdp_rs_FF g1435 (.Q(w1290), .R(w1273), .S(w1500) );
	vdp_dff g1436 (.Q(w1293), .R(w1249), .C(w1239), .D(w1232) );
	vdp_dff g1437 (.Q(w1292), .R(w1249), .C(w1239), .D(w1231) );
	vdp_dff g1438 (.Q(w1294), .R(w1249), .C(w1239), .D(w1233) );
	vdp_rs_FF g1439 (.Q(w1550), .R(w1288), .S(w1549) );
	vdp_rs_FF g1440 (.Q(w1260), .R(w1261), .S(w1547) );
	vdp_dlatch_inv g1441 (.D(w1267), .Q(w1268), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g1442 (.D(w1261), .C(DCLK1), .Q(w1267), .nC(nDCLK1) );
	vdp_dlatch_inv g1443 (.D(w1271), .Q(w1245), .C(HCLK1), .nC(nHCLK1) );
	vdp_not g1444 (.A(w1284), .nZ(w1257) );
	vdp_not g1445 (.A(w671), .nZ(w1235) );
	vdp_not g1446 (.A(w1238), .nZ(w1233) );
	vdp_not g1447 (.A(w1237), .nZ(w1232) );
	vdp_not g1448 (.A(w1247), .nZ(w1249) );
	vdp_not g1449 (.A(w1264), .nZ(w1239) );
	vdp_not g1450 (.A(w1240), .nZ(w50) );
	vdp_not g1451 (.A(w1242), .nZ(w1241) );
	vdp_sr_bit g1452 (.D(w1269), .C2(HCLK2), .C1(HCLK1), .Q(w1288), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and g1453 (.A(M5), .B(w1260), .Z(w1264) );
	vdp_and g1454 (.A(w406), .B(w1259), .Z(w1080) );
	vdp_and g1455 (.A(w1240), .B(w1080), .Z(w1548) );
	vdp_or g1456 (.A(w427), .B(w1548), .Z(w1547) );
	vdp_or g1457 (.A(w1004), .B(SYSRES), .Z(w1549) );
	vdp_and g1458 (.A(w1243), .B(w1245), .Z(w1272) );
	vdp_or g1459 (.A(w1292), .B(w1272), .Z(w1273) );
	vdp_and g1460 (.A(M5), .B(w473), .Z(w1500) );
	vdp_and g1461 (.A(w1146), .B(M5), .Z(w1234) );
	vdp_or g1462 (.A(w1294), .B(w1272), .Z(w1244) );
	vdp_or g1463 (.A(w1293), .B(w1272), .Z(w1289) );
	vdp_comp_DFF g1464 (.D(w1550), .C2(HCLK2), .C1(HCLK1), .Q(w1269), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_comp_DFF g1465 (.D(w1264), .C2(DCLK2), .C1(DCLK1), .Q(w1261), .nC2(nDCLK2), .nC1(nDCLK1) );
	vdp_nor g1466 (.A(w1269), .B(SYSRES), .Z(w1270) );
	vdp_nand g1467 (.A(w1288), .B(w1270), .Z(w1271) );
	vdp_nand g1468 (.A(w1201), .B(w1145), .Z(w1238) );
	vdp_and3 g1469 (.A(w1234), .B(w930), .Z(w1283), .C(w1235) );
	vdp_and3 g1470 (.A(w1234), .B(w930), .Z(w1282), .C(w671) );
	vdp_and4 g1471 (.A(w1237), .B(w1144), .C(w1238), .D(w1290), .Z(w1231) );
	vdp_nand3 g1472 (.C(w1236), .A(w1238), .B(w1177), .Z(w1237) );
	vdp_aoi21 g1473 (.A1(w1268), .B(SYSRES), .Z(w1247), .A2(w1267) );
	vdp_dff g1474 (.Q(w1313), .R(w1299), .C(w1296), .D(w1281) );
	vdp_dff g1475 (.Q(w1309), .R(w1299), .C(w1296), .D(w1308) );
	vdp_dff g1476 (.Q(w1278), .R(w1299), .C(w1296), .D(w1276) );
	vdp_dff g1477 (.Q(w1286), .R(w1299), .C(w1296), .D(w1285) );
	vdp_dff g1478 (.Q(w1287), .R(w1299), .C(w1296), .D(w1275) );
	vdp_dff g1479 (.Q(w1265), .R(w1299), .C(w1296), .D(w1304) );
	vdp_dff g1480 (.Q(w1262), .R(w1299), .C(w1296), .D(w1302) );
	vdp_dff g1481 (.Q(w1295), .R(1'b0), .C(w1296), .D(w1258) );
	vdp_ha g1482 (.SUM(w1302), .A(w1262), .B(w1257), .CO(w1263) );
	vdp_ha g1483 (.SUM(w1304), .A(w1265), .B(w1263), .CO(w1266) );
	vdp_ha g1484 (.SUM(w1275), .A(w1287), .B(w1266), .CO(w1274) );
	vdp_ha g1485 (.SUM(w1285), .A(w1286), .B(w1274), .CO(w1279) );
	vdp_ha g1486 (.SUM(w1276), .A(w1278), .B(w1279), .CO(w1277) );
	vdp_ha g1487 (.SUM(w1281), .A(w1313), .B(w1277), .CO(w1280) );
	vdp_ha g1488 (.SUM(w1308), .A(w1309), .B(w1280) );
	vdp_and3 g1489 (.A(w1309), .B(w1278), .Z(w1306), .C(w1313) );
	vdp_and4 g1490 (.C(w1265), .A(w1286), .B(w1306), .Z(w1312), .D(w1287) );
	vdp_nand g1491 (.A(w1295), .B(w406), .Z(w1436) );
	vdp_dff g1492 (.Q(w1321), .R(1'b0), .C(w1296), .D(w1301) );
	vdp_dff g1493 (.Q(w1301), .R(w1303), .C(w1296), .D(w1326) );
	vdp_dff g1494 (.Q(w1326), .R(w1303), .C(w1324), .D(w1305) );
	vdp_dff g1495 (.Q(w1305), .R(w1303), .C(w1296), .D(w1330) );
	vdp_dff g1496 (.Q(w1330), .R(w1303), .C(w1296), .D(w1331) );
	vdp_dff g1497 (.Q(w1331), .R(w1303), .C(w1296), .D(1'b1) );
	vdp_dff g1498 (.Q(w1537), .R(w1340), .C(w1314), .D(w1306) );
	vdp_dff g1499 (.Q(w1314), .R(1'b0), .C(w1296), .D(w1312) );
	vdp_dff g1500 (.Q(w1333), .R(w1311), .C(w1334), .D(w1306) );
	vdp_dff g1501 (.Q(w1310), .R(w1325), .C(w1338), .D(1'b1) );
	vdp_or g1502 (.A(SYSRES), .B(w1310), .Z(w1311) );
	vdp_or g1503 (.A(w1303), .B(w1321), .Z(w1336) );
	vdp_not g1504 (.A(w1321), .nZ(w1298) );
	vdp_not g1505 (.A(w1537), .nZ(w1303) );
	vdp_nand3 g1506 (.A(w406), .B(w1319), .Z(w1299), .C(w1298) );
	vdp_not g1507 (.nZ(w1324), .A(w1320) );
	vdp_not g1508 (.nZ(w1296), .A(w1297) );
	vdp_dff g1509 (.Q(w1323), .R(1'b0), .C(w1324), .D(w1346) );
	vdp_dff g1510 (.Q(w1349), .R(w1325), .C(w1324), .D(w1329) );
	vdp_dff g1511 (.Q(w1329), .R(w1325), .C(w1296), .D(w1351) );
	vdp_dff g1512 (.Q(w1351), .R(w1325), .C(w1324), .D(w1328) );
	vdp_dff g1513 (.Q(w1328), .R(w1325), .C(w1324), .D(w1339) );
	vdp_dff g1514 (.Q(w1339), .R(w1325), .C(w1296), .D(w47) );
	vdp_dff g1515 (.Q(w1356), .R(w1355), .C(w1324), .D(w1134) );
	vdp_dff g1516 (.Q(w1134), .R(w1355), .C(w1296), .D(w1335) );
	vdp_not g1517 (.A(w1343), .nZ(w113) );
	vdp_not g1518 (.A(w1002), .nZ(w1318) );
	vdp_not g1519 (.A(w1329), .nZ(w1327) );
	vdp_not g1520 (.A(w1326), .nZ(w1545) );
	vdp_not g1521 (.A(w1335), .nZ(w1355) );
	vdp_not g1522 (.A(w1080), .nZ(w1338) );
	vdp_not g1523 (.A(w1240), .nZ(w1538) );
	vdp_and g1524 (.A(w1336), .B(w1080), .Z(w1335) );
	vdp_and g1525 (.A(w1337), .B(w1335), .Z(w1334) );
	vdp_and g1526 (.A(w1356), .B(w1334), .Z(w47) );
	vdp_and g1527 (.A(w1330), .B(w1545), .Z(w1347) );
	vdp_and g1528 (.A(w1331), .B(w1545), .Z(w1348) );
	vdp_and g1529 (.A(w1322), .B(w993), .Z(w1345) );
	vdp_and g1530 (.A(w1322), .B(w1035), .Z(w1317) );
	vdp_and g1531 (.A(w1002), .B(w1323), .Z(w1322) );
	vdp_and g1532 (.A(w113), .B(w1134), .Z(w1068) );
	vdp_nand g1533 (.A(w1328), .B(w1327), .Z(w1319) );
	vdp_nor g1534 (.A(w1325), .B(w1339), .Z(w1350) );
	vdp_or3 g1535 (.C(w1333), .A(SYSRES), .B(w1321), .Z(w1340) );
	vdp_oai21 g1536 (.A1(w1035), .B(w1318), .Z(w1343), .A2(w993) );
	vdp_dff g1537 (.Q(w1364), .R(1'b0), .C(w1296), .D(w1242) );
	vdp_rs_FF g1538 (.nQ(w1077), .R(w1365), .S(w1362) );
	vdp_not g1539 (.A(w1370), .nZ(w1058) );
	vdp_not g1540 (.A(REG_BUS[7]), .nZ(w1361) );
	vdp_and3 g1541 (.C(w1361), .A(w828), .B(M5), .Z(w1362) );
	vdp_or g1542 (.A(w1242), .B(SYSRES), .Z(w1365) );
	vdp_and g1543 (.A(w1382), .B(w592), .Z(w1383) );
	vdp_not g1544 (.A(w1337), .nZ(w1385) );
	vdp_and4 g1545 (.C(CA[21]), .A(w1207), .B(CA[20]), .Z(w1337), .D(w1538) );
	vdp_dff g1546 (.Q(w1425), .R(1'b0), .C(w1370), .D(w1410) );
	vdp_dff g1547 (.Q(w1405), .R(1'b0), .C(w1370), .D(w1404) );
	vdp_dff g1548 (.Q(w1344), .R(1'b0), .C(w1391), .D(w1392) );
	vdp_dff g1549 (.Q(w1404), .R(1'b0), .C(w1391), .D(w1344) );
	vdp_dff g1550 (.Q(w1417), .R(w1418), .C(HCLK2), .D(w1420) );
	vdp_dff g1551 (.Q(DMA_BUSY), .R(w1418), .C(HCLK2), .D(w1417) );
	vdp_rs_FF g1552 (.Q(w1284), .R(w1418), .S(w1353) );
	vdp_rs_FF g1553 (.Q(w1539), .R(w1418), .S(w1282) );
	vdp_rs_FF g1554 (.Q(w1258), .R(w1354), .S(w1283) );
	vdp_sr_bit g1555 (.D(w592), .Q(w1382), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1556 (.D(w1546), .Q(w1416), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_dlatch_inv g1557 (.D(w1381), .nQ(w1359), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g1558 (.D(w1380), .nQ(w1381), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g1559 (.D(w1367), .C(HCLK1), .nQ(w1380), .nC(nHCLK1) );
	vdp_aon22 g1560 (.Z(w1412), .A2(w1358), .B1(w1380), .B2(w1421), .A1(w1359) );
	vdp_sr_bit g1561 (.D(w1422), .Q(w1427), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1562 (.D(w1384), .Q(w1422), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g1563 (.D(VRAM_REFRESH), .C2(HCLK2), .C1(HCLK1), .Q(w1384), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_aon22 g1564 (.Z(w1400), .A2(w1350), .B1(w1428), .B2(w1431), .A1(w1398) );
	vdp_not g1565 (.A(w1536), .nZ(w1070) );
	vdp_not g1566 (.A(w1350), .nZ(w1431) );
	vdp_not g1567 (.A(w1416), .nZ(w1421) );
	vdp_not g1568 (.A(w1357), .nZ(w1399) );
	vdp_not g1569 (.A(w1333), .nZ(w1325) );
	vdp_or g1570 (.A(w1284), .B(w1539), .Z(w1420) );
	vdp_or g1571 (.A(SYSRES), .B(w594), .Z(w1418) );
	vdp_or g1572 (.A(w1353), .B(w1418), .Z(w1354) );
	vdp_or g1573 (.A(w1233), .B(w1231), .Z(w279) );
	vdp_or g1574 (.A(w1233), .B(w1232), .Z(w254) );
	vdp_and g1575 (.A(w1416), .B(w645), .Z(w1358) );
	vdp_or g1576 (.A(w1359), .B(w1422) );
	vdp_and g1577 (.A(w1319), .B(w1334), .Z(w1398) );
	vdp_and g1578 (.A(w1351), .B(w1334), .Z(w1428) );
	vdp_and g1579 (.A(w1334), .B(w1325), .Z(w115) );
	vdp_and g1580 (.A(w997), .B(w116), .Z(w1411) );
	vdp_or g1581 (.A(w1345), .B(w1001), .Z(w1407) );
	vdp_aon22 g1582 (.Z(w1415), .A2(w1071), .B1(w1352), .B2(w1403), .A1(w1402) );
	vdp_and g1583 (.A(w1410), .B(w1425), .Z(w1133) );
	vdp_and g1584 (.A(w1423), .B(w1432), .Z(w1413) );
	vdp_and g1585 (.A(w1432), .B(w1426), .Z(w1410) );
	vdp_not g1586 (.A(w1426), .nZ(w1423) );
	vdp_not g1587 (.A(w1424), .nZ(w1432) );
	vdp_not g1588 (.A(w1381), .nZ(w1419) );
	vdp_not g1589 (.A(w1396), .nZ(w1414) );
	vdp_and g1590 (.A(w1408), .B(w1372), .Z(w1371) );
	vdp_and g1591 (.A(w1408), .B(w1374), .Z(w996) );
	vdp_and g1592 (.A(w1408), .B(w1376), .Z(w1001) );
	vdp_and g1593 (.A(w1408), .B(w1373), .Z(w997) );
	vdp_and g1594 (.A(w1408), .B(w1375), .Z(w1392) );
	vdp_and g1595 (.A(w996), .B(w1392), .Z(w427) );
	vdp_and g1596 (.A(w406), .B(w1386), .Z(w993) );
	vdp_and g1597 (.A(w406), .B(w1377), .Z(w1035) );
	vdp_not g1598 (.A(w406), .nZ(w1408) );
	vdp_nand g1599 (.A(w1404), .B(w1405), .Z(w1426) );
	vdp_nand g1600 (.A(w1038), .B(w1369), .Z(w1368) );
	vdp_nand g1601 (.A(w406), .B(w254), .Z(w1379) );
	vdp_nand g1602 (.A(w279), .B(w406), .Z(w1378) );
	vdp_or3 g1603 (.C(w1233), .A(w1232), .B(w1231), .Z(w1063) );
	vdp_and3 g1604 (.C(w1359), .A(w592), .B(w1416), .Z(w597) );
	vdp_aoi21 g1605 (.A2(w1358), .B(w1419), .Z(w1357), .A1(w1380) );
	vdp_nor g1606 (.A(w1384), .B(w1427), .Z(w1369) );
	vdp_nand g1607 (.A(w113), .B(w1385), .Z(w1396) );
	vdp_nand3 g1608 (.C(w1368), .A(w3), .B(w1383), .Z(w1367) );
	vdp_2a3oi g1609 (.A1(w1419), .B(w672), .Z(w1366), .A2(w1380), .C(w1416) );
	vdp_nor4 g1610 (.C(VRAM_REFRESH), .A(w1422), .B(w1384), .Z(w1546), .D(w1427) );
	vdp_comb1 g1611 (.A1(CA[15]), .B(w1423), .Z(w1424), .A2(CA[14]), .C(w1371) );
	vdp_aon22 g1612 (.Z(w1342), .A2(w1071), .B1(w1352), .B2(w1397), .A1(w1535) );
	vdp_not g1613 (.A(w1071), .nZ(w1352) );
	vdp_or4 g1614 (.C(w1399), .A(w1432), .B(w1398), .Z(w1535), .D(w1347) );
	vdp_or4 g1615 (.C(w1359), .A(w1414), .B(w1411), .Z(w1403), .D(w1359) );
	vdp_or3 g1616 (.C(w1400), .A(w1410), .B(w1401), .Z(w1397) );
	vdp_comb1 g1617 (.A1(w1134), .B(w1329), .Z(w1536), .A2(w1350), .C(w1334) );
	vdp_and6 g1618 (.C(w1394), .A(w1295), .B(w1393), .Z(w1353), .D(w1364), .E(w406), .F(w1338) );
	vdp_or5 g1619 (.C(w1412), .A(w1404), .B(w47), .Z(w1402), .D(w1348), .E(w1135) );
	vdp_or5 g1620 (.C(w1359), .A(w1413), .B(w114), .Z(w1406), .D(w1347), .E(w1411) );
	vdp_aoi22 g1621 (.Z(w1346), .A2(w47), .B1(w1349), .B2(w1334), .A1(w1350) );
	vdp_g1622 g1622 (.Z(w308), .A(w426) );
	vdp_g1623 g1623 (.Z(w264), .A(w426) );
	vdp_g1624 g1624 (.A(w426), .Z(w300) );
	vdp_g1625 g1625 (.A(w426), .Z(w256) );
	vdp_g1626 g1626 (.Z(w290), .A(w426) );
	vdp_g1627 g1627 (.Z(w247), .A(w426) );
	vdp_g1628 g1628 (.Z(w281), .A(w426) );
	vdp_g1629 g1629 (.Z(w239), .A(w426) );
	vdp_aon22 g1630 (.Z(w1401), .A2(w1358), .B1(w1358), .B2(w1419), .A1(w1359) );
	vdp_comp_we g1631 (.nZ(w1370), .Z(w1391), .A(w1409) );
	vdp_comp_we g1632 (.nZ(w1297), .Z(w1320), .A(w1437) );
	vdp_not g1633 (.nZ(w1626), .A(w1982) );
	vdp_not g1634 (.nZ(w1628), .A(w1629) );
	vdp_sr_bit g1635 (.Q(w5), .D(w1977), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1636 (.Q(w1634), .D(w1831), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1637 (.Q(w1610), .D(w1832), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1638 (.Q(w1666), .D(w1631), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1639 (.Q(w1611), .D(w1833), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1640 (.Q(w1615), .D(w1834), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1641 (.Q(w1810), .D(w1821), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1642 (.Q(w1642), .D(w1640), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1643 (.Q(w1639), .D(w1822), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1644 (.Q(w1616), .D(w1823), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1645 (.Q(w1649), .D(w1848), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1646 (.Q(w1647), .D(w1644), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1647 (.Q(w1644), .D(w1993), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1648 (.Q(w1648), .D(w1651), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1649 (.Q(w1621), .D(w1943), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_not g1650 (.nZ(w1640), .A(w1650) );
	vdp_not g1651 (.nZ(w58), .A(w1639) );
	vdp_not g1652 (.nZ(w1625), .A(w1639) );
	vdp_not g1653 (.nZ(w1618), .A(ODD/EVEN) );
	vdp_not g1654 (.nZ(w1627), .A(LS0) );
	vdp_not g1655 (.nZ(w1993), .A(w1978) );
	vdp_not g1656 (.nZ(w1653), .A(w1654) );
	vdp_not g1657 (.nZ(w1641), .A(w1979) );
	vdp_not g1658 (.nZ(w1646), .A(w1647) );
	vdp_not g1659 (.nZ(w1623), .A(w53) );
	vdp_and g1660 (.Z(w1645), .A(w1844), .B(w1649) );
	vdp_nor g1661 (.Z(w1643), .A(SYSRES), .B(w1615) );
	vdp_oai21 g1662 (.Z(w1978), .B(w1643), .A2(w1653), .A1(w1644) );
	vdp_oai21 g1663 (.Z(w1654), .B(w1652), .A2(w1651), .A1(w1848) );
	vdp_aoi21 g1664 (.Z(w1979), .B(SYSRES), .A2(w1648), .A1(w1844) );
	vdp_and g1665 (.Z(w1622), .A(w1625), .B(w27) );
	vdp_and3 g1666 (.Z(w1844), .A(w1646), .B(w53), .C(w1644) );
	vdp_or g1667 (.Z(w1624), .A(SYSRES), .B(w1625) );
	vdp_and g1668 (.Z(w1943), .A(w1619), .B(w1629) );
	vdp_and g1669 (.Z(w1630), .A(w1622), .B(w1623) );
	vdp_and g1670 (.Z(w1619), .A(w1622), .B(w53) );
	vdp_and g1671 (.Z(w1614), .A(w1609), .B(w1616) );
	vdp_or g1672 (.Z(w1613), .A(SYSRES), .B(w1614) );
	vdp_2?3?I g1673 (.Z(w1982), .A1(w1628), .A2(w1619), .C(SYSRES), .B(w1627) );
	vdp_or g1674 (.Z(w1609), .A(w1617), .B(w1618) );
	vdp_or g1675 (.Z(w1612), .A(SYSRES), .B(w1664) );
	vdp_and g1676 (.Z(w1664), .A(w1609), .B(w1611) );
	vdp_and g1677 (.Z(w1635), .A(w1609), .B(w1634) );
	vdp_and g1678 (.Z(w1633), .A(w1609), .B(w1610) );
	vdp_or g1679 (.Z(w1932), .A(w1664), .B(SYSRES) );
	vdp_and g1680 (.Z(w1850), .A(w1631), .B(M5) );
	vdp_not g1681 (.nZ(w46), .A(w1637) );
	vdp_not g1682 (.nZ(w1637), .A(w1636) );
	vdp_not g1683 (.nZ(w1670), .A(w1636) );
	vdp_not g1684 (.nZ(w1977), .A(w1820) );
	vdp_and g1685 (.Z(w1736), .A(M5), .B(w1632) );
	vdp_or g1686 (.Z(w1638), .A(SYSRES), .B(w1635) );
	vdp_oai21 g1687 (.Z(w1636), .B(w1116), .A2(w31), .A1(w5) );
	vdp_RS g1688 (.Q(w1632), .S(w1633), .R(w1638) );
	vdp_RS g1689 (.Q(w1620), .R(w1612), .S(w1614) );
	vdp_RS g1690 (.Q(w31), .S(w1642), .R(w1624) );
	vdp_RS g1691 (.Q(w20), .R(w1615), .S(w1613) );
	vdp_TFF g1692 (.C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .CI(w1630), .R(w1626), .A(w1621), .Q(ODD/EVEN) );
	vdp_cnt_bit_load g1693 (.D(w1840), .Q(w1702), .nL(w1960), .L(w1825), .CI(w1842), .nC1(nHCLK1), .CO(w1930), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g1694 (.Q(w1617), .D(w1921), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1695 (.Q(w1991), .D(w1939), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1696 (.Q(w32), .D(w2006), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1697 (.Q(w27), .D(w1917), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1698 (.Q(VRAM_REFRESH), .D(w1689), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1699 (.Q(w1704), .D(w1688), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1700 (.Q(w1698), .D(w1687), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1701 (.Q(w1674), .D(w1918), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1702 (.Q(w1699), .D(w1713), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1703 (.Q(w1651), .D(w1920), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1704 (.Q(w1847), .D(w1922), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1705 (.Q(w1728), .D(w1916), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1706 (.Q(w1848), .D(w1912), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1707 (.Q(w1713), .D(w1970), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1708 (.Q(w1866), .D(w1874), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1709 (.Q(w1708), .D(w1685), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1710 (.Q(w1727), .D(w1875), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1711 (.Q(w2004), .D(w2007), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1712 (.Q(w1762), .D(w1758), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1713 (.Q(w1710), .D(w1869), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1714 (.Q(w9), .D(w1868), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1715 (.Q(w1725), .D(w1772), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1716 (.Q(w1722), .D(w1919), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1717 (.Q(w1741), .D(w1873), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1718 (.Q(w1733), .D(w1749), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1719 (.Q(w1793), .D(w1737), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1720 (.Q(w29), .D(w1764), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1721 (.Q(w22), .D(w1671), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1722 (.Q(w1757), .D(w1771), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1723 (.Q(w1972), .D(w1799), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1724 (.Q(w1795), .D(w1870), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1725 (.Q(w1753), .D(w1910), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1726 (.Q(w1779), .D(w1802), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1727 (.Q(w30), .D(w1941), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1728 (.Q(w1781), .D(w1872), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1729 (.Q(w1782), .D(w1871), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1730 (.Q(w1808), .D(w1751), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1731 (.Q(w1754), .D(w1913), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1732 (.Q(w1665), .D(w1998), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1733 (.Q(w1739), .D(w1997), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1734 (.Q(w1794), .D(w1750), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1735 (.Q(w1755), .D(w1752), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1736 (.Q(w1798), .D(w1914), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1737 (.Q(w1776), .D(w1911), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1738 (.Q(w25), .D(w1672), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1739 (.Q(w1777), .D(w1665), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2) );
	vdp_sr_bit g1740 (.Q(w1809), .D(w1763), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_sr_bit g1741 (.Q(w1860), .D(w1909), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_not g1742 (.nZ(w1694), .A(M5) );
	vdp_not g1743 (.nZ(w6), .A(w1945) );
	vdp_not g1744 (.nZ(w7), .A(w1674) );
	vdp_not g1745 (.nZ(w1867), .A(w1669) );
	vdp_not g1746 (.nZ(w1678), .A(w53) );
	vdp_not g1747 (.nZ(w1680), .A(w1940) );
	vdp_not g1748 (.nZ(w1768), .A(w1) );
	vdp_not g1749 (.nZ(w1718), .A(w1686) );
	vdp_not g1750 (.nZ(w1700), .A(w1699) );
	vdp_not g1751 (.nZ(w1711), .A(w1674) );
	vdp_not g1752 (.nZ(w1712), .A(w44) );
	vdp_not g1753 (.nZ(w8), .A(w1706) );
	vdp_not g1754 (.nZ(w1696), .A(w39) );
	vdp_not g1755 (.nZ(w2003), .A(w53) );
	vdp_not g1756 (.nZ(w13), .A(w1966) );
	vdp_not g1757 (.nZ(w1967), .A(w1722) );
	vdp_not g1758 (.nZ(w1970), .A(w1732) );
	vdp_not g1759 (.nZ(w1767), .A(w1691) );
	vdp_not g1760 (.nZ(w1989), .A(w1690) );
	vdp_not g1761 (.nZ(w1716), .A(H40) );
	vdp_not g1762 (.nZ(w14), .A(w1765) );
	vdp_not g1763 (.nZ(w1959), .A(w1677) );
	vdp_not g1764 (.nZ(w1805), .A(w1735) );
	vdp_not g1765 (.nZ(w1783), .A(w1769) );
	vdp_not g1766 (.nZ(w1800), .A(w52) );
	vdp_not g1767 (.nZ(w1745), .A(w1915) );
	vdp_not g1768 (.nZ(w12), .A(w1946) );
	vdp_not g1769 (.nZ(w1811), .A(w1809) );
	vdp_not g1770 (.nZ(w1709), .A(w42) );
	vdp_not g1771 (.nZ(w1726), .A(w51) );
	vdp_not g1772 (.nZ(w1675), .A(w41) );
	vdp_not g1773 (.nZ(w1931), .A(w19) );
	vdp_not g1774 (.nZ(w1990), .A(w45) );
	vdp_not g1775 (.nZ(w1992), .A(M5) );
	vdp_not g1776 (.nZ(w1985), .A(w1746) );
	vdp_not g1777 (.nZ(w1824), .A(w1774) );
	vdp_not g1778 (.nZ(w1963), .A(w1938) );
	vdp_not g1779 (.nZ(w1826), .A(w1092) );
	vdp_not g1780 (.nZ(w1843), .A(w1841) );
	vdp_not g1781 (.nZ(w1837), .A(w1495) );
	vdp_not g1782 (.nZ(w1838), .A(PAL) );
	vdp_aon22 g1783 (.Z(w2012), .B1(w1828), .A1(w1827), .A2(DB[4]), .B2(w1826) );
	vdp_aon22 g1784 (.Z(w1952), .B1(w1828), .A1(w1827), .A2(DB[5]), .B2(w1815) );
	vdp_aon22 g1785 (.Z(w1953), .B1(w1828), .A1(w1827), .B2(w1963), .A2(DB[6]) );
	vdp_aon22 g1786 (.Z(w1949), .B2(1'b1), .A2(DB[7]), .B1(w1828), .A1(w1827) );
	vdp_aon22 g1787 (.Z(w1948), .B2(1'b1), .A2(DB[8]), .B1(w1828), .A1(w1827) );
	vdp_aon22 g1788 (.Z(w1817), .B2(1'b1), .B1(w1676), .A2(DB[8]), .A1(w1942) );
	vdp_aon22 g1789 (.Z(w1962), .B2(w1814), .A2(DB[3]), .B1(w1828), .A1(w1827) );
	vdp_aon22 g1790 (.Z(w1835), .A2(DB[2]), .B2(w1838), .B1(w1828), .A1(w1827) );
	vdp_aon22 g1791 (.Z(w1836), .A2(DB[1]), .B2(w1813), .B1(w1828), .A1(w1827) );
	vdp_aon22 g1792 (.Z(w1954), .A1(w1942), .B1(w1676), .B2(1'b1), .A2(DB[7]) );
	vdp_aon22 g1793 (.Z(w21), .A1(w1992), .B2(w1816), .B1(M5), .A2(w1793) );
	vdp_aon22 g1794 (.Z(w1786), .B1(w1676), .A1(w1942), .A2(DB[6]), .B2(1'b1) );
	vdp_aon22 g1795 (.Z(w1761), .B1(w1777), .B2(w1778), .A2(w1861), .A1(w1775) );
	vdp_not g1796 (.nZ(w1778), .A(w1775) );
	vdp_aon22 g1797 (.Z(w1955), .B1(w1676), .A1(w1942), .B2(1'b0), .A2(DB[5]) );
	vdp_not g1798 (.nZ(w1806), .A(w1803) );
	vdp_aon22 g1799 (.Z(w1999), .B1(w1942), .A1(w1676), .B2(w1959), .A2(DB[4]) );
	vdp_aon22 g1800 (.Z(w1956), .B2(w1958), .B1(w1676), .A2(DB[3]), .A1(w1942) );
	vdp_aon22 g1801 (.Z(w1759), .A2(w1694), .B2(M5), .A1(w1761), .B1(w1760) );
	vdp_aon22 g1802 (.Z(w1957), .A2(DB[2]), .B2(w1729), .A1(w1942), .B1(w1676) );
	vdp_aon22 g1803 (.Z(w1968), .B2(w1866), .B1(w44), .A2(w1712), .A1(w1711) );
	vdp_aon22 g1804 (.Z(w1703), .B1(w1944), .A1(HCLK2), .B2(w1696), .A2(w39) );
	vdp_aon22 g1805 (.Z(w1983), .A1(w1942), .B1(w1676), .B2(w1714), .A2(DB[1]) );
	vdp_aon22 g1806 (.Z(w1681), .A2(DB[0]), .B1(w1676), .B2(w1677), .A1(w1942) );
	vdp_not g1807 (.nZ(w4), .A(w1847) );
	vdp_not g1808 (.nZ(w3), .A(w1710) );
	vdp_RS g1809 (.Q(w1756), .S(w1807), .R(w1934) );
	vdp_RS g1810 (.Q(w1804), .R(w1795), .S(w1797) );
	vdp_RS g1811 (.Q(w1737), .S(w1973), .R(w1755) );
	vdp_RS g1812 (.Q(w1933), .R(w2002), .S(w1733) );
	vdp_RS g1813 (.Q(w1738), .R(w1728), .S(w1996) );
	vdp_aon22 g1814 (.Z(w1840), .A2(DB[0]), .B2(w1812), .B1(w1828), .A1(w1827) );
	vdp_notif0 g1815 (.nZ(DB[1]), .A(VRAM_REFRESH), .nE(w1692) );
	vdp_notif0 g1816 (.nZ(DB[0]), .A(w32), .nE(w1692) );
	vdp_notif0 g1817 (.nZ(DB[7]), .A(w27), .nE(w1693) );
	vdp_notif0 g1818 (.A(w7), .nZ(DB[6]), .nE(w1693) );
	vdp_notif0 g1819 (.A(w6), .nZ(DB[2]), .nE(w1692) );
	vdp_notif0 g1820 (.A(w8), .nZ(DB[3]), .nE(w1692) );
	vdp_notif0 g1821 (.nZ(DB[5]), .A(w14), .nE(w1692) );
	vdp_notif0 g1822 (.A(w13), .nZ(DB[4]), .nE(w1692) );
	vdp_notif0 g1823 (.A(w16), .nZ(DB[5]), .nE(w1693) );
	vdp_notif0 g1824 (.nZ(DB[7]), .A(w9), .nE(w1692) );
	vdp_notif0 g1825 (.nZ(DB[6]), .A(w3), .nE(w1692) );
	vdp_notif0 g1826 (.nZ(DB[4]), .A(w17), .nE(w1693) );
	vdp_notif0 g1827 (.nZ(DB[9]), .A(w29), .nE(w1692) );
	vdp_notif0 g1828 (.nZ(DB[8]), .A(w22), .nE(w1692) );
	vdp_notif0 g1829 (.nZ(DB[3]), .A(w11), .nE(w1693) );
	vdp_notif0 g1830 (.nZ(DB[2]), .A(w28), .nE(w1693) );
	vdp_notif0 g1831 (.nZ(DB[10]), .A(w30), .nE(w1692) );
	vdp_notif0 g1832 (.nZ(DB[11]), .A(w12), .nE(w1692) );
	vdp_notif0 g1833 (.nZ(DB[12]), .A(w24), .nE(w1692) );
	vdp_notif0 g1834 (.nZ(DB[13]), .A(w25), .nE(w1692) );
	vdp_notif0 g1835 (.nZ(DB[1]), .A(w15), .nE(w1693) );
	vdp_notif0 g1836 (.nZ(DB[0]), .A(w10), .nE(w1693) );
	vdp_not g1837 (.nZ(VPOS[9]), .A(w1951) );
	vdp_not g1838 (.nZ(VPOS[8]), .A(w1950) );
	vdp_not g1839 (.nZ(VPOS[7]), .A(w1747) );
	vdp_not g1840 (.nZ(HPOS[7]), .A(w1985) );
	vdp_not g1841 (.nZ(HPOS[8]), .A(w1824) );
	vdp_not g1842 (.nZ(HPOS[6]), .A(w1745) );
	vdp_not g1843 (.nZ(VPOS[6]), .A(w1986) );
	vdp_not g1844 (.nZ(VPOS[5]), .A(w1987) );
	vdp_not g1845 (.nZ(HPOS[5]), .A(w1783) );
	vdp_not g1846 (.nZ(HPOS[4]), .A(w1805) );
	vdp_not g1847 (.nZ(VPOS[4]), .A(w1988) );
	vdp_not g1848 (.nZ(HPOS[3]), .A(w1989) );
	vdp_not g1849 (.nZ(VPOS[3]), .A(w1730) );
	vdp_not g1850 (.nZ(HPOS[2]), .A(w1767) );
	vdp_not g1851 (.nZ(VPOS[2]), .A(w1719) );
	vdp_not g1852 (.nZ(HPOS[1]), .A(w1718) );
	vdp_not g1853 (.nZ(VPOS[1]), .A(w1679) );
	vdp_not g1854 (.nZ(HPOS[0]), .A(w1680) );
	vdp_not g1855 (.nZ(VPOS[0]), .A(w1673) );
	vdp_aoi22 g1856 (.Z(w1944), .A1(w1666), .B1(w1695), .B2(M5), .A2(w1694) );
	vdp_aon22 g1857 (.Z(w1720), .A2(w1694), .B1(w1721), .B2(M5), .A1(w1763) );
	vdp_aoi22 g1858 (.Z(w1673), .B2(w1768), .B1(w1702), .A1(ODD/EVEN), .A2(w1) );
	vdp_aoi22 g1859 (.Z(w1679), .B2(w1768), .B1(w1845), .A1(w1702), .A2(w1) );
	vdp_aoi22 g1860 (.Z(w1719), .A2(w1), .A1(w1845), .B2(w1768), .B1(w1937) );
	vdp_aoi22 g1861 (.Z(w1730), .A1(w1937), .B2(w1768), .A2(w1), .B1(w1830) );
	vdp_aoi22 g1862 (.Z(w1988), .B1(w1936), .A1(w1830), .A2(w1), .B2(w1768) );
	vdp_aoi22 g1863 (.Z(w1987), .B1(w1785), .A1(w1936), .A2(w1), .B2(w1768) );
	vdp_aoi22 g1864 (.Z(w1986), .A2(w1), .B2(w1768), .B1(w1748), .A1(w1785) );
	vdp_aoi22 g1865 (.Z(w1747), .B2(w1768), .A1(w1748), .B1(w1819), .A2(w1) );
	vdp_aoi22 g1866 (.Z(w1950), .B2(w1768), .A2(w1), .A1(w1819), .B1(w1846) );
	vdp_aoi22 g1867 (.Z(w1951), .B1(1'b0), .A2(w1), .B2(w1768), .A1(w1846) );
	vdp_comp_ g1868 (.Q(w1652), .D(w1697), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_comp_ g1869 (.Q(w1801), .D(w1974), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2) );
	vdp_cnt_bit g1870 (.CI(w1976), .Q(w1861), .nEN(SYSRES), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_not g1871 (.nZ(w1947), .A(w55) );
	vdp_and g1872 (.Z(w1788), .A(w1803), .B(w1738) );
	vdp_and g1873 (.Z(w1789), .A(w1803), .B(w1738) );
	vdp_and g1874 (.Z(w1791), .A(w2001), .B(w1804) );
	vdp_and g1875 (.Z(w1792), .A(w1804), .B(w1806) );
	vdp_and g1876 (.Z(w1790), .A(w1850), .B(w1756) );
	vdp_and g1877 (.Z(w2001), .A(w1849), .B(w1736) );
	vdp_and g1878 (.Z(w1729), .A(w53), .B(w1716) );
	vdp_and g1879 (.Z(w16), .A(w1968), .B(w1707) );
	vdp_and g1880 (.Z(w1714), .A(w1678), .B(w1716) );
	vdp_and g1881 (.Z(w26), .A(w1637), .B(w1933) );
	vdp_and g1882 (.Z(w1715), .A(w52), .B(w1801) );
	vdp_and g1883 (.Z(w1740), .A(w1931), .B(w53) );
	vdp_and g1884 (.Z(w15), .A(w1707), .B(w1798) );
	vdp_and g1885 (.Z(w1773), .A(w1990), .B(w1740) );
	vdp_and g1886 (.Z(w10), .A(w1860), .B(w1707) );
	vdp_and g1887 (.Z(w1961), .A(w1810), .B(w4) );
	vdp_or g1888 (.Z(w1815), .A(w1935), .B(w1938) );
	vdp_or g1889 (.Z(w1814), .A(w1964), .B(w1938) );
	vdp_and g1890 (.Z(w1775), .A(M5), .B(w23) );
	vdp_and g1891 (.Z(w1976), .A(w1811), .B(w1763) );
	vdp_or g1892 (.Z(w1797), .A(SYSRES), .B(w1796) );
	vdp_or g1893 (.Z(w28), .A(w1782), .B(w1781) );
	vdp_or g1894 (.Z(w24), .A(w1776), .B(w1782) );
	vdp_or g1895 (.Z(w1998), .A(w1788), .B(w1792) );
	vdp_or g1896 (.Z(w1807), .A(w1794), .B(w1753) );
	vdp_or g1897 (.Z(w1934), .A(SYSRES), .B(w1796) );
	vdp_or g1898 (.Z(w1796), .A(w1741), .B(w1808) );
	vdp_or g1899 (.Z(w1973), .A(w1754), .B(SYSRES) );
	vdp_or g1900 (.Z(w1958), .A(w1677), .B(w2000) );
	vdp_or g1901 (.Z(w2002), .A(SYSRES), .B(w1753) );
	vdp_or g1902 (.Z(w1971), .A(w1715), .B(w1652) );
	vdp_or g1903 (.Z(w1919), .A(w1972), .B(w1799) );
	vdp_and g1904 (.Z(w11), .A(w1757), .B(w1707) );
	vdp_and g1905 (.Z(w1799), .A(w1667), .B(w1740) );
	vdp_or g1906 (.Z(w1996), .A(SYSRES), .B(w1741) );
	vdp_not g1907 (.nZ(w1693), .A(w54) );
	vdp_not g1908 (.nZ(w1692), .A(w48) );
	vdp_aon33 g1909 (.Z(w1842), .A3(w1841), .A2(w1947), .A1(w4), .B1(w55), .B3(1'b1), .B2(w1241) );
	vdp_aoi21 g1910 (.Z(w1945), .A1(w1698), .A2(w1707), .B(w1668) );
	vdp_aoi21 g1911 (.Z(w1706), .A1(w1704), .B(w1705), .A2(w1707) );
	vdp_aoi21 g1912 (.Z(w1669), .A1(w40), .A2(w50), .B(w1701) );
	vdp_aoi21 g1913 (.Z(w1732), .A1(w1713), .B(w1969), .A2(w1971) );
	vdp_aoi21 g1914 (.Z(w1966), .A1(w1707), .B(w1965), .A2(w1708) );
	vdp_aoi21 g1915 (.Z(w1765), .B(w1975), .A1(w1707), .A2(w1727) );
	vdp_aoi21 g1916 (.Z(w1946), .A1(w1707), .A2(w1779), .B(w1780) );
	vdp_xor g1917 (.Z(w1763), .B(w1666), .A(w1739) );
	vdp_xor g1918 (.Z(w1812), .A(ODD/EVEN), .B(w1838) );
	vdp_and3 g1919 (.Z(w1668), .A(w1726), .B(w42), .C(w1675) );
	vdp_and3 g1920 (.Z(w2006), .A(w2005), .B(w1865), .C(w1723) );
	vdp_and3 g1921 (.Z(w1705), .A(w1709), .B(w51), .C(w1675) );
	vdp_and3 g1922 (.Z(w1965), .A(w51), .B(w1675), .C(w42) );
	vdp_and3 g1923 (.Z(w1975), .A(w1709), .B(w1726), .C(w1782) );
	vdp_and3 g1924 (.Z(w1780), .A(w42), .B(w1726), .C(w41) );
	vdp_or3 g1925 (.Z(w1997), .A(w1790), .B(w1791), .C(w1789) );
	vdp_and3 g1926 (.Z(w2000), .A(w53), .B(w1716), .C(M5) );
	vdp_and3 g1927 (.Z(w1876), .A(w1713), .B(w53), .C(w1700) );
	vdp_and3 g1928 (.Z(w1677), .A(H40), .B(M5), .C(w1678) );
	vdp_nor4 g1929 (.Z(w1723), .A(w1766), .B(w1802), .C(w1671), .D(w1764) );
	vdp_nor4 g1930 (.Z(w1841), .A(w56), .B(w1844), .D(w1961), .C(SYSRES) );
	vdp_comp_we g1931 (.Z(w1825), .nZ(w1960), .A(w1843) );
	vdp_comp_we g1932 (.Z(w1827), .nZ(w1828), .A(w56) );
	vdp_comp_we g1933 (.Z(w1942), .nZ(w1676), .A(w57) );
	vdp_comp_we g1934 (.Z(w1683), .nZ(w1682), .A(w1667) );
	vdp_and3 g1935 (.Z(w18), .A(w1116), .B(w1933), .C(w31) );
	vdp_or4 g1936 (.Z(w1667), .A(w57), .B(SYSRES), .C(w1876), .D(w1991) );
	vdp_nor3 g1937 (.Z(w1865), .A(w1868), .B(w1724), .C(w1875) );
	vdp_nor3 g1938 (.Z(w1803), .A(w1736), .B(w1850), .C(w1849) );
	vdp_nand g1939 (.Z(w1758), .A(w1759), .B(w1800) );
	vdp_nand g1940 (.Z(w2007), .A(w1720), .B(w2003) );
	vdp_nand g1941 (.Z(w1869), .A(w1967), .B(w1724) );
	vdp_nor3 g1942 (.Z(w1707), .A(w42), .B(w51), .C(w41) );
	vdp_nor g1943 (.Z(w1938), .A(w1838), .B(M5) );
	vdp_nor g1944 (.Z(w1813), .A(ODD/EVEN), .B(w1838) );
	vdp_nor g1945 (.Z(w1935), .A(w1826), .B(PAL) );
	vdp_nor g1946 (.Z(w1964), .A(w1826), .B(w1838) );
	vdp_nor g1947 (.Z(w1969), .A(w1651), .B(SYSRES) );
	vdp_SDELAY8 g1948 (.Q(w1816), .D(w1793), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2), .nC3(nHCLK1), .C3(HCLK1), .nC4(nHCLK2), .C4(HCLK2), .nC5(nHCLK1), .C5(HCLK1), .nC6(nHCLK2), .C6(HCLK2), .nC7(nHCLK1), .C7(HCLK1), .nC8(nHCLK2), .C8(HCLK2), .nC9(nHCLK1), .C9(HCLK1), .nC10(nHCLK2), .C10(HCLK2), .nC11(nHCLK1), .C11(HCLK1), .nC12(nHCLK2), .C12(HCLK2), .nC13(nHCLK1), .C13(HCLK1), .nC14(nHCLK2), .C14(HCLK2), .nC15(nHCLK1), .C15(HCLK1), .nC16(nHCLK2), .C16(HCLK2) );
	vdp_SDELAY7 g1949 (.Q(w1760), .D(w1761), .C1(HCLK1), .nC1(nHCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .nC4(nHCLK2), .C5(HCLK1), .nC5(nHCLK1), .C6(HCLK2), .nC6(nHCLK2), .C7(HCLK1), .nC7(nHCLK1), .C8(HCLK2), .nC8(nHCLK2), .C9(HCLK1), .nC9(nHCLK1), .C10(HCLK2), .nC10(nHCLK2), .C11(HCLK1), .nC11(nHCLK1), .C12(HCLK2), .nC12(nHCLK2), .C13(HCLK1), .nC13(nHCLK1), .C14(HCLK2), .nC14(nHCLK2), .C3(HCLK1) );
	vdp_SDELAY8 g1950 (.Q(w1721), .D(w1763), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2), .C3(HCLK1), .nC4(nHCLK2), .C4(HCLK2), .nC5(nHCLK1), .C5(HCLK1), .nC6(nHCLK2), .C6(HCLK2), .nC7(nHCLK1), .C7(HCLK1), .nC8(nHCLK2), .C8(HCLK2), .nC9(nHCLK1), .C9(HCLK1), .nC10(nHCLK2), .C10(HCLK2), .C11(HCLK1), .nC12(nHCLK2), .C12(HCLK2), .nC13(nHCLK1), .C13(HCLK1), .nC14(nHCLK2), .C14(HCLK2), .nC15(nHCLK1), .C15(HCLK1), .nC16(nHCLK2), .C16(HCLK2), .nC3(nHCLK1), .nC11(nHCLK1) );
	vdp_SDELAY8 g1951 (.Q(w1695), .D(w1666), .nC1(nHCLK1), .C1(HCLK1), .nC2(nHCLK2), .C2(HCLK2), .C3(HCLK1), .nC4(nHCLK2), .C4(HCLK2), .nC5(nHCLK1), .C5(HCLK1), .nC6(nHCLK2), .C6(HCLK2), .nC7(nHCLK1), .C7(HCLK1), .nC8(nHCLK2), .C8(HCLK2), .nC9(nHCLK1), .C9(HCLK1), .nC10(nHCLK2), .C10(HCLK2), .nC11(nHCLK1), .C11(HCLK1), .nC12(nHCLK2), .C12(HCLK2), .nC13(nHCLK1), .C13(HCLK1), .nC14(nHCLK2), .C14(HCLK2), .nC15(nHCLK1), .C15(HCLK1), .nC16(nHCLK2), .C16(HCLK2), .nC3(nHCLK1) );
	vdp_cnt_bit_load g1952 (.D(w1836), .Q(w1845), .nL(w1960), .L(w1825), .CI(w1930), .nC1(nHCLK1), .CO(w2009), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1953 (.D(w1835), .Q(w1937), .nL(w1960), .L(w1825), .CI(w2009), .nC1(nHCLK1), .CO(w2010), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1954 (.D(w1962), .Q(w1830), .nL(w1960), .L(w1825), .CI(w2010), .nC1(nHCLK1), .CO(w2011), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1955 (.D(w2012), .Q(w1936), .nL(w1960), .L(w1825), .CI(w2011), .nC1(nHCLK1), .CO(w1864), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1956 (.D(w1952), .Q(w1785), .nL(w1960), .L(w1825), .CI(w1864), .nC1(nHCLK1), .CO(w1863), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1957 (.D(w1953), .Q(w1748), .nL(w1960), .L(w1825), .CI(w1863), .nC1(nHCLK1), .CO(w2013), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1958 (.D(w1949), .Q(w1819), .nL(w1960), .L(w1825), .CI(w2013), .nC1(nHCLK1), .CO(w1862), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1959 (.D(w1948), .Q(w1846), .nL(w1960), .L(w1825), .CI(w1862), .nC1(nHCLK1), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1960 (.D(w1817), .Q(w1774), .nL(w1742), .L(w1683), .CI(w1818), .nC1(nHCLK1), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1961 (.D(w1954), .Q(w1746), .nL(w1742), .L(w1683), .CI(w1744), .nC1(nHCLK1), .CO(w1818), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1962 (.D(w1786), .Q(w1915), .nL(w1742), .L(w1683), .CI(w1784), .nC1(nHCLK1), .CO(w1744), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1963 (.D(w1955), .Q(w1769), .nL(w1742), .L(w1683), .CI(w1770), .nC1(nHCLK1), .CO(w1784), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1964 (.D(w1999), .Q(w1735), .nL(w1742), .L(w1683), .CI(w1734), .nC1(nHCLK1), .CO(w1770), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1965 (.D(w1956), .Q(w1690), .nL(w1682), .L(w1683), .CI(w1731), .nC1(nHCLK1), .CO(w1734), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1966 (.D(w1957), .Q(w1691), .nL(w1682), .L(w1683), .CI(w1717), .nC1(nHCLK1), .CO(w1731), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1967 (.D(w1983), .Q(w1686), .nL(w1682), .L(w1683), .CI(w2008), .nC1(nHCLK1), .CO(w1717), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g1968 (.D(w1681), .Q(w1940), .nL(w1682), .L(w1683), .CI(w1867), .nC1(nHCLK1), .CO(w2008), .R(1'b0), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_or8 g1969 (.Z(w1831), .A(w1877), .B(w1878), .C(w1879), .D(w1880), .E(w1927), .F(w1928), .G(w1929), .H(w1882) );
	vdp_or8 g1970 (.Z(w1832), .A(w1883), .B(w1926), .C(w1925), .D(w1908), .E(w1924), .F(w1884), .G(w1885), .H(w1923) );
	vdp_or8 g1971 (.Z(w1833), .A(w2014), .B(w1994), .C(w1995), .D(w1981), .E(w1907), .F(w1906), .G(w1980), .H(w1905) );
	vdp_or5 g1972 (.Z(w1834), .A(w1901), .B(w1902), .C(w1903), .D(w1904), .E(w6821) );
	vdp_or7 g1973 (.Z(w1823), .A(w1897), .B(w1898), .C(w1899), .D(w1900), .E(w6818), .F(w6819), .G(w6820) );
	vdp_or7 g1974 (.Z(w1821), .A(w1886), .B(w1887), .C(w1888), .D(w1889), .E(w1890), .F(w1891), .G(w1892) );
	vdp_nor g1975 (.Z(w1701), .A(w1667), .B(w40) );
	vdp_and g1976 (.Z(w17), .A(w1707), .B(w1725) );
	vdp_not g1977 (.nZ(w1650), .A(w1893) );
	vdp_nor3 g1978 (.Z(w1822), .A(w1896), .B(w1895), .C(w1894) );
	vdp_RS g1979 (.S(w1932), .R(w1633), .Q(w1631) );
	vdp_RS g1980 (.S(w1645), .R(w1641), .Q(w1629) );
	vdp_and g1981 (.Z(w1849), .A(w1620), .B(M5) );
	vdp_nor4 g1982 (.Z(w2005), .A(w1689), .B(w1688), .C(w1687), .D(w1685) );
	vdp_nand3 g1983 (.A(w2135), .B(w2134), .C(w2132), .Z(w2128) );
	vdp_nand3 g1984 (.A(w2132), .B(w2134), .C(w2137), .Z(w2123) );
	vdp_nand3 g1985 (.A(w2132), .B(w2135), .C(w2136), .Z(w2124) );
	vdp_nand3 g1986 (.A(w2136), .B(w2132), .C(w2137), .Z(w2125) );
	vdp_nand3 g1987 (.A(w2136), .B(w2133), .C(w2137), .Z(w2120) );
	vdp_nand3 g1988 (.A(w2133), .B(w2135), .C(w2136), .Z(w2119) );
	vdp_nand3 g1989 (.A(w2134), .B(w2133), .C(w2137), .Z(w2127) );
	vdp_nand3 g1990 (.A(w2135), .B(w2134), .C(w2133), .Z(w2126) );
	vdp_nand3 g1991 (.A(w2108), .B(w2109), .C(w2104), .Z(w2118) );
	vdp_nand3 g1992 (.A(w2104), .B(w2109), .C(w2107), .Z(w2117) );
	vdp_nand3 g1993 (.A(w2106), .B(w2105), .C(w2107), .Z(w2111) );
	vdp_nand3 g1994 (.A(w2105), .B(w2108), .C(w2106), .Z(w2112) );
	vdp_nand3 g1995 (.A(w2109), .B(w2105), .C(w2107), .Z(w2113) );
	vdp_nand3 g1996 (.A(w2108), .B(w2109), .C(w2105), .Z(w2114) );
	vdp_nand3 g1997 (.A(w2106), .B(w2104), .C(w2107), .Z(w2115) );
	vdp_nand3 g1998 (.A(w2104), .B(w2108), .C(w2106), .Z(w2116) );
	vdp_nand3 g1999 (.A(w2096), .B(w2094), .C(w2092), .Z(w2089) );
	vdp_nand3 g2000 (.A(w2092), .B(w2094), .C(w2097), .Z(w2088) );
	vdp_nand3 g2001 (.A(w2095), .B(w2093), .C(w2097), .Z(w2082) );
	vdp_nand3 g2002 (.A(w2093), .B(w2096), .C(w2095), .Z(w2083) );
	vdp_nand3 g2003 (.A(w2094), .B(w2093), .C(w2097), .Z(w2084) );
	vdp_nand3 g2004 (.A(w2096), .B(w2094), .C(w2093), .Z(w2085) );
	vdp_nand3 g2005 (.A(w2095), .B(w2092), .C(w2097), .Z(w2086) );
	vdp_nand3 g2006 (.A(w2092), .B(w2096), .C(w2095), .Z(w2087) );
	vdp_nand3 g2007 (.A(w2035), .B(w2032), .C(w2036), .Z(w2029) );
	vdp_nand3 g2008 (.A(w2036), .B(w2032), .C(w2034), .Z(w2028) );
	vdp_nand3 g2009 (.A(w2033), .B(w2031), .C(w2034), .Z(w2022) );
	vdp_nand3 g2010 (.A(w2031), .B(w2035), .C(w2033), .Z(w2023) );
	vdp_nand3 g2011 (.A(w2032), .B(w2031), .C(w2034), .Z(w2024) );
	vdp_nand3 g2012 (.A(w2035), .B(w2032), .C(w2031), .Z(w2025) );
	vdp_nand3 g2013 (.A(w2033), .B(w2036), .C(w2034), .Z(w2026) );
	vdp_nand3 g2014 (.A(w2036), .B(w2035), .C(w2033), .Z(w2027) );
	vdp_not g2015 (.nZ(w2030), .A(w2017) );
	vdp_not g2016 (.nZ(w2090), .A(w2016) );
	vdp_not g2017 (.nZ(w2098), .A(w2018) );
	vdp_not g2018 (.nZ(w2129), .A(w2015) );
	vdp_nand g2019 (.Z(w2020), .B(w2021), .A(w2030) );
	vdp_nand g2020 (.Z(w2021), .B(w2030), .A(w2037) );
	vdp_nand g2021 (.Z(w2080), .B(w2081), .A(w2090) );
	vdp_nand g2022 (.Z(w2081), .B(w2090), .A(w2041) );
	vdp_comp_we g2023 (.A(w2091), .Z(w2093), .nZ(w2092) );
	vdp_comp_we g2024 (.A(w2151), .Z(w2095), .nZ(w2094) );
	vdp_comp_we g2025 (.A(w2150), .Z(w2097), .nZ(w2096) );
	vdp_comp_we g2026 (.A(w2038), .Z(w2031), .nZ(w2036) );
	vdp_comp_we g2027 (.A(w2039), .Z(w2033), .nZ(w2032) );
	vdp_comp_we g2028 (.A(w2040), .Z(w2034), .nZ(w2035) );
	vdp_nand g2029 (.Z(w2099), .B(w2098), .A(w2102) );
	vdp_comp_we g2030 (.A(w2101), .Z(w2105), .nZ(w2104) );
	vdp_comp_we g2031 (.A(w2103), .Z(w2106), .nZ(w2109) );
	vdp_comp_we g2032 (.A(w2110), .Z(w2107), .nZ(w2108) );
	vdp_nand g2033 (.Z(w2100), .B(w2099), .A(w2098) );
	vdp_nand g2034 (.Z(w2121), .B(w2129), .A(w2130) );
	vdp_comp_we g2035 (.A(w2131), .Z(w2133), .nZ(w2132) );
	vdp_comp_we g2036 (.A(w2138), .Z(w2136), .nZ(w2134) );
	vdp_comp_we g2037 (.A(w2139), .Z(w2137), .nZ(w2135) );
	vdp_nand g2038 (.Z(w2122), .B(w2121), .A(w2129) );
	vdp_comp_str g2039 (.A(w2162), .Z(w2163), .nZ(w2161) );
	vdp_comp_str g2040 (.A(w2179), .Z(w2152), .nZ(w2153) );
	vdp_comp_str g2041 (.A(w2188), .Z(w2143), .nZ(w2142) );
	vdp_comp_str g2042 (.A(w2189), .Z(w2044), .nZ(w2043) );
	vdp_comp_str g2043 (.A(w2052), .Z(w2053), .nZ(w2054) );
	vdp_comp_str g2044 (.A(w2226), .Z(w2412), .nZ(w2289) );
	vdp_comp_str g2045 (.A(w2437), .Z(w2405), .nZ(w2404) );
	vdp_comp_str g2046 (.A(w2408), .Z(w2418), .nZ(w2406) );
	vdp_comp_str g2047 (.A(w2197), .Z(w2409), .nZ(w2407) );
	vdp_comp_str g2048 (.A(w2317), .Z(w2060), .nZ(w2064) );
	vdp_comp_str g2049 (.A(w2438), .Z(w2061), .nZ(w2065) );
	vdp_comp_str g2050 (.A(w2195), .Z(w2063), .nZ(w2066) );
	vdp_dlatch g2051 (.Q(w2422), .C(w2063), .D(w2190), .nC(w2066) );
	vdp_dlatch g2052 (.Q(w2421), .C(w2061), .D(w2190), .nC(w2065) );
	vdp_dlatch g2053 (.Q(w2384), .C(w2063), .D(w2324), .nC(w2066) );
	vdp_dlatch g2054 (.Q(w2420), .C(w2060), .D(w2190), .nC(w2064) );
	vdp_dlatch g2055 (.Q(w2425), .C(w2063), .D(w2325), .nC(w2066) );
	vdp_dlatch g2056 (.Q(w2383), .C(w2060), .D(w2324), .nC(w2064) );
	vdp_dlatch g2057 (.Q(w2385), .C(w2061), .D(w2324), .nC(w2065) );
	vdp_dlatch g2058 (.Q(w2319), .C(w2063), .D(w2327), .nC(w2066) );
	vdp_dlatch g2059 (.Q(w2423), .C(w2060), .D(w2325), .nC(w2064) );
	vdp_dlatch g2060 (.Q(w2424), .C(w2061), .D(w2325), .nC(w2065) );
	vdp_dlatch g2061 (.Q(w2073), .C(w2063), .D(w2062), .nC(w2066) );
	vdp_dlatch g2062 (.Q(w2318), .C(w2060), .D(w2327), .nC(w2064) );
	vdp_dlatch g2063 (.Q(w2320), .C(w2061), .D(w2327), .nC(w2065) );
	vdp_dlatch g2064 (.Q(w2070), .C(w2060), .D(w2062), .nC(w2064) );
	vdp_dlatch g2065 (.Q(w2072), .C(w2061), .D(w2062), .nC(w2065) );
	vdp_dlatch g2066 (.Q(w2067), .C(w2063), .D(w2059), .nC(w2066) );
	vdp_dlatch g2067 (.Q(w2079), .C(w2060), .D(w2059), .nC(w2064) );
	vdp_dlatch g2068 (.Q(w2068), .C(w2061), .D(w2059), .nC(w2065) );
	vdp_dlatch g2069 (.Q(w2398), .C(w2409), .D(w2190), .nC(w2407) );
	vdp_dlatch g2070 (.Q(w2397), .C(w2418), .D(w2190), .nC(w2406) );
	vdp_dlatch g2071 (.Q(w2403), .C(w2409), .D(w2324), .nC(w2407) );
	vdp_dlatch g2072 (.Q(w2399), .C(w2405), .D(w2190), .nC(w2404) );
	vdp_dlatch g2073 (.Q(w2391), .C(w2409), .D(w2325), .nC(w2407) );
	vdp_dlatch g2074 (.Q(w2401), .C(w2405), .D(w2324), .nC(w2404) );
	vdp_dlatch g2075 (.Q(w2402), .C(w2418), .D(w2324), .nC(w2406) );
	vdp_dlatch g2076 (.Q(w2388), .C(w2409), .D(w2327), .nC(w2407) );
	vdp_dlatch g2077 (.Q(w2389), .C(w2405), .D(w2325), .nC(w2404) );
	vdp_dlatch g2078 (.Q(w2390), .C(w2418), .D(w2325), .nC(w2406) );
	vdp_dlatch g2079 (.Q(w2386), .C(w2405), .D(w2327), .nC(w2404) );
	vdp_dlatch g2080 (.Q(w2387), .C(w2418), .D(w2327), .nC(w2406) );
	vdp_dlatch g2081 (.Q(w2273), .C(w2412), .D(w2325), .nC(w2289) );
	vdp_dlatch g2082 (.Q(w2415), .C(w2412), .D(w2324), .nC(w2289) );
	vdp_dlatch g2083 (.Q(w2416), .C(w2412), .D(w2190), .nC(w2289) );
	vdp_and g2084 (.Z(w2233), .A(w2416), .B(w2415) );
	vdp_and g2085 (.Z(w2400), .A(w2415), .B(w2413) );
	vdp_and g2086 (.Z(w2382), .A(w2416), .B(w2414) );
	vdp_and g2087 (.Z(w2328), .A(w2413), .B(w2414) );
	vdp_dlatch g2088 (.Q(w2165), .C(w2163), .D(w2159), .nC(w2161) );
	vdp_or g2089 (.Z(w2139), .A(w2164), .B(w2165) );
	vdp_notif0 g2090 (.A(w2139), .nZ(DB[0]), .nE(w2045) );
	vdp_dlatch g2091 (.Q(w2448), .C(w2163), .D(w2156), .nC(w2161) );
	vdp_or g2092 (.Z(w2138), .A(w2164), .B(w2448) );
	vdp_notif0 g2093 (.A(w2138), .nZ(DB[1]), .nE(w2045) );
	vdp_dlatch g2094 (.Q(w2449), .C(w2163), .D(w2158), .nC(w2161) );
	vdp_or g2095 (.Z(w2131), .A(w2164), .B(w2449) );
	vdp_notif0 g2096 (.A(w2131), .nZ(DB[2]), .nE(w2045) );
	vdp_dlatch g2097 (.Q(w2169), .C(w2163), .D(w2170), .nC(w2161) );
	vdp_or g2098 (.Z(w2130), .A(w2164), .B(w2169) );
	vdp_notif0 g2099 (.A(w2130), .nZ(DB[3]), .nE(w2045) );
	vdp_dlatch g2100 (.Q(w2160), .C(w2152), .D(w2159), .nC(w2153) );
	vdp_or g2101 (.Z(w2110), .A(w2157), .B(w2160) );
	vdp_notif0 g2102 (.A(w2110), .nZ(DB[4]), .nE(w2045) );
	vdp_dlatch g2103 (.Q(w2155), .C(w2152), .D(w2156), .nC(w2153) );
	vdp_or g2104 (.Z(w2103), .A(w2157), .B(w2155) );
	vdp_notif0 g2105 (.A(w2103), .nZ(DB[5]), .nE(w2045) );
	vdp_dlatch g2106 (.Q(w2154), .C(w2152), .D(w2158), .nC(w2153) );
	vdp_or g2107 (.Z(w2101), .A(w2157), .B(w2154) );
	vdp_notif0 g2108 (.A(w2101), .nZ(DB[6]), .nE(w2045) );
	vdp_dlatch g2109 (.Q(w2149), .C(w2152), .D(w2170), .nC(w2153) );
	vdp_or g2110 (.Z(w2102), .A(w2157), .B(w2149) );
	vdp_notif0 g2111 (.A(w2102), .nZ(DB[7]), .nE(w2045) );
	vdp_dlatch g2112 (.Q(w2447), .C(w2143), .D(w2159), .nC(w2142) );
	vdp_or g2113 (.Z(w2150), .A(w2144), .B(w2447) );
	vdp_notif0 g2114 (.A(w2150), .nZ(DB[8]), .nE(w2045) );
	vdp_dlatch g2115 (.Q(w2148), .C(w2143), .D(w2156), .nC(w2142) );
	vdp_or g2116 (.Z(w2151), .A(w2144), .B(w2148) );
	vdp_notif0 g2117 (.A(w2151), .nZ(DB[9]), .nE(w2045) );
	vdp_dlatch g2118 (.Q(w2141), .C(w2143), .D(w2158), .nC(w2142) );
	vdp_or g2119 (.Z(w2091), .A(w2144), .B(w2141) );
	vdp_notif0 g2120 (.A(w2091), .nZ(DB[10]), .nE(w2045) );
	vdp_dlatch g2121 (.Q(w2140), .C(w2143), .D(w2170), .nC(w2142) );
	vdp_or g2122 (.Z(w2041), .A(w2144), .B(w2140) );
	vdp_notif0 g2123 (.A(w2041), .nZ(DB[11]), .nE(w2045) );
	vdp_dlatch g2124 (.Q(w2046), .C(w2044), .D(w2159), .nC(w2043) );
	vdp_or g2125 (.Z(w2040), .A(w2042), .B(w2046) );
	vdp_notif0 g2126 (.A(w2040), .nZ(DB[12]), .nE(w2045) );
	vdp_dlatch g2127 (.Q(w2047), .C(w2044), .D(w2156), .nC(w2043) );
	vdp_or g2128 (.Z(w2039), .A(w2042), .B(w2047) );
	vdp_notif0 g2129 (.A(w2039), .nZ(DB[13]), .nE(w2045) );
	vdp_dlatch g2130 (.Q(w2048), .C(w2044), .D(w2158), .nC(w2043) );
	vdp_or g2131 (.Z(w2038), .A(w2042), .B(w2048) );
	vdp_notif0 g2132 (.A(w2038), .nZ(DB[14]), .nE(w2045) );
	vdp_dlatch g2133 (.Q(w2049), .C(w2044), .D(w2170), .nC(w2043) );
	vdp_or g2134 (.Z(w2037), .A(w2042), .B(w2049) );
	vdp_notif0 g2135 (.A(w2037), .nZ(DB[15]), .nE(w2045) );
	vdp_not g2136 (.A(PSG_TEST_OE), .nZ(w2045) );
	vdp_not g2137 (.nZ(w2218), .A(w1058) );
	vdp_clkgen g2138 (.PH(w2218), .CLK1(w2219), .nCLK1(w2220), .CLK2(w2221), .nCLK2(w2222) );
	vdp_comp_dff g2139 (.D(SYSRES), .nC1(w2220), .C1(w2219), .C2(w2221), .nC2(w2222), .Q(w2250) );
	vdp_sr_bit g2140 (.D(w2250), .nC1(w2220), .nC2(w2222), .C1(w2219), .C2(w2221), .Q(w2252) );
	vdp_sr_bit g2141 (.D(w2225), .nC1(w2220), .nC2(w2222), .C1(w2219), .C2(w2221), .Q(w2224) );
	vdp_not g2142 (.nZ(w2251), .A(w2252) );
	vdp_and g2143 (.Z(w2223), .A(w2250), .B(w2251) );
	vdp_nor g2144 (.Z(w2225), .A(w2224), .B(w2223) );
	vdp_cnt_bit g2145 (.CI(w2224), .R(w2223), .C1(w2219), .nC1(w2220), .nC2(w2222), .C2(w2221), .Q(w2249) );
	vdp_dlatch_inv g2146 (.nQ(w2248), .D(w2249), .nC(w2220), .C(w2219) );
	vdp_not g2147 (.nZ(w2247), .A(w2248) );
	vdp_nand g2148 (.Z(w2246), .A(w2224), .B(w2248) );
	vdp_not g2149 (.nZ(w2245), .A(w2246) );
	vdp_not g2150 (.nZ(w2244), .A(w2243) );
	vdp_not g2151 (.nZ(w2201), .A(w2246) );
	vdp_not g2152 (.nZ(w2211), .A(w2245) );
	vdp_not g2153 (.nZ(w2210), .A(w2244) );
	vdp_not g2154 (.nZ(w2200), .A(w2243) );
	vdp_nand g2155 (.Z(w2243), .A(w2224), .B(w2247) );
	vdp_sr_bit g2156 (.D(w2353), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2209) );
	vdp_sr_bit g2157 (.D(w2354), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2353) );
	vdp_sr_bit g2158 (.D(w2352), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2354) );
	vdp_sr_bit g2159 (.D(w2213), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2352) );
	vdp_sr_bit g2160 (.D(w2351), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2212) );
	vdp_sr_bit g2161 (.D(w2350), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2351) );
	vdp_sr_bit g2162 (.D(w2349), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2350) );
	vdp_sr_bit g2163 (.D(w2217), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2349) );
	vdp_sr_bit g2164 (.D(w2348), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2216) );
	vdp_sr_bit g2165 (.D(w2347), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2348) );
	vdp_sr_bit g2166 (.D(w2346), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2347) );
	vdp_sr_bit g2167 (.D(w2279), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2346) );
	vdp_sr_bit g2168 (.D(w2344), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2278) );
	vdp_sr_bit g2169 (.D(w2345), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2344) );
	vdp_sr_bit g2170 (.D(w2343), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2345) );
	vdp_sr_bit g2171 (.D(w2277), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2343) );
	vdp_sr_bit g2172 (.D(w2342), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2276) );
	vdp_sr_bit g2173 (.D(w2341), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2342) );
	vdp_sr_bit g2174 (.D(w2340), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2341) );
	vdp_sr_bit g2175 (.D(w2265), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2340) );
	vdp_sr_bit g2176 (.D(w2339), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2264) );
	vdp_sr_bit g2177 (.D(w2338), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2339) );
	vdp_sr_bit g2178 (.D(w2335), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2338) );
	vdp_sr_bit g2179 (.D(w2262), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2335) );
	vdp_sr_bit g2180 (.D(w2336), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2263) );
	vdp_sr_bit g2181 (.D(w2337), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2336) );
	vdp_sr_bit g2182 (.D(w2363), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2337) );
	vdp_sr_bit g2183 (.D(w2331), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2363) );
	vdp_sr_bit g2184 (.D(w2362), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2332) );
	vdp_sr_bit g2185 (.D(w2364), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2362) );
	vdp_sr_bit g2186 (.D(w2365), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2364) );
	vdp_sr_bit g2187 (.D(w2300), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2365) );
	vdp_sr_bit g2188 (.D(w2290), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2299) );
	vdp_sr_bit g2189 (.D(w2291), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2290) );
	vdp_sr_bit g2190 (.D(w2292), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2291) );
	vdp_sr_bit g2191 (.D(w2301), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2292) );
	vdp_sr_bit g2192 (.D(w2207), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2297) );
	vdp_sr_bit g2193 (.D(w2206), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2207) );
	vdp_sr_bit g2194 (.D(w2205), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2206) );
	vdp_sr_bit g2195 (.D(w2203), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2205) );
	vdp_aon2222 g2196 (.Z(w2075), .D2(1'b0), .C2(w2079), .C1(w2071), .D1(w2078), .B1(w2068), .A2(w2067), .A1(w2069), .B2(w2077) );
	vdp_cgi2a g2197 (.Z(w2417), .A(w2075), .C(w2429), .B(w2209) );
	vdp_aon2222 g2198 (.Z(w2076), .D2(1'b0), .C2(w2070), .C1(w2071), .D1(w2078), .B1(w2072), .A2(w2073), .A1(w2069), .B2(w2077) );
	vdp_cgi2a g2199 (.Z(w2429), .A(w2076), .C(w2428), .B(w2212) );
	vdp_aon2222 g2200 (.Z(w2323), .D2(1'b0), .C2(w2318), .C1(w2071), .D1(w2078), .B1(w2320), .A2(w2319), .A1(w2069), .B2(w2077) );
	vdp_cgi2a g2201 (.Z(w2428), .A(w2323), .C(w2427), .B(w2216) );
	vdp_aon2222 g2202 (.Z(w2322), .D2(w2400), .C2(w2423), .C1(w2071), .D1(w2078), .B1(w2424), .A2(w2425), .A1(w2069), .B2(w2077) );
	vdp_cgi2a g2203 (.Z(w2427), .A(w2322), .C(w2329), .B(w2278) );
	vdp_aon2222 g2204 (.Z(w2321), .D2(w2382), .C2(w2383), .C1(w2071), .D1(w2078), .B1(w2385), .A2(w2384), .A1(w2069), .B2(w2077) );
	vdp_cgi2a g2205 (.Z(w2329), .A(w2321), .C(w2330), .B(w2276) );
	vdp_aon2222 g2206 (.Z(w2393), .D2(w2328), .C2(w2420), .C1(w2071), .D1(w2078), .B1(w2421), .A2(w2422), .A1(w2069), .B2(w2077) );
	vdp_cgi2a g2207 (.Z(w2330), .A(w2393), .C(w2426), .B(w2264) );
	vdp_aon2222 g2208 (.Z(w2392), .D2(1'b0), .C2(w2386), .C1(w2071), .D1(w2078), .B1(w2387), .A2(w2388), .A1(w2069), .B2(w2077) );
	vdp_cgi2a g2209 (.Z(w2426), .A(w2392), .C(w2419), .B(w2263) );
	vdp_aon2222 g2210 (.Z(w2394), .D2(1'b0), .C2(w2389), .C1(w2071), .D1(w2078), .B1(w2390), .A2(w2391), .A1(w2069), .B2(w2077) );
	vdp_cgi2a g2211 (.Z(w2419), .A(w2394), .C(w2293), .B(w2332) );
	vdp_aon2222 g2212 (.Z(w2395), .D2(1'b0), .C2(w2401), .C1(w2071), .D1(w2078), .B1(w2402), .A2(w2403), .A1(w2069), .B2(w2077) );
	vdp_cgi2a g2213 (.Z(w2293), .A(w2395), .C(w2294), .B(w2299) );
	vdp_aon2222 g2214 (.Z(w2296), .D2(1'b0), .C2(w2399), .C1(w2071), .D1(w2078), .B1(w2397), .A2(w2398), .A1(w2069), .B2(w2077) );
	vdp_cgi2a g2215 (.Z(w2294), .A(w2296), .C(1'b1), .B(w2297) );
	vdp_not g2216 (.nZ(w2078), .A(w2396) );
	vdp_sr_bit g2217 (.D(w2377), .C1(w2201), .C2(w2200), .nC1(w2211), .nC2(w2210), .Q(w2298) );
	vdp_nand g2218 (.Z(w2396), .A(w2372), .B(w2298) );
	vdp_not g2219 (.nZ(w2071), .A(w2378) );
	vdp_sr_bit g2220 (.D(w2373), .Q(w2377), .C1(w2201), .C2(w2200), .nC1(w2211), .nC2(w2210) );
	vdp_nand g2221 (.Z(w2378), .A(w2372), .B(w2377) );
	vdp_not g2222 (.nZ(w2077), .A(w2376) );
	vdp_sr_bit g2223 (.D(w2309), .Q(w2373), .C1(w2201), .C2(w2200), .nC1(w2211), .nC2(w2210) );
	vdp_nand g2224 (.Z(w2376), .A(w2372), .B(w2373) );
	vdp_not g2225 (.nZ(w2069), .A(w2374) );
	vdp_sr_bit g2226 (.D(w2375), .Q(w2309), .C1(w2201), .C2(w2200), .nC1(w2211), .nC2(w2210) );
	vdp_nand g2227 (.Z(w2374), .A(w2372), .B(w2309) );
	vdp_sr_bit g2228 (.D(w2199), .Q(w2280), .C1(w2201), .C2(w2200), .nC1(w2211), .nC2(w2210) );
	vdp_sr_bit g2229 (.D(w2381), .Q(w2379), .C1(w2201), .C2(w2200), .nC1(w2211), .nC2(w2210) );
	vdp_sr_bit g2230 (.D(w2380), .Q(w2381), .C1(w2201), .C2(w2200), .nC1(w2211), .nC2(w2210) );
	vdp_sr_bit g2231 (.D(w2308), .Q(w2380), .C1(w2201), .C2(w2200), .nC1(w2211), .nC2(w2210) );
	vdp_sr_bit g2232 (.D(w2417), .Q(w2308), .C1(w2201), .C2(w2200), .nC1(w2211), .nC2(w2210) );
	vdp_not g2233 (.nZ(w2372), .A(w2280) );
	vdp_nor4 g2234 (.Z(w2375), .A(w2377), .B(w2373), .D(w2309), .C(w2199) );
	vdp_nor4 g2235 (.Z(w2270), .A(w2312), .B(w2313), .D(w2310), .C(w2311) );
	vdp_nor4 g2236 (.Z(w2272), .A(w2305), .B(w2306), .D(w2285), .C(w2286) );
	vdp_nor3 g2237 (.Z(w2271), .A(w2281), .B(w2282), .C(w2283) );
	vdp_not g2238 (.nZ(w2057), .A(w2280) );
	vdp_nand4 g2239 (.Z(w2269), .A(w2270), .B(w2272), .D(w2240), .C(w2271) );
	vdp_nand g2240 (.Z(w2274), .A(w2208), .B(w2273) );
	vdp_nand g2241 (.Z(w2275), .A(w2269), .B(w2274) );
	vdp_lfsr_bit g2242 (.Q(w2305), .A(w2275), .C2(w2200), .C1(w2201), .nC2(w2210), .nC1(w2211), .C(w2303), .B(w2304) );
	vdp_lfsr_bit g2243 (.Q(w2306), .A(w2305), .C2(w2200), .C1(w2201), .nC2(w2210), .nC1(w2211), .C(w2303), .B(w2304) );
	vdp_lfsr_bit g2244 (.Q(w2286), .A(w2306), .C2(w2200), .C1(w2201), .nC2(w2210), .nC1(w2211), .C(w2303), .B(w2304) );
	vdp_lfsr_bit g2245 (.Q(w2285), .A(w2286), .C2(w2200), .C1(w2201), .nC2(w2210), .nC1(w2211), .C(w2303), .B(w2304) );
	vdp_lfsr_bit g2246 (.Q(w2281), .A(w2285), .C2(w2200), .C1(w2201), .nC2(w2210), .nC1(w2211), .C(w2303), .B(w2304) );
	vdp_lfsr_bit g2247 (.Q(w2282), .A(w2281), .C2(w2200), .C1(w2201), .nC2(w2210), .nC1(w2211), .C(w2303), .B(w2304) );
	vdp_lfsr_bit g2248 (.Q(w2283), .A(w2282), .C2(w2200), .C1(w2201), .nC2(w2210), .nC1(w2211), .C(w2303), .B(w2304) );
	vdp_lfsr_bit g2249 (.Q(w2310), .A(w2283), .C2(w2200), .C1(w2201), .nC2(w2210), .nC1(w2211), .C(w2303), .B(w2304) );
	vdp_lfsr_bit g2250 (.Q(w2311), .A(w2310), .C2(w2200), .C1(w2201), .nC2(w2210), .nC1(w2211), .C(w2303), .B(w2304) );
	vdp_lfsr_bit g2251 (.Q(w2312), .A(w2311), .C2(w2200), .C1(w2201), .nC2(w2210), .nC1(w2211), .C(w2303), .B(w2304) );
	vdp_lfsr_bit g2252 (.Q(w2313), .A(w2312), .C2(w2200), .C1(w2201), .nC2(w2210), .nC1(w2211), .C(w2303), .B(w2304) );
	vdp_lfsr_bit g2253 (.Q(w2314), .A(w2313), .C2(w2200), .C1(w2201), .nC2(w2210), .nC1(w2211), .C(w2303), .B(w2304) );
	vdp_lfsr_bit g2254 (.Q(w2315), .A(w2314), .C2(w2200), .C1(w2201), .nC2(w2210), .nC1(w2211), .C(w2303), .B(w2304) );
	vdp_lfsr_bit g2255 (.Q(w2302), .A(w2315), .C2(w2201), .C1(w2201), .nC2(w2210), .nC1(w2211), .C(w2303), .B(w2304) );
	vdp_lfsr_bit g2256 (.Q(w2202), .A(w2302), .C2(w2200), .C1(w2201), .nC2(w2210), .nC1(w2211), .C(w2303), .B(w2304) );
	vdp_lfsr_bit g2257 (.Q(w2316), .A(w2202), .C2(w2200), .C1(w2201), .nC2(w2210), .nC1(w2211), .C(w2303), .B(w2304) );
	vdp_xor g2258 (.Z(w2208), .A(w2315), .B(w2316) );
	vdp_and g2259 (.Z(w2361), .A(w2204), .B(w2297) );
	vdp_ha g2260 (.SUM(w2203), .CO(w2259), .B(w2361), .A(1'b1) );
	vdp_and g2261 (.Z(w2334), .A(w2204), .B(w2299) );
	vdp_ha g2262 (.SUM(w2301), .CO(w2258), .B(w2334), .A(w2259) );
	vdp_and g2263 (.Z(w2333), .A(w2204), .B(w2332) );
	vdp_ha g2264 (.SUM(w2300), .CO(w2257), .B(w2333), .A(w2258) );
	vdp_and g2265 (.Z(w2261), .A(w2204), .B(w2263) );
	vdp_ha g2266 (.SUM(w2331), .CO(w2256), .B(w2261), .A(w2257) );
	vdp_and g2267 (.Z(w2360), .A(w2204), .B(w2264) );
	vdp_ha g2268 (.SUM(w2262), .CO(w2255), .B(w2360), .A(w2256) );
	vdp_and g2269 (.Z(w2359), .A(w2204), .B(w2276) );
	vdp_ha g2270 (.SUM(w2265), .CO(w2254), .B(w2359), .A(w2255) );
	vdp_and g2271 (.Z(w2358), .A(w2204), .B(w2278) );
	vdp_ha g2272 (.SUM(w2277), .CO(w2253), .B(w2358), .A(w2254) );
	vdp_and g2273 (.Z(w2357), .A(w2204), .B(w2216) );
	vdp_ha g2274 (.SUM(w2279), .CO(w2215), .B(w2357), .A(w2253) );
	vdp_and g2275 (.Z(w2356), .A(w2204), .B(w2212) );
	vdp_ha g2276 (.SUM(w2217), .CO(w2214), .B(w2356), .A(w2215) );
	vdp_and g2277 (.Z(w2355), .A(w2204), .B(w2209) );
	vdp_ha g2278 (.SUM(w2213), .B(w2355), .A(w2214) );
	vdp_and g2279 (.Z(w2284), .A(w2309), .B(w2379) );
	vdp_cnt_bit g2280 (.CI(w2284), .R(w2280), .C1(w2201), .nC1(w2211), .nC2(w2210), .C2(w2200), .Q(w2410) );
	vdp_and g2281 (.Z(w2288), .A(w2309), .B(w2381) );
	vdp_cnt_bit g2282 (.CI(w2288), .R(w2280), .C1(w2201), .nC1(w2211), .nC2(w2210), .C2(w2200), .Q(w2411) );
	vdp_and g2283 (.Z(w2287), .A(w2309), .B(w2380) );
	vdp_cnt_bit g2284 (.CI(w2287), .R(w2280), .C1(w2201), .nC1(w2211), .nC2(w2210), .C2(w2200), .Q(w2234) );
	vdp_and g2285 (.Z(w2307), .A(w2309), .B(w2308) );
	vdp_cnt_bit g2286 (.CI(w2307), .R(w2280), .C1(w2201), .nC1(w2211), .nC2(w2210), .C2(w2200), .Q(w2227) );
	vdp_nor g2287 (.Z(w2204), .A(w2417), .B(w2280) );
	vdp_dlatch g2288 (.Q(w2058), .C(w2055), .D(DB[7]), .nC(w2056) );
	vdp_comp_str g2289 (.A(w1065), .Z(w2055), .nZ(w2056) );
	vdp_and g2290 (.Z(w2050), .A(w2057), .B(w2058) );
	vdp_and g2291 (.Z(w2052), .A(w2051), .B(w2050) );
	vdp_and g2292 (.Z(w2436), .A(w2057), .B(w2435) );
	vdp_dlatch g2293 (.Q(w2435), .C(w2055), .D(DB[6]), .nC(w2056) );
	vdp_dlatch g2294 (.Q(w2178), .C(w2053), .D(w2436), .nC(w2054) );
	vdp_and g2295 (.Z(w2059), .A(w2057), .B(w2146) );
	vdp_dlatch g2296 (.Q(w2146), .C(w2055), .D(DB[5]), .nC(w2056) );
	vdp_dlatch g2297 (.Q(w2147), .C(w2053), .D(w2059), .nC(w2054) );
	vdp_and g2298 (.Z(w2062), .A(w2057), .B(w2145) );
	vdp_dlatch g2299 (.Q(w2145), .C(w2055), .D(DB[4]), .nC(w2056) );
	vdp_dlatch g2300 (.Q(w2177), .C(w2053), .D(w2062), .nC(w2054) );
	vdp_and g2301 (.Z(w2327), .A(w2057), .B(w2184) );
	vdp_dlatch g2302 (.Q(w2184), .C(w2055), .D(DB[3]), .nC(w2056) );
	vdp_or g2303 (.Z(w2170), .A(w2185), .B(w2327) );
	vdp_and g2304 (.Z(w2325), .A(w2057), .B(w2434) );
	vdp_or g2305 (.Z(w2158), .A(w2185), .B(w2325) );
	vdp_dlatch g2306 (.Q(w2434), .C(w2055), .D(DB[2]), .nC(w2056) );
	vdp_not g2307 (.nZ(w2185), .A(w2057) );
	vdp_and g2308 (.Z(w2324), .A(w2057), .B(w2326) );
	vdp_or g2309 (.Z(w2156), .A(w2185), .B(w2324) );
	vdp_dlatch g2310 (.Q(w2326), .C(w2055), .D(DB[1]), .nC(w2056) );
	vdp_and g2311 (.Z(w2190), .A(w2057), .B(w2191) );
	vdp_or g2312 (.Z(w2159), .A(w2185), .B(w2190) );
	vdp_dlatch g2313 (.Q(w2191), .C(w2055), .D(DB[0]), .nC(w2056) );
	vdp_not g2314 (.nZ(w2189), .A(w2187) );
	vdp_aoi21 g2315 (.Z(w2187), .B(w2199), .A1(w2192), .A2(w2186) );
	vdp_and3 g2316 (.Z(w2186), .A(w2167), .B(w2166), .C(w2177) );
	vdp_not g2317 (.nZ(w2188), .A(w2432) );
	vdp_aoi21 g2318 (.Z(w2432), .B(w2199), .A1(w2192), .A2(w2433) );
	vdp_and3 g2319 (.Z(w2433), .A(w2167), .B(w2147), .C(w2177) );
	vdp_not g2320 (.nZ(w2450), .A(w2431) );
	vdp_aoi21 g2321 (.Z(w2431), .B(w2199), .A1(w2192), .A2(w2430) );
	vdp_and3 g2322 (.Z(w2430), .A(w2178), .B(w2166), .C(w2168) );
	vdp_not g2323 (.nZ(w2196), .A(w2050) );
	vdp_or g2324 (.Z(w2198), .A(w2050), .B(w2199) );
	vdp_and g2325 (.Z(w2437), .A(w2198), .B(w2450) );
	vdp_and g2326 (.Z(w2317), .A(w2196), .B(w2450) );
	vdp_and g2327 (.Z(w2408), .A(w2198), .B(w2183) );
	vdp_and g2328 (.Z(w2438), .A(w2196), .B(w2183) );
	vdp_not g2329 (.nZ(w2183), .A(w2182) );
	vdp_aoi21 g2330 (.Z(w2182), .B(w2199), .A1(w2192), .A2(w2181) );
	vdp_and3 g2331 (.Z(w2181), .A(w2167), .B(w2147), .C(w2168) );
	vdp_not g2332 (.nZ(w2179), .A(w2180) );
	vdp_aoi21 g2333 (.Z(w2180), .B(w2199), .A1(w2192), .A2(w2194) );
	vdp_and3 g2334 (.Z(w2194), .A(w2178), .B(w2166), .C(w2177) );
	vdp_and g2335 (.Z(w2197), .A(w2198), .B(w2193) );
	vdp_and g2336 (.Z(w2195), .A(w2196), .B(w2193) );
	vdp_not g2337 (.nZ(w2193), .A(w2176) );
	vdp_aoi21 g2338 (.Z(w2176), .B(w2199), .A1(w2192), .A2(w2175) );
	vdp_and3 g2339 (.Z(w2175), .A(w2167), .B(w2166), .C(w2168) );
	vdp_and3 g2340 (.Z(w2174), .A(w2178), .B(w2147), .C(w2177) );
	vdp_not g2341 (.nZ(w2162), .A(w2173) );
	vdp_aoi21 g2342 (.Z(w2173), .B(w2199), .A1(w2192), .A2(w2174) );
	vdp_and3 g2343 (.Z(w2171), .A(w2178), .B(w2147), .C(w2168) );
	vdp_not g2344 (.nZ(w2226), .A(w2172) );
	vdp_aoi21 g2345 (.Z(w2172), .B(w2199), .A1(w2192), .A2(w2171) );
	vdp_not g2346 (.nZ(w2413), .A(w2416) );
	vdp_not g2347 (.nZ(w2414), .A(w2415) );
	vdp_not g2348 (.nZ(w2168), .A(w2177) );
	vdp_not g2349 (.nZ(w2166), .A(w2147) );
	vdp_not g2350 (.nZ(w2167), .A(w2178) );
	vdp_nor g2351 (.Z(w2042), .A(w2410), .B(w1162) );
	vdp_nor g2352 (.Z(w2144), .A(w2411), .B(w1162) );
	vdp_nor g2353 (.Z(w2157), .A(w2234), .B(w1162) );
	vdp_nor g2354 (.Z(w2164), .A(w2202), .B(w1162) );
	vdp_aon22 g2355 (.Z(w2229), .A2(w2234), .A1(w2233), .B2(w2228), .B1(w2227) );
	vdp_sr_bit g2356 (.D(w2229), .nC1(w2211), .nC2(w2210), .C1(w2201), .C2(w2200), .Q(w2230) );
	vdp_not g2357 (.nZ(w2228), .A(w2233) );
	vdp_not g2358 (.nZ(w2231), .A(w2230) );
	vdp_not g2359 (.nZ(w2367), .A(w1163) );
	vdp_not g2360 (.nZ(w2366), .A(w1164) );
	vdp_not g2361 (.nZ(w2267), .A(w2266) );
	vdp_sr_bit g2362 (.D(w2051), .nC1(w2220), .nC2(w2222), .C1(w2219), .C2(w2221), .Q(w2192) );
	vdp_nand g2363 (.Z(w2368), .A(w1163), .B(w2366) );
	vdp_nand g2364 (.Z(w2232), .A(w1164), .B(w1163) );
	vdp_nand g2365 (.Z(w2369), .A(w2366), .B(w2367) );
	vdp_nand g2366 (.Z(w2370), .A(w1164), .B(w2367) );
	vdp_and g2367 (.Z(w2236), .A(w2229), .B(w2231) );
	vdp_and g2368 (.Z(w2015), .A(w1162), .B(w2232) );
	vdp_and g2369 (.Z(w2016), .A(w1162), .B(w2368) );
	vdp_and g2370 (.Z(w2017), .A(w1162), .B(w2369) );
	vdp_and g2371 (.Z(w2018), .A(w1162), .B(w2370) );
	vdp_nor4 g2372 (.Z(w2240), .A(w2302), .B(w2315), .D(w2314), .C(w2202) );
	vdp_not g2373 (.nZ(w2237), .A(w2236) );
	vdp_not g2374 (.nZ(w2304), .A(w2238) );
	vdp_not g2375 (.nZ(w2303), .A(w2371) );
	vdp_not g2376 (.nZ(w2199), .A(w2267) );
	vdp_nand g2377 (.Z(w2238), .A(w2235), .B(w2237) );
	vdp_nand g2378 (.Z(w2371), .A(w2235), .B(w2236) );
	vdp_nor g2379 (.Z(w2235), .A(w2199), .B(w2239) );
	vdp_rs_ff g2380 (.S(w2226), .R(w2239), .Q(w2268) );
	vdp_rs_ff g2381 (.S(w2051), .R(w1065), .Q(w2241) );
	vdp_nor g2382 (.Z(w2242), .A(w1065), .B(w2241) );
	vdp_comp_dff g2383 (.D(w2242), .nC1(w2220), .C1(w2219), .C2(w2221), .nC2(w2222), .Q(w2051) );
	vdp_comp_dff g2384 (.D(SYSRES), .nC1(w2211), .C1(w2201), .C2(w2200), .nC2(w2210), .Q(w2266) );
	vdp_comp_dff g2385 (.D(w2268), .nC1(w2211), .C1(w2201), .C2(w2200), .nC2(w2210), .Q(w2239) );
	vdp_sr_bit g2386 (.Q(w2623), .D(w2617), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2387 (.nZ(AD_RD_DIR), .A(w2616) );
	vdp_sr_bit g2388 (.Q(w2624), .D(w2485), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2389 (.Q(w2551), .D(w2498), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2390 (.Q(w2607), .D(w33), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2391 (.Q(w2477), .D(w35), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2392 (.nZ(w2619), .A(w2475) );
	vdp_or g2393 (.Z(w2485), .A(w35), .B(w2477) );
	vdp_sr_bit g2394 (.Q(w2494), .D(w2496), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_sr_bit g2395 (.Q(w2620), .D(w2609), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2396 (.nZ(w2550), .A(w2620) );
	vdp_or g2397 (.Z(w2473), .A(w2477), .B(w2476) );
	vdp_sr_bit g2398 (.Q(w2476), .D(w555), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2399 (.Q(w2474), .D(w32), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2400 (.Q(w2611), .D(w2474), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2401 (.Q(w2610), .D(w2486), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2402 (.Q(w2605), .D(w2607), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_sr_bit g2403 (.Q(w2622), .D(w2627), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_not g2404 (.nZ(w2601), .A(w2682) );
	vdp_not g2405 (.nZ(w2497), .A(128k) );
	vdp_sr_bit g2406 (.Q(w2486), .D(VRAM_REFRESH), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2407 (.nZ(w2558), .A(w2472) );
	vdp_not g2408 (.nZ(w2625), .A(w2612) );
	vdp_not g2409 (.nZ(w2492), .A(w2484) );
	vdp_oai21 g2410 (.Z(w2472), .B(w2492), .A1(w2625), .A2(w2613) );
	vdp_or g2411 (.Z(w2484), .A(w2619), .B(w2618) );
	vdp_or g2412 (.Z(w2617), .A(w2476), .B(w555) );
	vdp_not g2413 (.nZ(w2626), .A(w2478) );
	vdp_not g2414 (.nZ(w2674), .A(w2627) );
	vdp_dlatch_inv g2415 (.nQ(w2627), .D(w3), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2416 (.nQ(w2621), .D(w2493), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g2417 (.nQ(w2493), .D(w2622), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g2418 (.nQ(w2475), .D(w2473), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2419 (.nQ(w2618), .D(w2475), .C(HCLK2), .nC(nHCLK2) );
	vdp_dlatch_inv g2420 (.nQ(w2615), .D(w2614), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2421 (.nQ(w2612), .D(w2611), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g2422 (.nQ(w2613), .D(w2612), .C(HCLK2), .nC(nHCLK2) );
	vdp_aon22 g2423 (.Z(nCAS1), .A1(w2493), .B1(w2482), .B2(1'b1), .A2(w2620) );
	vdp_and3 g2424 (.Z(nWE1), .A(w2481), .B(w2624), .C(w2482) );
	vdp_and3 g2425 (.Z(nWE0), .A(w2482), .B(w2481), .C(w2623) );
	vdp_aoi222 g2426 (.Z(w2616), .A1(1'b1), .B1(w2479), .B2(1'b1), .A2(w100), .C1(w2484), .C2(w2482) );
	vdp_aon333 g2427 (.Z(nOE1), .A1(w2558), .A2(w2622), .A3(w2482), .B1(w2615), .B2(w2615), .B3(w2626), .C1(w2615), .C2(w2615), .C3(w2479) );
	vdp_or3 g2428 (.Z(w2614), .A(w2609), .B(w2611), .C(w2474) );
	vdp_sr_bit g2429 (.Q(w2479), .D(w2674), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_dlatch_inv g2430 (.nQ(w2481), .D(w2479), .C(DCLK1), .nC(nDCLK1) );
	vdp_dlatch_inv g2431 (.nQ(w2608), .D(w2481), .C(DCLK2), .nC(nDCLK2) );
	vdp_dlatch_inv g2432 (.nQ(w2482), .D(w2480), .C(DCLK1), .nC(nDCLK1) );
	vdp_not g2433 (.nZ(w2480), .A(w2608) );
	vdp_nand g2434 (.Z(w2702), .A(w2608), .B(w2479) );
	vdp_nand g2435 (.Z(w2701), .A(w2479), .B(w2621) );
	vdp_nand g2436 (.Z(w2488), .A(w2622), .B(1'b1) );
	vdp_aoi33 g2437 (.Z(w2688), .A1(w2605), .A2(w34), .A3(w34), .B1(w2499), .B2(w2500), .B3(w3) );
	vdp_and g2438 (.Z(w2495), .A(w2482), .B(w2481) );
	vdp_not g2439 (.nZ(w2489), .A(w2551) );
	vdp_comp_strong g2440 (.nZ(w2506), .Z(w2505), .A(w2512) );
	vdp_comp_strong g2441 (.nZ(w2573), .Z(w2596), .A(w2597) );
	vdp_comp_strong g2442 (.nZ(w2507), .Z(w2552), .A(w2597) );
	vdp_comp_strong g2443 (.nZ(w2556), .Z(w2555), .A(w2512) );
	vdp_comp_strong g2444 (.nZ(w2513), .Z(w2557), .A(w2509) );
	vdp_comp_strong g2445 (.nZ(w2560), .Z(w2602), .A(w2509) );
	vdp_not g2446 (.nZ(w2515), .A(w2479) );
	vdp_not g2447 (.nZ(w2500), .A(w34) );
	vdp_not g2448 (.nZ(w2499), .A(w36) );
	vdp_comp_strong g2449 (.nZ(w2554), .Z(w6817), .A(w2495) );
	vdp_comp_strong g2450 (.nZ(w2490), .Z(w2598), .A(w2495) );
	vdp_or g2451 (.Z(w2609), .A(w2486), .B(w2610) );
	vdp_and g2452 (.Z(w2496), .A(128k), .B(HCLK1) );
	vdp_comp_we g2453 (.nZ(w2599), .Z(w2600), .A(w100) );
	vdp_comp_we g2454 (.nZ(w2508), .Z(w2686), .A(w2516) );
	vdp_not g2455 (.nZ(w2687), .A(w2551) );
	vdp_not g2456 (.nZ(w2511), .A(w2702) );
	vdp_not g2457 (.nZ(w6822), .A(w2701) );
	vdp_not g2458 (.nZ(w6823), .A(w2488) );
	vdp_comp_we g2459 (.nZ(w6824), .Z(w2604), .A(M5) );
	vdp_comp_we g2460 (.nZ(w2559), .Z(w2514), .A(128k) );
	vdp_and g2461 (.Z(w2498), .A(w110), .B(w3) );
	vdp_and g2462 (.Z(w2509), .A(w3), .B(HCLK1) );
	vdp_and g2463 (.Z(w2512), .A(HCLK2), .B(w2606) );
	vdp_and g2464 (.Z(w2597), .A(w3), .B(HCLK1) );
	vdp_oai21 g2465 (.Z(w2682), .A1(HCLK2), .A2(w2497), .B(DCLK1) );
	vdp_notif0 g2466 (.nZ(AD_DATA[0]), .A(w2503), .nE(w2489) );
	vdp_aon22 g2467 (.Z(nYS), .A1(VRAMA[16]), .A2(w2600), .B1(w2599), .B2(w2666) );
	vdp_aon22 g2468 (.Z(w2642), .A1(VRAMA[15]), .B1(w2599), .A2(w2600), .B2(w2580) );
	vdp_aon22 g2469 (.Z(w2640), .A1(VRAMA[14]), .B1(w2599), .A2(w2600), .B2(w2463) );
	vdp_aon22 g2470 (.Z(w2462), .A1(VRAMA[6]), .B1(w2599), .A2(w2600), .B2(w2641) );
	vdp_aon22 g2471 (.Z(w2454), .A1(VRAMA[7]), .B1(w2599), .A2(w2600), .B2(w2453) );
	vdp_aon22 g2472 (.Z(w2670), .A1(VRAMA[13]), .B1(w2599), .A2(w2600), .B2(w2471) );
	vdp_aon22 g2473 (.Z(w2639), .A1(VRAMA[5]), .B1(w2599), .A2(w2600), .B2(w2690) );
	vdp_aon22 g2474 (.Z(w2645), .A1(VRAMA[12]), .B1(w2599), .A2(w2600), .B2(w2540) );
	vdp_aon22 g2475 (.Z(w2469), .A1(VRAMA[4]), .B1(w2599), .A2(w2600), .B2(w2547) );
	vdp_aon22 g2476 (.Z(w2644), .A1(VRAMA[11]), .B1(w2599), .A2(w2600), .B2(w2695) );
	vdp_aon22 g2477 (.Z(w2579), .A1(VRAMA[3]), .B1(w2599), .A2(w2600), .B2(w2691) );
	vdp_aon22 g2478 (.Z(w2672), .A1(VRAMA[10]), .B1(w2599), .A2(w2600), .B2(w2592) );
	vdp_aon22 g2479 (.Z(w2578), .A1(VRAMA[2]), .B1(w2599), .A2(w2600), .B2(w2536) );
	vdp_aon22 g2480 (.Z(w2501), .A1(VRAMA[8]), .B1(w2599), .A2(w2600), .B2(w2504) );
	vdp_aon22 g2481 (.Z(w2693), .A1(VRAMA[0]), .B1(w2599), .A2(w2600), .B2(w2527) );
	vdp_aon22 g2482 (.Z(w2694), .A1(VRAMA[9]), .B1(w2599), .A2(w2600), .B2(w2574) );
	vdp_aon22 g2483 (.Z(w2530), .A1(VRAMA[1]), .B1(w2599), .A2(w2600), .B2(w2532) );
	vdp_notif0 g2484 (.nZ(AD_DATA[1]), .A(w2522), .nE(w2489) );
	vdp_notif0 g2485 (.nZ(AD_DATA[2]), .A(w2576), .nE(w2489) );
	vdp_notif0 g2486 (.nZ(AD_DATA[3]), .A(w2533), .nE(w2489) );
	vdp_notif0 g2487 (.nZ(AD_DATA[5]), .A(w2470), .nE(w2489) );
	vdp_notif0 g2488 (.nZ(AD_DATA[4]), .A(w2553), .nE(w2489) );
	vdp_notif0 g2489 (.nZ(AD_DATA[6]), .A(w2464), .nE(w2489) );
	vdp_notif0 g2490 (.nZ(AD_DATA[7]), .A(w2461), .nE(w2489) );
	vdp_slatch g2491 (.nQ(w2503), .D(w2502), .nC(w2490), .C(w2598) );
	vdp_slatch g2492 (.nQ(w2522), .D(w2521), .nC(w2490), .C(w2598) );
	vdp_slatch g2493 (.nQ(w2576), .D(w2529), .nC(w2490), .C(w2598) );
	vdp_slatch g2494 (.nQ(w2533), .D(w2534), .nC(w2490), .C(w2598) );
	vdp_slatch g2495 (.nQ(w2553), .D(w2487), .nC(w2490), .C(w2598) );
	vdp_slatch g2496 (.nQ(w2470), .D(w2671), .nC(w2490), .C(w2598) );
	vdp_slatch g2497 (.nQ(w2464), .D(w2542), .nC(w2490), .C(w2598) );
	vdp_slatch g2498 (.nQ(w2461), .D(w2643), .nC(w2490), .C(w2598) );
	vdp_slatch g2499 (.nQ(w2456), .D(w2455), .nC(w2554), .C(w6817) );
	vdp_slatch g2500 (.nQ(w2545), .D(w2541), .nC(w2554), .C(w6817) );
	vdp_slatch g2501 (.nQ(w2583), .D(w2683), .nC(w2554), .C(w6817) );
	vdp_slatch g2502 (.nQ(w2584), .D(w2468), .nC(w2554), .C(w6817) );
	vdp_slatch g2503 (.nQ(w2646), .D(w2543), .nC(w2554), .C(w6817) );
	vdp_slatch g2504 (.nQ(w2537), .D(w2535), .nC(w2554), .C(w6817) );
	vdp_slatch g2505 (.nQ(w2531), .D(w2577), .nC(w2554), .C(w6817) );
	vdp_slatch g2506 (.nQ(w2561), .D(w2673), .nC(w2554), .C(w6817) );
	vdp_slatch g2507 (.Q(w2504), .D(w2564), .nC(w2506), .C(w2505) );
	vdp_slatch g2508 (.Q(w2574), .D(w2697), .nC(w2506), .C(w2505) );
	vdp_slatch g2509 (.Q(w2695), .D(w2649), .nC(w2506), .C(w2505) );
	vdp_slatch g2510 (.Q(w2592), .D(w2575), .nC(w2506), .C(w2505) );
	vdp_slatch g2511 (.Q(w2471), .D(w2563), .nC(w2506), .C(w2505) );
	vdp_slatch g2512 (.Q(w2540), .D(w2650), .nC(w2506), .C(w2505) );
	vdp_slatch g2513 (.Q(w2580), .D(w2653), .nC(w2506), .C(w2505) );
	vdp_slatch g2514 (.Q(w2463), .D(w2562), .nC(w2506), .C(w2505) );
	vdp_slatch g2515 (.nQ(w2652), .D(w358), .nC(w2573), .C(w2596) );
	vdp_slatch g2516 (.nQ(w2654), .D(RD_DATA[6]), .nC(w2573), .C(w2596) );
	vdp_slatch g2517 (.nQ(w2651), .D(RD_DATA[5]), .nC(w2573), .C(w2596) );
	vdp_slatch g2518 (.nQ(w2699), .D(RD_DATA[4]), .nC(w2573), .C(w2596) );
	vdp_slatch g2519 (.nQ(w2648), .D(w324), .nC(w2573), .C(w2596) );
	vdp_slatch g2520 (.nQ(w2700), .D(RD_DATA[2]), .nC(w2573), .C(w2596) );
	vdp_slatch g2521 (.nQ(w2698), .D(RD_DATA[0]), .nC(w2573), .C(w2596) );
	vdp_slatch g2522 (.nQ(w2647), .D(RD_DATA[1]), .nC(w2573), .C(w2596) );
	vdp_notif0 g2523 (.nZ(w358), .A(w2456), .nE(w2687) );
	vdp_notif0 g2524 (.nZ(RD_DATA[6]), .A(w2545), .nE(w2687) );
	vdp_notif0 g2525 (.nZ(RD_DATA[5]), .A(w2583), .nE(w2687) );
	vdp_notif0 g2526 (.nZ(RD_DATA[4]), .A(w2584), .nE(w2687) );
	vdp_notif0 g2527 (.nZ(w324), .A(w2646), .nE(w2687) );
	vdp_notif0 g2528 (.nZ(RD_DATA[2]), .A(w2537), .nE(w2687) );
	vdp_notif0 g2529 (.nZ(RD_DATA[1]), .A(w2531), .nE(w2687) );
	vdp_notif0 g2530 (.nZ(RD_DATA[0]), .A(w2561), .nE(w2687) );
	vdp_slatch g2531 (.nQ(w2676), .D(AD_DATA[7]), .nC(w2507), .C(w2552) );
	vdp_slatch g2532 (.nQ(w2675), .D(AD_DATA[6]), .nC(w2507), .C(w2552) );
	vdp_slatch g2533 (.nQ(w2696), .D(AD_DATA[5]), .nC(w2507), .C(w2552) );
	vdp_slatch g2534 (.nQ(w2678), .D(AD_DATA[3]), .nC(w2507), .C(w2552) );
	vdp_slatch g2535 (.nQ(w2679), .D(AD_DATA[2]), .nC(w2507), .C(w2552) );
	vdp_slatch g2536 (.nQ(w2681), .D(AD_DATA[1]), .nC(w2507), .C(w2552) );
	vdp_slatch g2537 (.nQ(w2680), .D(AD_DATA[0]), .nC(w2507), .C(w2552) );
	vdp_slatch g2538 (.Q(w2460), .D(w2572), .nC(w2556), .C(w2555) );
	vdp_slatch g2539 (.Q(w2467), .D(w2571), .nC(w2556), .C(w2555) );
	vdp_slatch g2540 (.Q(w2544), .D(w2570), .nC(w2556), .C(w2555) );
	vdp_slatch g2541 (.Q(w2684), .D(w2567), .nC(w2556), .C(w2555) );
	vdp_slatch g2542 (.Q(w2595), .D(w2568), .nC(w2556), .C(w2555) );
	vdp_slatch g2543 (.Q(w2528), .D(w2566), .nC(w2556), .C(w2555) );
	vdp_slatch g2544 (.Q(w2582), .D(w2459), .nC(w2513), .C(w2557) );
	vdp_slatch g2545 (.Q(w2689), .D(w2466), .nC(w2513), .C(w2557) );
	vdp_slatch g2546 (.Q(w2656), .D(w2520), .nC(w2513), .C(w2557) );
	vdp_slatch g2547 (.Q(w2586), .D(w2519), .nC(w2513), .C(w2557) );
	vdp_slatch g2548 (.Q(w2593), .D(w2594), .nC(w2513), .C(w2557) );
	vdp_slatch g2549 (.Q(w2685), .D(w2525), .nC(w2513), .C(w2557) );
	vdp_slatch g2550 (.Q(w2591), .D(w2491), .nC(w2513), .C(w2557) );
	vdp_slatch g2551 (.Q(w2692), .D(w2526), .nC(w2513), .C(w2557) );
	vdp_slatch g2552 (.Q(w2603), .D(w2524), .nC(w2560), .C(w2602) );
	vdp_slatch g2553 (.Q(w2590), .D(w2707), .nC(w2560), .C(w2602) );
	vdp_slatch g2554 (.Q(w2538), .D(w2518), .nC(w2560), .C(w2602) );
	vdp_slatch g2555 (.Q(w2587), .D(w2703), .nC(w2560), .C(w2602) );
	vdp_slatch g2556 (.Q(w2548), .D(w2465), .nC(w2560), .C(w2602) );
	vdp_slatch g2557 (.Q(w2585), .D(w2517), .nC(w2560), .C(w2602) );
	vdp_slatch g2558 (.Q(w2546), .D(w2458), .nC(w2560), .C(w2602) );
	vdp_slatch g2559 (.Q(w2581), .D(w2457), .nC(w2560), .C(w2602) );
	vdp_sr_bit g2560 (.Q(w2516), .D(w34), .C2(HCLK2), .C1(HCLK1), .nC1(nHCLK1), .nC2(nHCLK2) );
	vdp_not g2561 (.nZ(w2714), .A(w111) );
	vdp_not g2562 (.nZ(w2588), .A(w2589) );
	vdp_not g2563 (.nZ(w6825), .A(M5) );
	vdp_not g2564 (.nZ(w2523), .A(w2515) );
	vdp_not g2565 (.nZ(w2478), .A(w2523) );
	vdp_aoi21 g2566 (.Z(w2589), .B(w2657), .A2(VRAMA[9]), .A1(w6825) );
	vdp_aoi22 g2567 (.Z(w2697), .A1(w2531), .B1(w2508), .B2(w2647), .A2(w2686) );
	vdp_aoi22 g2568 (.Z(w2649), .A1(w2646), .B1(w2508), .B2(w2648), .A2(w2686) );
	vdp_aoi22 g2569 (.Z(w2575), .A1(w2537), .B1(w2508), .B2(w2700), .A2(w2686) );
	vdp_aoi22 g2570 (.Z(w2563), .A1(w2583), .B1(w2508), .B2(w2651), .A2(w2686) );
	vdp_aoi22 g2571 (.Z(w2650), .A1(w2584), .B1(w2508), .B2(w2699), .A2(w2686) );
	vdp_aoi22 g2572 (.Z(w2653), .A1(w2456), .B1(w2508), .B2(w2652), .A2(w2686) );
	vdp_aoi22 g2573 (.Z(w2562), .A1(w2545), .B1(w2508), .B2(w2654), .A2(w2686) );
	vdp_slatch g2574 (.Q(w2510), .D(w2565), .nC(w2556), .C(w2555) );
	vdp_slatch g2575 (.nQ(w2677), .D(AD_DATA[4]), .nC(w2507), .C(w2552) );
	vdp_slatch g2576 (.Q(w2539), .D(w2569), .nC(w2556), .C(w2555) );
	vdp_aoi22 g2577 (.Z(w2565), .A1(w2503), .B1(w2508), .B2(w2680), .A2(w2686) );
	vdp_aoi22 g2578 (.Z(w2566), .A1(w2522), .B1(w2508), .B2(w2681), .A2(w2686) );
	vdp_aoi22 g2579 (.Z(w2567), .A1(w2576), .B1(w2508), .B2(w2679), .A2(w2686) );
	vdp_aoi22 g2580 (.Z(w2568), .A1(w2533), .B1(w2508), .B2(w2678), .A2(w2686) );
	vdp_aoi22 g2581 (.Z(w2569), .A1(w2553), .B1(w2508), .B2(w2677), .A2(w2686) );
	vdp_aoi22 g2582 (.Z(w2570), .A1(w2470), .B1(w2508), .B2(w2696), .A2(w2686) );
	vdp_aoi22 g2583 (.Z(w2572), .A1(w2461), .B1(w2508), .B2(w2676), .A2(w2686) );
	vdp_aoi22 g2584 (.Z(w2571), .A1(w2464), .B1(w2508), .B2(w2675), .A2(w2686) );
	vdp_aon22 g2585 (.Z(w2526), .A1(VRAMA[2]), .B1(w6824), .B2(VRAMA[1]), .A2(w2604) );
	vdp_aon22 g2586 (.Z(w2525), .A1(VRAMA[3]), .B1(w6824), .B2(VRAMA[2]), .A2(w2604) );
	vdp_aon22 g2587 (.Z(w2491), .A1(VRAMA[4]), .B1(w6824), .B2(VRAMA[3]), .A2(w2604) );
	vdp_aon22 g2588 (.Z(w2594), .A1(VRAMA[5]), .B1(w6824), .B2(VRAMA[4]), .A2(w2604) );
	vdp_aon22 g2589 (.Z(w2519), .A1(VRAMA[6]), .B1(w6824), .B2(VRAMA[5]), .A2(w2604) );
	vdp_aon22 g2590 (.Z(w2520), .A1(VRAMA[7]), .B1(w6824), .B2(VRAMA[6]), .A2(w2604) );
	vdp_aon22 g2591 (.Z(w2466), .A1(VRAMA[8]), .B1(w6824), .B2(VRAMA[7]), .A2(w2604) );
	vdp_aon22 g2592 (.Z(w2459), .A1(VRAMA[9]), .B1(w6824), .B2(VRAMA[8]), .A2(w2604) );
	vdp_and g2593 (.Z(w2657), .A(VRAMA[1]), .B(M5) );
	vdp_aon22 g2594 (.Z(w2457), .A1(w2655), .B1(w2559), .B2(VRAMA[15]), .A2(w2514) );
	vdp_aon22 g2595 (.Z(w2458), .A1(VRAMA[15]), .B1(w2559), .B2(VRAMA[14]), .A2(w2514) );
	vdp_aon22 g2596 (.Z(w2465), .A1(VRAMA[14]), .B1(w2559), .B2(VRAMA[13]), .A2(w2514) );
	vdp_aon22 g2597 (.Z(w2703), .A1(VRAMA[12]), .B1(w2559), .B2(VRAMA[11]), .A2(w2514) );
	vdp_aon22 g2598 (.Z(w2517), .A1(VRAMA[13]), .B1(w2559), .B2(VRAMA[12]), .A2(w2514) );
	vdp_aon22 g2599 (.Z(w2518), .A1(VRAMA[11]), .B1(w2559), .B2(VRAMA[10]), .A2(w2514) );
	vdp_aon22 g2600 (.Z(w2707), .A1(VRAMA[10]), .B1(w2559), .B2(w2588), .A2(w2514) );
	vdp_aon22 g2601 (.Z(w2524), .A1(w2657), .B1(w2559), .B2(VRAMA[0]), .A2(w2514) );
	vdp_aon22 g2602 (.Z(w2655), .A1(w2714), .B1(w111), .B2(w94), .A2(VRAMA[16]) );
	vdp_aon222 g2603 (.Z(w2527), .A1(w2511), .A2(w2510), .B1(w6822), .B2(w2692), .C1(w6823), .C2(w2603) );
	vdp_aon222 g2604 (.Z(w2532), .A1(w2511), .A2(w2528), .B1(w6822), .B2(w2685), .C1(w6823), .C2(w2590) );
	vdp_aon222 g2605 (.Z(w2536), .A1(w2511), .A2(w2684), .B1(w6822), .B2(w2591), .C1(w6823), .C2(w2538) );
	vdp_aon222 g2606 (.Z(w2691), .A1(w2511), .A2(w2595), .B1(w6822), .B2(w2593), .C1(w6823), .C2(w2587) );
	vdp_aon222 g2607 (.Z(w2547), .A1(w2511), .A2(w2539), .B1(w6822), .B2(w2586), .C1(w6823), .C2(w2585) );
	vdp_aon222 g2608 (.Z(w2690), .A1(w2511), .A2(w2544), .B1(w6822), .B2(w2656), .C1(w6823), .C2(w2548) );
	vdp_aon222 g2609 (.Z(w2641), .A1(w2511), .A2(w2467), .B1(w6822), .B2(w2689), .C1(w6823), .C2(w2546) );
	vdp_aon222 g2610 (.Z(w2453), .A1(w2511), .A2(w2460), .B1(w6822), .B2(w2582), .C1(w6823), .C2(w2581) );
	vdp_dlatch_inv g2611 (.nQ(w2606), .D(w2688), .C(HCLK1), .nC(nHCLK1) );
	vdp_comp_we g2612 (.Z(w2549), .A(w2608) );
	vdp_aon22 g2613 (.Z(nRAS1), .A1(1'b1), .B1(w2550), .B2(w2493), .A2(w2549) );
	vdp_aoi22 g2614 (.Z(w2564), .A1(w2561), .B1(w2508), .B2(w2698), .A2(w2686) );
	vdp_and g2615 (.Z(w2628), .B(w2712), .A(DCLK2) );
	vdp_nor g2616 (.Z(w2708), .A(w2630), .B(RES) );
	vdp_sr_bit g2617 (.Q(w2630), .D(w2708), .C2(DCLK2), .C1(DCLK1), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_dlatch_inv g2618 (.nQ(w2709), .D(w2631), .C(DCLK1), .nC(nDCLK1) );
	vdp_and g2619 (.Z(w2710), .A(DCLK2), .B(w2709) );
	vdp_dlatch_inv g2620 (.nQ(w2712), .D(w2630), .C(DCLK1), .nC(nDCLK1) );
	vdp_not g2621 (.nZ(w2634), .A(w2636) );
	vdp_not g2622 (.nZ(w2633), .A(w2711) );
	vdp_neg_dff g2623 (.Q(w2636), .C(DCLK1), .D(1'b1), .R(w2628) );
	vdp_not g2624 (.A(w2630), .nZ(w2631) );
	vdp_neg_dff g2625 (.Q(w2711), .R(w2710), .C(DCLK1), .D(1'b1) );
	vdp_sr_bit g2626 (.Q(w2790), .D(w2782), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2627 (.Q(w2786), .D(w2785), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2628 (.Q(w2980), .D(w2786), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2629 (.Q(w2803), .D(w2980), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2630 (.Q(w2758), .D(RD_DATA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2631 (.Q(w2759), .D(RD_DATA[2]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2632 (.Q(w2760), .D(w324), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2633 (.Q(w2961), .D(w2983), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2634 (.Q(w2983), .D(w2984), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2635 (.Q(w2984), .D(w2985), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2636 (.Q(w2985), .D(w2986), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2637 (.Q(w2986), .D(w2987), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2638 (.Q(w2987), .D(w2988), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2639 (.Q(w2988), .D(w2989), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2640 (.Q(w2989), .D(w18), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2641 (.Q(w2768), .D(w2761), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2642 (.Q(w2766), .D(w2992), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g2643 (.Q(w3020), .D(w2994), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2644 (.Q(w2994), .D(w2741), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2645 (.Q(w2741), .D(w108), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2646 (.Q(w2716), .D(w2715), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2647 (.Q(w2721), .D(w2864), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2648 (.Q(w2780), .D(w2976), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2649 (.Q(w2784), .D(w2991), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2650 (.Q(w2799), .D(w2792), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2651 (.Q(w2715), .D(w2795), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2652 (.Q(w2820), .D(w2797), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2653 (.Q(w2819), .D(w2865), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2654 (.Q(PLANE_A_PRIO), .D(w2811), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2655 (.Q(PLANE_B_PRIO), .D(w2812), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2656 (.Q(w2776), .D(w2813), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2657 (.Q(w2818), .D(w2817), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2658 (.Q(w2737), .D(w2816), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2659 (.Q(w2816), .D(w130), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2660 (.Q(w2738), .D(w3022), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2661 (.Q(w3022), .D(w129), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2662 (.Q(w2829), .D(w2802), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2663 (.Q(w2815), .D(w2814), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2664 (.Q(SPR_PRIO), .D(w2968), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2665 (.Q(w2826), .D(w175), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2666 (.Q(w2825), .D(w174), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2667 (.Q(w2730), .D(w2746), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2668 (.Q(w2735), .D(w2747), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2669 (.Q(w2732), .D(w2757), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2670 (.Q(w2723), .D(w2748), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2671 (.Q(w2742), .D(w2755), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2672 (.Q(w2722), .D(w2749), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2673 (.Q(w2717), .D(w2852), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2674 (.Q(w2727), .D(w2750), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2675 (.Q(w2733), .D(w2744), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_slatch g2676 (.nQ(w3018), .D(w2746), .C(w2743), .nC(w2740) );
	vdp_slatch g2677 (.nQ(w3019), .D(w2744), .C(w2743), .nC(w2740) );
	vdp_slatch g2678 (.nQ(w3017), .D(w2747), .C(w2743), .nC(w2740) );
	vdp_slatch g2679 (.nQ(w3016), .D(w2757), .C(w2743), .nC(w2740) );
	vdp_slatch g2680 (.nQ(w3015), .D(w2748), .C(w2743), .nC(w2740) );
	vdp_slatch g2681 (.nQ(w3014), .D(w2755), .C(w2743), .nC(w2740) );
	vdp_slatch g2682 (.nQ(w3013), .D(w2749), .C(w2743), .nC(w2740) );
	vdp_slatch g2683 (.nQ(w3012), .D(w2852), .C(w2743), .nC(w2740) );
	vdp_slatch g2684 (.nQ(w3011), .D(w2750), .C(w2743), .nC(w2740) );
	vdp_slatch g2685 (.Q(w2801), .D(REG_BUS[7]), .nC(w2779), .C(w2789) );
	vdp_slatch g2686 (.Q(w2798), .D(REG_BUS[5]), .nC(w2779), .C(w2789) );
	vdp_slatch g2687 (.Q(w2791), .D(REG_BUS[4]), .nC(w2779), .C(w2789) );
	vdp_slatch g2688 (.Q(w2787), .D(REG_BUS[3]), .nC(w2779), .C(w2789) );
	vdp_slatch g2689 (.Q(w2783), .D(REG_BUS[2]), .nC(w2779), .C(w2789) );
	vdp_slatch g2690 (.Q(w2979), .D(REG_BUS[1]), .nC(w2779), .C(w2789) );
	vdp_slatch g2691 (.Q(w2781), .D(REG_BUS[0]), .nC(w2779), .C(w2789) );
	vdp_slatch g2692 (.Q(w2954), .D(REG_BUS[6]), .nC(w2779), .C(w2789) );
	vdp_aon2222 g2693 (.Z(w2931), .B2(w2870), .B1(w2875), .A2(w3006), .A1(w2870), .D2(w2866), .D1(w2875), .C2(w2875), .C1(w2867) );
	vdp_aon22 g2694 (.Z(w2896), .B2(w2866), .B1(w2880), .A2(w3007), .A1(w2871) );
	vdp_aon22 g2695 (.Z(w2901), .B2(w2866), .B1(w2876), .A2(w3006), .A1(w2871) );
	vdp_not g2696 (.nZ(w2884), .A(w2930) );
	vdp_not g2697 (.nZ(w2878), .A(w2879) );
	vdp_not g2698 (.nZ(w2883), .A(w2882) );
	vdp_not g2699 (.nZ(w2902), .A(w2931) );
	vdp_not g2700 (.nZ(w2895), .A(w2888) );
	vdp_buf g2701 (.Z(w2870), .A(w2766) );
	vdp_not g2702 (.nZ(w2965), .A(w2923) );
	vdp_not g2703 (.nZ(w2926), .A(w2924) );
	vdp_not g2704 (.nZ(w2927), .A(w2928) );
	vdp_not g2705 (.nZ(w2891), .A(w2867) );
	vdp_sr_bit g2706 (.Q(w2890), .D(w2738), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2707 (.Q(w2928), .D(w2736), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2708 (.Q(w2867), .D(w2737), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2709 (.Q(w2923), .D(w2925), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2710 (.Q(w2924), .D(w2762), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g2711 (.Z(w3002), .A(w2927), .B(w2965), .C(w2924) );
	vdp_and3 g2712 (.Z(w3004), .A(w2926), .B(w2928), .C(w2965) );
	vdp_and3 g2713 (.Z(w3003), .A(w2927), .B(w2965), .C(w2926) );
	vdp_and3 g2714 (.Z(w2889), .A(w2965), .B(w2924), .C(w2928) );
	vdp_and3 g2715 (.Z(w2887), .A(w2927), .B(w2923), .C(w2926) );
	vdp_and3 g2716 (.Z(w2885), .A(w2923), .B(w2924), .C(w2928) );
	vdp_and3 g2717 (.Z(w3005), .A(w2927), .B(w2924), .C(w2923) );
	vdp_and3 g2718 (.Z(w2886), .A(w2926), .B(w2928), .C(w2923) );
	vdp_sr_bit g2719 (.Q(w2882), .D(w2929), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2720 (.Q(w2879), .D(w2726), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2721 (.Q(w2930), .D(w2763), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g2722 (.Z(w2881), .A(w2883), .B(w2884), .C(w2878) );
	vdp_and3 g2723 (.Z(w2880), .A(w2878), .B(w2882), .C(w2884) );
	vdp_and3 g2724 (.Z(w3007), .A(w2883), .B(w2884), .C(w2879) );
	vdp_and3 g2725 (.Z(w2876), .A(w2884), .B(w2879), .C(w2882) );
	vdp_and3 g2726 (.Z(w2877), .A(w2878), .B(w2882), .C(w2930) );
	vdp_and3 g2727 (.Z(w2874), .A(w2883), .B(w2930), .C(w2878) );
	vdp_and3 g2728 (.Z(w3006), .A(w2883), .B(w2879), .C(w2930) );
	vdp_and3 g2729 (.Z(w2875), .A(w2930), .B(w2879), .C(w2882) );
	vdp_not g2730 (.nZ(w2964), .A(w3021) );
	vdp_not g2731 (.nZ(w2919), .A(w2921) );
	vdp_not g2732 (.nZ(w2920), .A(w2922) );
	vdp_sr_bit g2733 (.Q(w2921), .D(w2960), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2734 (.Q(w2922), .D(w2958), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g2735 (.Q(w3021), .D(w2724), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and3 g2736 (.Z(w2873), .A(w2920), .B(w2964), .C(w2919) );
	vdp_and3 g2737 (.Z(w2872), .A(w2919), .B(w2922), .C(w2964) );
	vdp_and3 g2738 (.A(w2920), .B(w2964), .C(w2921), .Z(w2869) );
	vdp_and3 g2739 (.Z(w3008), .A(w2964), .B(w2921), .C(w2922) );
	vdp_and3 g2740 (.Z(w2868), .A(w2920), .B(w3021), .C(w2919) );
	vdp_and3 g2741 (.Z(w3010), .A(w2919), .B(w2922), .C(w3021) );
	vdp_and3 g2742 (.Z(w2963), .A(w3021), .B(w2921), .C(w2922) );
	vdp_and3 g2743 (.Z(w3009), .A(w2920), .B(w2921), .C(w3021) );
	vdp_aon22 g2744 (.nZ(w2953), .B2(w2866), .B1(w3009), .A2(w3010), .A1(w2867) );
	vdp_aon22 g2745 (.nZ(w2918), .B2(w2866), .B1(w2868), .A2(w2872), .A1(w2867) );
	vdp_aon22 g2746 (.nZ(w2952), .B2(w2867), .B1(w2873), .A2(w2963), .A1(w2871) );
	vdp_and g2747 (.nZ(w2917), .B(w2867), .A(w2868) );
	vdp_and g2748 (.nZ(w2951), .B(w2867), .A(w3009) );
	vdp_and g2749 (.nZ(w2950), .B(w2867), .A(w2869) );
	vdp_aon22 g2750 (.nZ(w2949), .B2(w2870), .B1(w3010), .A2(w2868), .A1(w2870) );
	vdp_aon22 g2751 (.nZ(w2948), .B2(w2866), .B1(w3010), .A2(w3008), .A1(w2867) );
	vdp_aon2222 g2752 (.Z(w2932), .B2(w2870), .B1(w2963), .A2(w3009), .A1(w2870), .D2(w2866), .D1(w2963), .C2(w2963), .C1(w2867) );
	vdp_aon22 g2753 (.Z(w2915), .B2(w2866), .B1(w2872), .A2(w2869), .A1(w2871) );
	vdp_aon22 g2754 (.Z(w2912), .B2(w2866), .B1(w3008), .A2(w3009), .A1(w2871) );
	vdp_and g2755 (.Z(w2916), .B(w3010), .A(w2871) );
	vdp_and g2756 (.Z(w2911), .B(w2871), .A(w3008) );
	vdp_and g2757 (.Z(w2913), .B(w2872), .A(w2871) );
	vdp_aon22 g2758 (.Z(w2910), .B2(w2870), .B1(w3008), .A2(w2869), .A1(w2870) );
	vdp_aon22 g2759 (.Z(w2909), .B2(w2866), .B1(w2869), .A2(w2868), .A1(w2871) );
	vdp_aon2222 g2760 (.Z(w2947), .B2(w2870), .B1(w2872), .A2(w2873), .A1(w2870), .D2(w2866), .D1(w2873), .C2(w2873), .C1(w2871) );
	vdp_not g2761 (.nZ(w2914), .A(w2932) );
	vdp_aon22 g2762 (.nZ(w2946), .B2(w2866), .B1(w3006), .A2(w2877), .A1(w2867) );
	vdp_aon22 g2763 (.nZ(w2945), .B2(w2866), .B1(w2874), .A2(w2880), .A1(w2867) );
	vdp_aon22 g2764 (.nZ(w2908), .B2(w2867), .B1(w2881), .A2(w2875), .A1(w2871) );
	vdp_and g2765 (.nZ(w2907), .B(w2867), .A(w2874) );
	vdp_and g2766 (.nZ(w2906), .B(w2867), .A(w3006) );
	vdp_and g2767 (.nZ(w2905), .B(w2867), .A(w3007) );
	vdp_aon22 g2768 (.nZ(w2904), .B2(w2870), .B1(w2877), .A2(w2874), .A1(w2870) );
	vdp_aon22 g2769 (.nZ(w2903), .B2(w2866), .B1(w2877), .A2(w2876), .A1(w2867) );
	vdp_and g2770 (.Z(w2900), .B(w2877), .A(w2871) );
	vdp_and g2771 (.Z(w2999), .B(w2871), .A(w2876) );
	vdp_and g2772 (.Z(w2899), .B(w2880), .A(w2871) );
	vdp_aon22 g2773 (.Z(w2898), .B2(w2870), .B1(w2876), .A2(w3007), .A1(w2870) );
	vdp_aon22 g2774 (.Z(w2897), .B2(w2866), .B1(w3007), .A2(w2874), .A1(w2871) );
	vdp_aon2222 g2775 (.Z(w3000), .B2(w2870), .B1(w2880), .A2(w2881), .A1(w2870), .D2(w2866), .D1(w2881), .C2(w2881), .C1(w2871) );
	vdp_aon22 g2776 (.nZ(w2894), .B2(w2866), .B1(w3005), .A2(w2886), .A1(w2867) );
	vdp_aon22 g2777 (.nZ(w2944), .B2(w2866), .B1(w2887), .A2(w3004), .A1(w2867) );
	vdp_aon22 g2778 (.nZ(w2940), .B2(w2867), .B1(w3003), .A2(w2885), .A1(w2871) );
	vdp_and g2779 (.nZ(w2941), .B(w2867), .A(w2887) );
	vdp_and g2780 (.nZ(w2942), .B(w2867), .A(w3005) );
	vdp_and g2781 (.nZ(w2939), .B(w2867), .A(w3002) );
	vdp_aon22 g2782 (.nZ(w2943), .B2(w2870), .B1(w2886), .A2(w2887), .A1(w2870) );
	vdp_aon22 g2783 (.nZ(w3001), .B2(w2866), .B1(w2886), .A2(w2889), .A1(w2867) );
	vdp_aon2222 g2784 (.Z(w2888), .B2(w2870), .B1(w2885), .A2(w3005), .A1(w2870), .D2(w2866), .D1(w2885), .C2(w2885), .C1(w2867) );
	vdp_aon22 g2785 (.Z(w2892), .B2(w2866), .B1(w3004), .A2(w3002), .A1(w2871) );
	vdp_aon22 g2786 (.Z(w2893), .B2(w2870), .B1(w2889), .A2(w3002), .A1(w2870) );
	vdp_aon22 g2787 (.Z(w2938), .B2(w2866), .B1(w2889), .A2(w3005), .A1(w2871) );
	vdp_and g2788 (.Z(w2937), .B(w2871), .A(w2889) );
	vdp_and g2789 (.Z(w2936), .B(w3004), .A(w2871) );
	vdp_and g2790 (.Z(w2935), .B(w2871), .A(w2886) );
	vdp_aon22 g2791 (.Z(w2933), .B2(w2866), .B1(w3002), .A2(w2887), .A1(w2871) );
	vdp_aon2222 g2792 (.Z(w2934), .B2(w2870), .B1(w3004), .A2(w3003), .A1(w2870), .D2(w2866), .D1(w3003), .C2(w3003), .C1(w2871) );
	vdp_nor3 g2793 (.Z(w2866), .A(w2870), .B(w2890), .C(w2867) );
	vdp_and g2794 (.Z(w2871), .A(w2890), .B(w2891) );
	vdp_bufif0 g2795 (.A(w2781), .nE(w2788), .Z(COL[0]) );
	vdp_bufif0 g2796 (.A(w2979), .nE(w2788), .Z(COL[1]) );
	vdp_bufif0 g2797 (.A(w2783), .nE(w2788), .Z(COL[2]) );
	vdp_bufif0 g2798 (.A(w2787), .nE(w2788), .Z(COL[3]) );
	vdp_bufif0 g2799 (.A(w2800), .nE(w2788), .Z(COL[4]) );
	vdp_bufif0 g2800 (.A(w2978), .nE(w2788), .Z(COL[5]) );
	vdp_and g2801 (.Z(w2978), .A(M5), .B(w2798) );
	vdp_or g2802 (.Z(w2800), .A(w2771), .B(w2791) );
	vdp_not g2803 (.nZ(w2666), .A(M5) );
	vdp_not g2804 (.nZ(w2769), .A(w2977) );
	vdp_not g2805 (.nZ(w2770), .A(w2772) );
	vdp_not g2806 (.nZ(w2771), .A(M5) );
	vdp_not g2807 (.nZ(w2767), .A(w2773) );
	vdp_not g2808 (.nZ(w2788), .A(w2776) );
	vdp_comp_strong g2809 (.nZ(w2779), .Z(w2789), .A(w73) );
	vdp_not g2810 (.nZ(w2777), .A(w101) );
	vdp_not g2811 (.nZ(w2990), .A(w19) );
	vdp_aon222 g2812 (.Z(w2976), .B2(w2769), .A2(w2770), .A1(VRAMA[0]), .B1(VRAMA[1]), .C2(w2767), .C1(COL[0]) );
	vdp_aon222 g2813 (.Z(w2991), .B2(w2769), .A2(w2770), .A1(VRAMA[1]), .B1(VRAMA[2]), .C2(w2767), .C1(COL[1]) );
	vdp_aon222 g2814 (.Z(w2782), .B2(w2769), .A2(w2770), .A1(VRAMA[2]), .B1(VRAMA[3]), .C2(w2767), .C1(COL[2]) );
	vdp_aon222 g2815 (.Z(w2792), .B2(w2769), .A2(w2770), .A1(VRAMA[3]), .B1(VRAMA[4]), .C2(w2767), .C1(COL[3]) );
	vdp_aon222 g2816 (.Z(w2797), .B2(w2769), .A2(w2770), .A1(VRAMA[4]), .B1(VRAMA[5]), .C2(w2767), .C1(COL[4]) );
	vdp_aon222 g2817 (.Z(w2865), .B2(w2769), .A2(w2770), .A1(1'b0), .B1(VRAMA[6]), .C2(w2767), .C1(COL[5]) );
	vdp_nand g2818 (.Z(w2977), .A(w2773), .B(M5) );
	vdp_nand g2819 (.Z(w2772), .A(w2773), .B(w2771) );
	vdp_and g2820 (.Z(w2802), .A(w2803), .B(w3029) );
	vdp_aon222 g2821 (.Z(w3029), .B2(w3024), .A2(w2808), .A1(w2764), .B1(w2810), .C2(w3023), .C1(w2831) );
	vdp_not g2822 (.nZ(w3024), .A(w2975) );
	vdp_not g2823 (.nZ(w3023), .A(w2765) );
	vdp_not g2824 (.nZ(w2836), .A(w2821) );
	vdp_nor g2825 (.Z(w2810), .A(w2765), .B(w2968) );
	vdp_nor g2826 (.Z(w2975), .A(w2831), .B(w2830) );
	vdp_and g2827 (.Z(w2809), .A(w2804), .B(w2844) );
	vdp_and g2828 (.Z(w2808), .A(w2821), .B(w2835) );
	vdp_and g2829 (.Z(w2838), .A(w2835), .B(w2836) );
	vdp_or g2830 (.Z(w2968), .A(w2839), .B(w2838) );
	vdp_or g2831 (.Z(w2807), .A(w2764), .B(w2765) );
	vdp_and g2832 (.Z(w2778), .A(w2803), .B(w2777) );
	vdp_and g2833 (.Z(w2957), .A(w2804), .B(w2841) );
	vdp_and g2834 (.Z(w2967), .A(w2805), .B(w2843) );
	vdp_not g2835 (.nZ(w2849), .A(w101) );
	vdp_or g2836 (.Z(w2811), .A(w2842), .B(w2828) );
	vdp_not g2837 (.nZ(w3027), .A(w2805) );
	vdp_not g2838 (.nZ(w2955), .A(w2705) );
	vdp_not g2839 (.nZ(w2833), .A(w2822) );
	vdp_not g2840 (.nZ(w2832), .A(w2823) );
	vdp_not g2841 (.nZ(w2837), .A(w2706) );
	vdp_and g2842 (.Z(w2856), .A(w2805), .B(w2840) );
	vdp_and g2843 (.Z(w2834), .A(w2806), .B(w2846) );
	vdp_not g2844 (.nZ(w2966), .A(w98) );
	vdp_not g2845 (.nZ(w2973), .A(w99) );
	vdp_and g2846 (.Z(w2839), .A(w2973), .B(w98) );
	vdp_and g2847 (.Z(w2842), .A(w2966), .B(w99) );
	vdp_and g2848 (.Z(w2855), .A(w98), .B(w99) );
	vdp_or3 g2849 (.Z(w2773), .A(w108), .B(w174), .C(w175) );
	vdp_and3 g2850 (.Z(w2972), .A(w2806), .B(w2805), .C(w2843) );
	vdp_and3 g2851 (.Z(w2841), .A(w2832), .B(w2822), .C(w2706) );
	vdp_and3 g2852 (.Z(w2840), .A(w2833), .B(w2823), .C(w2837) );
	vdp_and3 g2853 (.Z(w2846), .A(w2832), .B(w2822), .C(w2837) );
	vdp_and3 g2854 (.Z(w2843), .A(w2822), .B(w2823), .C(w2837) );
	vdp_and g2855 (.Z(w2962), .A(M5), .B(w89) );
	vdp_or g2856 (.Z(w2804), .A(w2955), .B(w2821) );
	vdp_and3 g2857 (.Z(w2814), .A(w2808), .B(w2765), .C(w2975) );
	vdp_and3 g2858 (.Z(w2971), .A(w2806), .B(w2804), .C(w2841) );
	vdp_and3 g2859 (.Z(w2970), .A(w2806), .B(w2804), .C(w2846) );
	vdp_and3 g2860 (.Z(w2828), .A(w2827), .B(w2778), .C(w3027) );
	vdp_and3 g2861 (.Z(w2821), .A(w2807), .B(w2824), .C(w2962) );
	vdp_and3 g2862 (.Z(w2850), .A(w2805), .B(w2804), .C(w2844) );
	vdp_and3 g2863 (.Z(w3026), .A(w2805), .B(w2804), .C(w2840) );
	vdp_and3 g2864 (.Z(w2847), .A(w2806), .B(w2805), .C(w2804) );
	vdp_and3 g2865 (.Z(w2848), .A(w2778), .B(w2845), .C(w3025) );
	vdp_and g2866 (.Z(w2813), .A(w2956), .B(w2969) );
	vdp_not g2867 (.nZ(w2851), .A(w2778) );
	vdp_not g2868 (.nZ(w3025), .A(w2806) );
	vdp_or g2869 (.Z(w2812), .A(w2855), .B(w2848) );
	vdp_or g2870 (.Z(w2969), .A(w2851), .B(w2847) );
	vdp_not g2871 (.nZ(w2982), .A(M5) );
	vdp_notif0 g2872 (.A(w3019), .nE(w2745), .nZ(w324) );
	vdp_notif0 g2873 (.nZ(RD_DATA[2]), .A(w3018), .nE(w2745) );
	vdp_notif0 g2874 (.nZ(RD_DATA[1]), .A(w3017), .nE(w2745) );
	vdp_notif0 g2875 (.nZ(AD_DATA[7]), .A(w3016), .nE(w2745) );
	vdp_notif0 g2876 (.nZ(AD_DATA[6]), .A(w3015), .nE(w2745) );
	vdp_notif0 g2877 (.nZ(AD_DATA[5]), .A(w3014), .nE(w2745) );
	vdp_notif0 g2878 (.nZ(AD_DATA[3]), .A(w3013), .nE(w2745) );
	vdp_notif0 g2879 (.nZ(AD_DATA[2]), .A(w3012), .nE(w2745) );
	vdp_notif0 g2880 (.nZ(AD_DATA[1]), .A(w3011), .nE(w2745) );
	vdp_notif0 g2881 (.nZ(DB[1]), .A(w2738), .nE(w2729) );
	vdp_notif0 g2882 (.A(w2737), .nE(w2729) );
	vdp_notif0 g2883 (.nZ(DB[2]), .A(w2958), .nE(w2729) );
	vdp_notif0 g2884 (.nZ(DB[5]), .A(w2929), .nE(w2729) );
	vdp_notif0 g2885 (.nZ(DB[8]), .A(w2736), .nE(w2729) );
	vdp_notif0 g2886 (.nZ(DB[10]), .A(w2925), .nE(w2729) );
	vdp_notif0 g2887 (.nZ(DB[9]), .A(w2762), .nE(w2729) );
	vdp_notif0 g2888 (.nZ(DB[7]), .A(w2763), .nE(w2729) );
	vdp_notif0 g2889 (.nZ(DB[6]), .A(w2726), .nE(w2729) );
	vdp_notif0 g2890 (.nZ(DB[4]), .A(w2724), .nE(w2729) );
	vdp_comp_we g2891 (.A(M5), .nZ(w2719), .Z(w2718) );
	vdp_notif0 g2892 (.nZ(DB[3]), .A(w2960), .nE(w2729) );
	vdp_not g2893 (.A(w88), .nZ(w2729) );
	vdp_and g2894 (.Z(w2720), .A(w2721), .B(w2716) );
	vdp_and3 g2895 (.Z(w2960), .A(w97), .B(w2721), .C(w2959) );
	vdp_and3 g2896 (.Z(w2724), .A(w97), .B(w2721), .C(w2993) );
	vdp_and3 g2897 (.Z(w2726), .A(w97), .B(w2721), .C(w2725) );
	vdp_and3 g2898 (.Z(w2763), .A(w97), .B(w2721), .C(w2728) );
	vdp_and3 g2899 (.Z(w2762), .A(w97), .B(w2721), .C(w2731) );
	vdp_and3 g2900 (.Z(w2925), .A(w97), .B(w2721), .C(w2734) );
	vdp_and3 g2901 (.Z(w2736), .A(M5), .B(w2721), .C(w2735) );
	vdp_and3 g2902 (.Z(w2929), .A(M5), .B(w2721), .C(w2742) );
	vdp_and3 g2903 (.Z(w2958), .A(M5), .B(w2721), .C(w2727) );
	vdp_comp_strong g2904 (.nZ(w2740), .A(w2739), .Z(w2743) );
	vdp_and g2905 (.Z(w2739), .A(w2741), .B(HCLK1) );
	vdp_not g2906 (.nZ(w2745), .A(w3020) );
	vdp_aon22 g2907 (.Z(w2981), .B2(FIFOo[5]), .A2(FIFOo[7]), .A1(w2794), .B1(w2793) );
	vdp_aon22 g2908 (.Z(w2756), .B2(FIFOo[4]), .A2(FIFOo[6]), .A1(w2794), .B1(w2793) );
	vdp_aon22 g2909 (.Z(w2754), .B2(FIFOo[3]), .A2(FIFOo[5]), .A1(w2794), .B1(w2793) );
	vdp_aon22 g2910 (.Z(w2753), .B2(FIFOo[2]), .A2(FIFOo[3]), .A1(w2794), .B1(w2793) );
	vdp_aon22 g2911 (.Z(w2752), .B2(FIFOo[1]), .A2(FIFOo[2]), .A1(w2794), .B1(w2793) );
	vdp_aon22 g2912 (.Z(w2751), .B2(FIFOo[0]), .A2(FIFOo[1]), .A1(w2794), .B1(w2793) );
	vdp_comp_we g2913 (.Z(w2794), .nZ(w2793), .A(M5) );
	vdp_aon22 g2914 (.Z(w2785), .B2(w2982), .A2(M5), .A1(w2961), .B1(w18) );
	vdp_aon22 g2915 (.Z(w130), .B2(w2815), .A2(w2801), .A1(w101), .B1(w2849) );
	vdp_aon22 g2916 (.Z(w129), .B2(w2829), .A2(w2954), .A1(w101), .B1(w2849) );
	vdp_and3 g2917 (.Z(w2835), .A(w2778), .B(w2705), .C(w3028) );
	vdp_aon22 g2918 (.Z(w2844), .B2(w2832), .A2(w2823), .A1(w2706), .B1(w2833) );
	vdp_aon22 g2919 (.Z(w2728), .B2(w2742), .A2(w2732), .A1(w2718), .B1(w2719) );
	vdp_aon22 g2920 (.Z(w2725), .B2(w2722), .A2(w2723), .A1(w2718), .B1(w2719) );
	vdp_aon22 g2921 (.Z(w2959), .B2(w2727), .A2(w2717), .A1(w2718), .B1(w2719) );
	vdp_aon22 g2922 (.Z(w2993), .B2(w2717), .A2(w2722), .A1(w2718), .B1(w2719) );
	vdp_aon22 g2923 (.Z(w2731), .B2(w2723), .A2(w2730), .A1(w2718), .B1(w2719) );
	vdp_aon22 g2924 (.Z(w2734), .B2(w2732), .A2(w2733), .A1(w2718), .B1(w2719) );
	vdp_g2925 g2925 (.Z(w2830), .A(w2833), .B(w2706), .C(w2962), .D(w2832) );
	vdp_or5 g2926 (.Z(w2827), .A(w2809), .B(w2840), .C(w2843), .D(w2971), .E(w2970) );
	vdp_or5 g2927 (.Z(w2845), .A(w2850), .B(w2846), .C(w2957), .D(w2967), .E(w3026) );
	vdp_or5 g2928 (.Z(w3028), .A(w2841), .B(w2844), .C(w2856), .D(w2834), .E(w2972) );
	vdp_nor4 g2929 (.Z(w2795), .A(COL[2]), .B(COL[3]), .C(COL[1]), .D(COL[0]) );
	vdp_nor g2930 (.Z(w2956), .A(w98), .B(w99) );
	vdp_nor g2931 (.Z(w2805), .A(w2974), .B(w2854) );
	vdp_nor g2932 (.Z(w2974), .A(w2705), .B(M5) );
	vdp_nand g2933 (.Z(w2806), .A(M5), .B(w2853) );
	vdp_nand g2934 (.Z(w2817), .A(SPR_PRIO), .B(w19) );
	vdp_and4 g2935 (.Z(w2831), .A(w2832), .B(w2962), .C(w2833), .D(w2837) );
	vdp_aoi21 g2936 (.Z(w2992), .B(w2720), .A2(w2990), .A1(w2768) );
	vdp_nor g2937 (.Z(w2864), .A(w21), .B(w20) );
	vdp_g2938 g2938 (.A(w2776), .Z(COL[6]) );
	vdp_slatch g2939 (.Q(w4136), .D(S[3]), .C(w3156), .nC(w3146) );
	vdp_slatch g2940 (.Q(w4138), .D(S[3]), .C(w3137), .nC(w3136) );
	vdp_slatch g2941 (.Q(w4140), .D(S[3]), .C(w3138), .nC(w3134) );
	vdp_slatch g2942 (.Q(w4142), .D(S[3]), .C(w3155), .nC(w3147) );
	vdp_slatch g2943 (.Q(w4144), .D(S[7]), .C(w3156), .nC(w3146) );
	vdp_slatch g2944 (.Q(w4147), .D(S[7]), .C(w3137), .nC(w3136) );
	vdp_slatch g2945 (.Q(w4146), .D(S[7]), .C(w3138), .nC(w3134) );
	vdp_slatch g2946 (.Q(w4151), .D(S[7]), .C(w3155), .nC(w3147) );
	vdp_slatch g2947 (.Q(w4150), .D(S[2]), .C(w3156), .nC(w3146) );
	vdp_slatch g2948 (.Q(w4157), .D(S[2]), .C(w3137), .nC(w3136) );
	vdp_slatch g2949 (.Q(w4156), .D(S[2]), .C(w3138), .nC(w3134) );
	vdp_slatch g2950 (.Q(w4159), .D(S[2]), .C(w3155), .nC(w3147) );
	vdp_slatch g2951 (.Q(w4158), .D(S[6]), .C(w3156), .nC(w3146) );
	vdp_slatch g2952 (.Q(w4163), .D(S[6]), .C(w3137), .nC(w3136) );
	vdp_slatch g2953 (.Q(w4162), .D(S[6]), .C(w3138), .nC(w3134) );
	vdp_slatch g2954 (.Q(w4167), .D(S[6]), .C(w3155), .nC(w3147) );
	vdp_slatch g2955 (.Q(w4166), .D(S[1]), .C(w3156), .nC(w3146) );
	vdp_slatch g2956 (.Q(w4171), .D(S[1]), .C(w3137), .nC(w3136) );
	vdp_slatch g2957 (.Q(w4170), .D(S[1]), .C(w3138), .nC(w3134) );
	vdp_slatch g2958 (.Q(w4175), .D(S[1]), .C(w3155), .nC(w3147) );
	vdp_slatch g2959 (.Q(w4174), .D(S[5]), .C(w3156), .nC(w3146) );
	vdp_slatch g2960 (.Q(w4179), .D(S[5]), .C(w3137), .nC(w3136) );
	vdp_slatch g2961 (.Q(w4178), .D(S[5]), .C(w3138), .nC(w3134) );
	vdp_slatch g2962 (.Q(w4183), .D(S[5]), .C(w3155), .nC(w3147) );
	vdp_slatch g2963 (.Q(w4182), .D(S[0]), .C(w3156), .nC(w3146) );
	vdp_slatch g2964 (.Q(w4187), .D(S[0]), .C(w3137), .nC(w3136) );
	vdp_slatch g2965 (.Q(w4186), .D(S[0]), .C(w3138), .nC(w3134) );
	vdp_slatch g2966 (.Q(w4191), .D(S[0]), .C(w3155), .nC(w3147) );
	vdp_slatch g2967 (.Q(w4190), .D(S[4]), .C(w3156), .nC(w3146) );
	vdp_slatch g2968 (.Q(w4195), .D(S[4]), .C(w3137), .nC(w3136) );
	vdp_slatch g2969 (.Q(w4194), .D(S[4]), .C(w3138), .nC(w3134) );
	vdp_slatch g2970 (.Q(w4198), .D(S[4]), .C(w3155), .nC(w3147) );
	vdp_slatch g2971 (.Q(w4137), .D(w4136), .C(w3126), .nC(w3143) );
	vdp_slatch g2972 (.Q(w4139), .D(w4138), .C(w3144), .nC(w3135) );
	vdp_slatch g2973 (.Q(w4141), .D(w4140), .C(w3145), .nC(w3133) );
	vdp_slatch g2974 (.Q(w4143), .D(w4142), .C(w3141), .nC(w3142) );
	vdp_slatch g2975 (.Q(w4145), .D(w4144), .C(w3126), .nC(w3143) );
	vdp_slatch g2976 (.Q(w4149), .D(w4147), .C(w3144), .nC(w3135) );
	vdp_slatch g2977 (.Q(w4148), .D(w4146), .C(w3145), .nC(w3133) );
	vdp_slatch g2978 (.Q(w4153), .D(w4151), .C(w3141), .nC(w3142) );
	vdp_slatch g2979 (.Q(w4152), .D(w4150), .C(w3126), .nC(w3143) );
	vdp_slatch g2980 (.Q(w4155), .D(w4157), .C(w3144), .nC(w3135) );
	vdp_slatch g2981 (.Q(w4154), .D(w4156), .C(w3145), .nC(w3133) );
	vdp_slatch g2982 (.Q(w4161), .D(w4159), .C(w3141), .nC(w3142) );
	vdp_slatch g2983 (.Q(w4160), .D(w4158), .C(w3126), .nC(w3143) );
	vdp_slatch g2984 (.Q(w4165), .D(w4163), .C(w3144), .nC(w3135) );
	vdp_slatch g2985 (.Q(w4164), .D(w4162), .C(w3145), .nC(w3133) );
	vdp_slatch g2986 (.Q(w4169), .D(w4167), .C(w3141), .nC(w3142) );
	vdp_slatch g2987 (.Q(w4168), .D(w4166), .C(w3126), .nC(w3143) );
	vdp_slatch g2988 (.Q(w4173), .D(w4171), .C(w3144), .nC(w3135) );
	vdp_slatch g2989 (.Q(w4172), .D(w4170), .C(w3145), .nC(w3133) );
	vdp_slatch g2990 (.Q(w4177), .D(w4175), .C(w3141), .nC(w3142) );
	vdp_slatch g2991 (.Q(w4176), .D(w4174), .C(w3126), .nC(w3143) );
	vdp_slatch g2992 (.Q(w4181), .D(w4179), .C(w3144), .nC(w3135) );
	vdp_slatch g2993 (.Q(w4180), .D(w4178), .C(w3145), .nC(w3133) );
	vdp_slatch g2994 (.Q(w4185), .D(w4183), .C(w3141), .nC(w3142) );
	vdp_slatch g2995 (.Q(w4184), .D(w4182), .C(w3126), .nC(w3143) );
	vdp_slatch g2996 (.Q(w4189), .D(w4187), .C(w3144), .nC(w3135) );
	vdp_slatch g2997 (.Q(w4188), .D(w4186), .C(w3145), .nC(w3133) );
	vdp_slatch g2998 (.Q(w4193), .D(w4191), .C(w3141), .nC(w3142) );
	vdp_slatch g2999 (.Q(w4192), .D(w4190), .C(w3126), .nC(w3143) );
	vdp_slatch g3000 (.Q(w4197), .D(w4195), .C(w3144), .nC(w3135) );
	vdp_slatch g3001 (.Q(w4196), .D(w4194), .C(w3145), .nC(w3133) );
	vdp_slatch g3002 (.Q(w4199), .D(w4198), .C(w3141), .nC(w3142) );
	vdp_slatch g3003 (.Q(w3183), .D(w4137), .C(w3148), .nC(w3174) );
	vdp_slatch g3004 (.Q(w3182), .D(w4139), .C(w3127), .nC(w3184) );
	vdp_slatch g3005 (.Q(w3181), .D(w4141), .C(w3139), .nC(w3185) );
	vdp_slatch g3006 (.Q(w3180), .D(w4143), .C(w3140), .nC(w3114) );
	vdp_slatch g3007 (.Q(w3179), .D(w4145), .C(w3148), .nC(w3174) );
	vdp_slatch g3008 (.Q(w3178), .D(w4149), .C(w3127), .nC(w3184) );
	vdp_slatch g3009 (.Q(w3177), .D(w4148), .C(w3139), .nC(w3185) );
	vdp_slatch g3010 (.Q(w3176), .D(w4153), .C(w3140), .nC(w3114) );
	vdp_slatch g3011 (.Q(w3175), .D(w4152), .C(w3148), .nC(w3174) );
	vdp_slatch g3012 (.Q(w3188), .D(w4155), .C(w3127), .nC(w3184) );
	vdp_slatch g3013 (.Q(w3192), .D(w4154), .C(w3139), .nC(w3185) );
	vdp_slatch g3014 (.Q(w3191), .D(w4161), .C(w3140), .nC(w3114) );
	vdp_slatch g3015 (.Q(w3190), .D(w4160), .C(w3148), .nC(w3174) );
	vdp_slatch g3016 (.Q(w3186), .D(w4165), .C(w3127), .nC(w3184) );
	vdp_slatch g3017 (.Q(w3187), .D(w4164), .C(w3139), .nC(w3185) );
	vdp_slatch g3018 (.D(w4169), .Q(w3189), .C(w3140), .nC(w3114) );
	vdp_slatch g3019 (.Q(w3193), .D(w4168), .C(w3148), .nC(w3174) );
	vdp_slatch g3020 (.Q(w3194), .D(w4173), .C(w3127), .nC(w3184) );
	vdp_slatch g3021 (.Q(w3196), .D(w4172), .C(w3139), .nC(w3185) );
	vdp_slatch g3022 (.Q(w3195), .D(w4177), .C(w3140), .nC(w3114) );
	vdp_slatch g3023 (.Q(w3237), .D(w4176), .C(w3148), .nC(w3174) );
	vdp_slatch g3024 (.Q(w3238), .D(w4181), .C(w3127), .nC(w3184) );
	vdp_slatch g3025 (.Q(w3234), .D(w4180), .C(w3139), .nC(w3185) );
	vdp_slatch g3026 (.Q(w3229), .D(w4185), .C(w3140), .nC(w3114) );
	vdp_slatch g3027 (.Q(w3241), .D(w4184), .C(w3148), .nC(w3174) );
	vdp_slatch g3028 (.Q(w3240), .D(w4189), .C(w3127), .nC(w3184) );
	vdp_slatch g3029 (.Q(w3239), .D(w4188), .C(w3139), .nC(w3185) );
	vdp_slatch g3030 (.Q(w3236), .D(w4193), .C(w3140), .nC(w3114) );
	vdp_slatch g3031 (.Q(w3222), .D(w4192), .C(w3148), .nC(w3174) );
	vdp_slatch g3032 (.Q(w3221), .D(w4197), .C(w3127), .nC(w3184) );
	vdp_slatch g3033 (.Q(w3223), .D(w4196), .C(w3139), .nC(w3185) );
	vdp_slatch g3034 (.Q(w3224), .D(w4199), .C(w3140), .nC(w3114) );
	vdp_slatch g3035 (.Q(w3301), .D(w4421), .C(w3298), .nC(w3299) );
	vdp_slatch g3036 (.Q(w3302), .D(w4422), .C(w3297), .nC(w3307) );
	vdp_slatch g3037 (.Q(w3303), .D(w4424), .C(w3296), .nC(w3308) );
	vdp_slatch g3038 (.Q(w3304), .D(w4423), .C(w3295), .nC(w3300) );
	vdp_slatch g3039 (.Q(w3305), .D(w4255), .C(w3298), .nC(w3299) );
	vdp_slatch g3040 (.Q(w3306), .D(w4254), .C(w3297), .nC(w3307) );
	vdp_slatch g3041 (.Q(w3312), .D(w4249), .C(w3296), .nC(w3308) );
	vdp_slatch g3042 (.Q(w3313), .D(w4248), .C(w3295), .nC(w3300) );
	vdp_slatch g3043 (.Q(w3314), .D(w4245), .C(w3298), .nC(w3299) );
	vdp_slatch g3044 (.Q(w3315), .D(w4244), .C(w3297), .nC(w3307) );
	vdp_slatch g3045 (.Q(w3316), .D(w4243), .C(w3296), .nC(w3308) );
	vdp_slatch g3046 (.Q(w3311), .D(w4240), .C(w3295), .nC(w3300) );
	vdp_slatch g3047 (.Q(w3317), .D(w4237), .C(w3298), .nC(w3299) );
	vdp_slatch g3048 (.Q(w3318), .D(w4238), .C(w3297), .nC(w3307) );
	vdp_slatch g3049 (.Q(w3319), .D(w4233), .C(w3296), .nC(w3308) );
	vdp_slatch g3050 (.Q(w3320), .D(w4234), .C(w3295), .nC(w3300) );
	vdp_slatch g3051 (.Q(w3245), .D(w4231), .C(w3298), .nC(w3299) );
	vdp_slatch g3052 (.Q(w4023), .D(w4230), .C(w3297), .nC(w3307) );
	vdp_slatch g3053 (.Q(w3247), .D(w4227), .C(w3296), .nC(w3308) );
	vdp_slatch g3054 (.Q(w3248), .D(w4226), .C(w3295), .nC(w3300) );
	vdp_slatch g3055 (.Q(w3321), .D(w4223), .C(w3298), .nC(w3299) );
	vdp_slatch g3056 (.Q(w3246), .D(w4222), .C(w3297), .nC(w3307) );
	vdp_slatch g3057 (.Q(w3226), .D(w4219), .C(w3296), .nC(w3308) );
	vdp_slatch g3058 (.Q(w3249), .D(w4218), .C(w3295), .nC(w3300) );
	vdp_slatch g3059 (.Q(w3252), .D(w4215), .C(w3298), .nC(w3299) );
	vdp_slatch g3060 (.Q(w3260), .D(w4214), .C(w3297), .nC(w3307) );
	vdp_slatch g3061 (.Q(w3259), .D(w4211), .C(w3296), .nC(w3308) );
	vdp_slatch g3062 (.Q(w3258), .D(w4210), .C(w3295), .nC(w3300) );
	vdp_slatch g3063 (.Q(w3256), .D(w4207), .C(w3298), .nC(w3299) );
	vdp_slatch g3064 (.Q(w3250), .D(w4206), .C(w3297), .nC(w3307) );
	vdp_slatch g3065 (.Q(w3257), .D(w4203), .C(w3296), .nC(w3308) );
	vdp_slatch g3066 (.Q(w3251), .D(w4202), .C(w3295), .nC(w3300) );
	vdp_slatch g3067 (.Q(w4421), .D(w4258), .C(w3291), .nC(w3285) );
	vdp_slatch g3068 (.Q(w4422), .D(w4259), .C(w3106), .nC(w3286) );
	vdp_slatch g3069 (.Q(w4424), .D(w4257), .C(w3293), .nC(w3094) );
	vdp_slatch g3070 (.Q(w4423), .D(w4256), .C(w3294), .nC(w3095) );
	vdp_slatch g3071 (.Q(w4255), .D(w4253), .C(w3291), .nC(w3285) );
	vdp_slatch g3072 (.Q(w4254), .D(w4252), .C(w3106), .nC(w3286) );
	vdp_slatch g3073 (.Q(w4249), .D(w4251), .C(w3293), .nC(w3094) );
	vdp_slatch g3074 (.Q(w4248), .D(w4250), .C(w3294), .nC(w3095) );
	vdp_slatch g3075 (.Q(w4245), .D(w4247), .C(w3291), .nC(w3285) );
	vdp_slatch g3076 (.Q(w4244), .D(w4246), .C(w3106), .nC(w3286) );
	vdp_slatch g3077 (.Q(w4243), .D(w4241), .C(w3293), .nC(w3094) );
	vdp_slatch g3078 (.Q(w4240), .D(w4242), .C(w3294), .nC(w3095) );
	vdp_slatch g3079 (.Q(w4237), .D(w4239), .C(w3291), .nC(w3285) );
	vdp_slatch g3080 (.Q(w4238), .D(w4236), .C(w3106), .nC(w3286) );
	vdp_slatch g3081 (.Q(w4233), .D(w4235), .C(w3293), .nC(w3094) );
	vdp_slatch g3082 (.Q(w4234), .D(w4232), .C(w3294), .nC(w3095) );
	vdp_slatch g3083 (.Q(w4231), .D(w4229), .C(w3291), .nC(w3285) );
	vdp_slatch g3084 (.Q(w4230), .D(w4228), .C(w3106), .nC(w3286) );
	vdp_slatch g3085 (.Q(w4227), .D(w4225), .C(w3293), .nC(w3094) );
	vdp_slatch g3086 (.Q(w4226), .D(w4224), .C(w3294), .nC(w3095) );
	vdp_slatch g3087 (.Q(w4223), .D(w4221), .C(w3291), .nC(w3285) );
	vdp_slatch g3088 (.Q(w4222), .D(w4220), .C(w3106), .nC(w3286) );
	vdp_slatch g3089 (.Q(w4219), .D(w4217), .C(w3293), .nC(w3094) );
	vdp_slatch g3090 (.Q(w4218), .D(w4216), .C(w3294), .nC(w3095) );
	vdp_slatch g3091 (.Q(w4215), .D(w4213), .C(w3291), .nC(w3285) );
	vdp_slatch g3092 (.Q(w4214), .D(w4212), .C(w3106), .nC(w3286) );
	vdp_slatch g3093 (.Q(w4211), .D(w4209), .C(w3293), .nC(w3094) );
	vdp_slatch g3094 (.Q(w4210), .D(w4208), .C(w3294), .nC(w3095) );
	vdp_slatch g3095 (.Q(w4207), .D(w4205), .C(w3291), .nC(w3285) );
	vdp_slatch g3096 (.Q(w4206), .D(w4204), .C(w3106), .nC(w3286) );
	vdp_slatch g3097 (.Q(w4203), .D(w4201), .C(w3293), .nC(w3094) );
	vdp_slatch g3098 (.Q(w4202), .D(w4200), .C(w3294), .nC(w3095) );
	vdp_slatch g3099 (.Q(w4258), .D(S[3]), .C(w3058), .nC(w3092) );
	vdp_slatch g3100 (.Q(w4259), .D(S[3]), .C(w3062), .nC(w3096) );
	vdp_slatch g3101 (.Q(w4257), .D(S[3]), .C(w3065), .nC(w3093) );
	vdp_slatch g3102 (.Q(w4256), .D(S[3]), .C(w3067), .nC(w3091) );
	vdp_slatch g3103 (.Q(w4253), .D(S[7]), .C(w3058), .nC(w3092) );
	vdp_slatch g3104 (.Q(w4252), .D(S[7]), .C(w3062), .nC(w3096) );
	vdp_slatch g3105 (.Q(w4251), .D(S[7]), .C(w3065), .nC(w3093) );
	vdp_slatch g3106 (.Q(w4250), .D(S[7]), .C(w3067), .nC(w3091) );
	vdp_slatch g3107 (.Q(w4247), .D(S[2]), .C(w3058), .nC(w3092) );
	vdp_slatch g3108 (.Q(w4246), .D(S[2]), .C(w3062), .nC(w3096) );
	vdp_slatch g3109 (.Q(w4241), .D(S[2]), .C(w3065), .nC(w3093) );
	vdp_slatch g3110 (.Q(w4242), .D(S[2]), .C(w3067), .nC(w3091) );
	vdp_slatch g3111 (.Q(w4239), .D(S[6]), .C(w3058), .nC(w3092) );
	vdp_slatch g3112 (.Q(w4236), .D(S[6]), .C(w3062), .nC(w3096) );
	vdp_slatch g3113 (.Q(w4235), .D(S[6]), .C(w3065), .nC(w3093) );
	vdp_slatch g3114 (.Q(w4232), .D(S[6]), .C(w3067), .nC(w3091) );
	vdp_slatch g3115 (.Q(w4229), .D(S[1]), .C(w3058), .nC(w3092) );
	vdp_slatch g3116 (.Q(w4228), .D(S[1]), .C(w3062), .nC(w3096) );
	vdp_slatch g3117 (.Q(w4225), .D(S[1]), .C(w3065), .nC(w3093) );
	vdp_slatch g3118 (.Q(w4224), .D(S[1]), .C(w3067), .nC(w3091) );
	vdp_slatch g3119 (.Q(w4221), .D(S[5]), .C(w3058), .nC(w3092) );
	vdp_slatch g3120 (.Q(w4220), .D(S[5]), .C(w3062), .nC(w3096) );
	vdp_slatch g3121 (.Q(w4217), .D(S[5]), .C(w3065), .nC(w3093) );
	vdp_slatch g3122 (.Q(w4216), .D(S[5]), .C(w3067), .nC(w3091) );
	vdp_slatch g3123 (.Q(w4213), .D(S[0]), .C(w3058), .nC(w3092) );
	vdp_slatch g3124 (.Q(w4212), .D(S[0]), .C(w3062), .nC(w3096) );
	vdp_slatch g3125 (.Q(w4209), .D(S[0]), .C(w3065), .nC(w3093) );
	vdp_slatch g3126 (.Q(w4208), .D(S[0]), .C(w3067), .nC(w3091) );
	vdp_slatch g3127 (.Q(w4205), .D(S[4]), .C(w3058), .nC(w3092) );
	vdp_slatch g3128 (.Q(w4204), .D(S[4]), .C(w3062), .nC(w3096) );
	vdp_slatch g3129 (.Q(w4201), .D(S[4]), .C(w3065), .nC(w3093) );
	vdp_slatch g3130 (.Q(w4200), .D(S[4]), .C(w3067), .nC(w3091) );
	vdp_slatch g3131 (.Q(w4263), .D(S[3]), .C(w3059), .nC(w3084) );
	vdp_slatch g3132 (.Q(w4262), .D(S[3]), .C(w3063), .nC(w3089) );
	vdp_slatch g3133 (.Q(w4267), .D(S[3]), .C(w3064), .nC(w3090) );
	vdp_slatch g3134 (.Q(w4266), .D(S[3]), .C(w3066), .nC(w3085) );
	vdp_slatch g3135 (.Q(w4271), .D(S[7]), .C(w3059), .nC(w3084) );
	vdp_slatch g3136 (.Q(w4270), .D(S[7]), .C(w3063), .nC(w3089) );
	vdp_slatch g3137 (.Q(w4275), .D(S[7]), .C(w3064), .nC(w3090) );
	vdp_slatch g3138 (.Q(w4274), .D(S[7]), .C(w3066), .nC(w3085) );
	vdp_slatch g3139 (.Q(w4279), .D(S[2]), .C(w3059), .nC(w3084) );
	vdp_slatch g3140 (.Q(w4278), .D(S[2]), .C(w3063), .nC(w3089) );
	vdp_slatch g3141 (.Q(w4283), .D(S[2]), .C(w3064), .nC(w3090) );
	vdp_slatch g3142 (.Q(w4282), .D(S[2]), .C(w3066), .nC(w3085) );
	vdp_slatch g3143 (.Q(w4285), .D(S[6]), .C(w3059), .nC(w3084) );
	vdp_slatch g3144 (.Q(w4286), .D(S[6]), .C(w3063), .nC(w3089) );
	vdp_slatch g3145 (.Q(w4322), .D(S[6]), .C(w3064), .nC(w3090) );
	vdp_slatch g3146 (.Q(w4321), .D(S[6]), .C(w3066), .nC(w3085) );
	vdp_slatch g3147 (.Q(w4318), .D(S[1]), .C(w3059), .nC(w3084) );
	vdp_slatch g3148 (.Q(w4317), .D(S[1]), .C(w3063), .nC(w3089) );
	vdp_slatch g3149 (.Q(w4314), .D(S[1]), .C(w3064), .nC(w3090) );
	vdp_slatch g3150 (.Q(w4313), .D(S[1]), .C(w3066), .nC(w3085) );
	vdp_slatch g3151 (.Q(w4310), .D(S[5]), .C(w3059), .nC(w3084) );
	vdp_slatch g3152 (.Q(w4309), .D(S[5]), .C(w3063), .nC(w3089) );
	vdp_slatch g3153 (.Q(w4306), .D(S[5]), .C(w3064), .nC(w3090) );
	vdp_slatch g3154 (.Q(w4305), .D(S[5]), .C(w3066), .nC(w3085) );
	vdp_slatch g3155 (.Q(w4302), .D(S[0]), .C(w3059), .nC(w3084) );
	vdp_slatch g3156 (.Q(w4301), .D(S[0]), .C(w3063), .nC(w3089) );
	vdp_slatch g3157 (.Q(w4298), .D(S[0]), .C(w3064), .nC(w3090) );
	vdp_slatch g3158 (.Q(w4297), .D(S[0]), .C(w3066), .nC(w3085) );
	vdp_slatch g3159 (.Q(w4294), .D(S[4]), .C(w3059), .nC(w3084) );
	vdp_slatch g3160 (.Q(w4293), .D(S[4]), .C(w3063), .nC(w3089) );
	vdp_slatch g3161 (.Q(w4290), .D(S[4]), .C(w3064), .nC(w3090) );
	vdp_slatch g3162 (.Q(w4289), .D(S[4]), .C(w3066), .nC(w3085) );
	vdp_slatch g3163 (.Q(w4261), .D(w4263), .C(w3046), .nC(w3086) );
	vdp_slatch g3164 (.Q(w4260), .D(w4262), .C(w3049), .nC(w3087) );
	vdp_slatch g3165 (.Q(w4265), .D(w4267), .C(w3054), .nC(w3088) );
	vdp_slatch g3166 (.Q(w4264), .D(w4266), .C(w3051), .nC(w3056) );
	vdp_slatch g3167 (.Q(w4269), .D(w4271), .C(w3046), .nC(w3086) );
	vdp_slatch g3168 (.Q(w4268), .D(w4270), .C(w3049), .nC(w3087) );
	vdp_slatch g3169 (.Q(w4273), .D(w4275), .C(w3054), .nC(w3088) );
	vdp_slatch g3170 (.Q(w4272), .D(w4274), .C(w3051), .nC(w3056) );
	vdp_slatch g3171 (.Q(w4277), .D(w4279), .C(w3046), .nC(w3086) );
	vdp_slatch g3172 (.Q(w4276), .D(w4278), .C(w3049), .nC(w3087) );
	vdp_slatch g3173 (.Q(w4387), .D(w4283), .C(w3054), .nC(w3088) );
	vdp_slatch g3174 (.Q(w4281), .D(w4282), .C(w3051), .nC(w3056) );
	vdp_slatch g3175 (.Q(w4280), .D(w4285), .C(w3046), .nC(w3086) );
	vdp_slatch g3176 (.Q(w4284), .D(w4286), .C(w3049), .nC(w3087) );
	vdp_slatch g3177 (.Q(w4320), .D(w4322), .C(w3054), .nC(w3088) );
	vdp_slatch g3178 (.Q(w4319), .D(w4321), .C(w3051), .nC(w3056) );
	vdp_slatch g3179 (.Q(w4316), .D(w4318), .C(w3046), .nC(w3086) );
	vdp_slatch g3180 (.Q(w4315), .D(w4317), .C(w3049), .nC(w3087) );
	vdp_slatch g3181 (.Q(w4312), .D(w4314), .C(w3054), .nC(w3088) );
	vdp_slatch g3182 (.Q(w4311), .D(w4313), .C(w3051), .nC(w3056) );
	vdp_slatch g3183 (.Q(w4308), .D(w4310), .C(w3046), .nC(w3086) );
	vdp_slatch g3184 (.Q(w4307), .D(w4309), .C(w3049), .nC(w3087) );
	vdp_slatch g3185 (.Q(w4304), .D(w4306), .C(w3054), .nC(w3088) );
	vdp_slatch g3186 (.Q(w4303), .D(w4305), .C(w3051), .nC(w3056) );
	vdp_slatch g3187 (.D(w4302), .Q(w4300), .C(w3046), .nC(w3086) );
	vdp_slatch g3188 (.Q(w4299), .D(w4301), .C(w3049), .nC(w3087) );
	vdp_slatch g3189 (.Q(w4296), .D(w4298), .C(w3054), .nC(w3088) );
	vdp_slatch g3190 (.Q(w4295), .D(w4297), .C(w3051), .nC(w3056) );
	vdp_slatch g3191 (.Q(w4292), .D(w4294), .C(w3046), .nC(w3086) );
	vdp_slatch g3192 (.Q(w4291), .D(w4293), .C(w3049), .nC(w3087) );
	vdp_slatch g3193 (.Q(w4288), .D(w4290), .C(w3054), .nC(w3088) );
	vdp_slatch g3194 (.Q(w4287), .D(w4289), .C(w3051), .nC(w3056) );
	vdp_slatch g3195 (.Q(w3367), .D(w4261), .C(w3047), .nC(w3048) );
	vdp_slatch g3196 (.Q(w3366), .D(w4260), .C(w3055), .nC(w3050) );
	vdp_slatch g3197 (.Q(w3354), .D(w4265), .C(w3052), .nC(w3053) );
	vdp_slatch g3198 (.Q(w3352), .D(w4264), .C(w3045), .nC(w3044) );
	vdp_slatch g3199 (.Q(w3365), .D(w4269), .C(w3047), .nC(w3048) );
	vdp_slatch g3200 (.Q(w3364), .D(w4268), .C(w3055), .nC(w3050) );
	vdp_slatch g3201 (.D(w4273), .C(w3052), .nC(w3053), .Q(w3363) );
	vdp_slatch g3202 (.Q(w3351), .D(w4272), .C(w3045), .nC(w3044) );
	vdp_slatch g3203 (.Q(w3362), .D(w4277), .C(w3047), .nC(w3048) );
	vdp_slatch g3204 (.Q(w3361), .D(w4276), .C(w3055), .nC(w3050) );
	vdp_slatch g3205 (.Q(w3360), .D(w4387), .C(w3052), .nC(w3053) );
	vdp_slatch g3206 (.Q(w3359), .D(w4281), .C(w3045), .nC(w3044) );
	vdp_slatch g3207 (.Q(w3358), .D(w4280), .C(w3047), .nC(w3048) );
	vdp_slatch g3208 (.Q(w3357), .D(w4284), .C(w3055), .nC(w3050) );
	vdp_slatch g3209 (.Q(w3356), .D(w4320), .C(w3052), .nC(w3053) );
	vdp_slatch g3210 (.Q(w3355), .D(w4319), .C(w3045), .nC(w3044) );
	vdp_slatch g3211 (.Q(w3347), .D(w4316), .C(w3047), .nC(w3048) );
	vdp_slatch g3212 (.Q(w3393), .D(w4315), .C(w3055), .nC(w3050) );
	vdp_slatch g3213 (.Q(w3348), .D(w4312), .C(w3052), .nC(w3053) );
	vdp_slatch g3214 (.Q(w3349), .D(w4311), .C(w3045), .nC(w3044) );
	vdp_slatch g3215 (.Q(w3397), .D(w4308), .C(w3047), .nC(w3048) );
	vdp_slatch g3216 (.Q(w3406), .D(w4307), .C(w3055), .nC(w3050) );
	vdp_slatch g3217 (.Q(w3398), .D(w4304), .C(w3052), .nC(w3053) );
	vdp_slatch g3218 (.Q(w3405), .D(w4303), .nC(w3044), .C(w3045) );
	vdp_slatch g3219 (.Q(w3404), .D(w4300), .C(w3047), .nC(w3048) );
	vdp_slatch g3220 (.Q(w3403), .D(w4299), .C(w3055), .nC(w3050) );
	vdp_slatch g3221 (.Q(w3399), .D(w4296), .C(w3052), .nC(w3053) );
	vdp_slatch g3222 (.Q(w3402), .D(w4295), .C(w3045), .nC(w3044) );
	vdp_slatch g3223 (.Q(w3401), .D(w4292), .C(w3047), .nC(w3048) );
	vdp_slatch g3224 (.Q(w3400), .D(w4291), .C(w3055), .nC(w3050) );
	vdp_slatch g3225 (.Q(w3353), .D(w4288), .C(w3052), .nC(w3053) );
	vdp_slatch g3226 (.Q(w3350), .D(w4287), .C(w3045), .nC(w3044) );
	vdp_slatch g3227 (.Q(w3385), .D(w4326), .nC(w3447), .C(w3446) );
	vdp_slatch g3228 (.Q(w3494), .D(w4325), .nC(w3450), .C(w3451) );
	vdp_slatch g3229 (.Q(w3387), .D(w4330), .nC(w3449), .C(w3448) );
	vdp_slatch g3230 (.Q(w3386), .D(w4329), .nC(w3453), .C(w3452) );
	vdp_slatch g3231 (.Q(w3493), .D(w4334), .nC(w3447), .C(w3446) );
	vdp_slatch g3232 (.Q(w3497), .D(w4333), .nC(w3450), .C(w3451) );
	vdp_slatch g3233 (.Q(w3496), .D(w4338), .nC(w3449), .C(w3448) );
	vdp_slatch g3234 (.Q(w3495), .D(w4337), .nC(w3453), .C(w3452) );
	vdp_slatch g3235 (.Q(w3388), .D(w4342), .nC(w3447), .C(w3446) );
	vdp_slatch g3236 (.Q(w3498), .D(w4341), .nC(w3450), .C(w3451) );
	vdp_slatch g3237 (.Q(w3492), .D(w4346), .nC(w3449), .C(w3448) );
	vdp_slatch g3238 (.Q(w3499), .D(w4345), .nC(w3453), .C(w3452) );
	vdp_slatch g3239 (.Q(w3500), .D(w4350), .nC(w3447), .C(w3446) );
	vdp_slatch g3240 (.Q(w3501), .D(w4349), .nC(w3450), .C(w3451) );
	vdp_slatch g3241 (.Q(w3389), .D(w4354), .nC(w3449), .C(w3448) );
	vdp_slatch g3242 (.Q(w3390), .D(w4353), .nC(w3453), .C(w3452) );
	vdp_slatch g3243 (.Q(w3484), .D(w4358), .nC(w3447), .C(w3446) );
	vdp_slatch g3244 (.Q(w3485), .D(w4357), .nC(w3450), .C(w3451) );
	vdp_slatch g3245 (.Q(w3486), .D(w4362), .nC(w3449), .C(w3448) );
	vdp_slatch g3246 (.Q(w3487), .D(w4361), .nC(w3453), .C(w3452) );
	vdp_slatch g3247 (.Q(w3488), .D(w4366), .nC(w3447), .C(w3446) );
	vdp_slatch g3248 (.Q(w3489), .D(w4365), .nC(w3450), .C(w3451) );
	vdp_slatch g3249 (.Q(w3490), .D(w4370), .nC(w3449), .C(w3448) );
	vdp_slatch g3250 (.Q(w3491), .D(w4369), .nC(w3453), .C(w3452) );
	vdp_slatch g3251 (.Q(w3483), .D(w4374), .nC(w3447), .C(w3446) );
	vdp_slatch g3252 (.Q(w3482), .D(w4373), .nC(w3450), .C(w3451) );
	vdp_slatch g3253 (.Q(w3481), .D(w4378), .nC(w3449), .C(w3448) );
	vdp_slatch g3254 (.Q(w3480), .D(w4377), .nC(w3453), .C(w3452) );
	vdp_slatch g3255 (.Q(w3479), .D(w4382), .nC(w3447), .C(w3446) );
	vdp_slatch g3256 (.Q(w3478), .D(w4381), .nC(w3450), .C(w3451) );
	vdp_slatch g3257 (.Q(w3476), .D(w4386), .nC(w3449), .C(w3448) );
	vdp_slatch g3258 (.Q(w3477), .D(w4385), .nC(w3453), .C(w3452) );
	vdp_slatch g3259 (.Q(w4326), .D(w4324), .C(w3411), .nC(w3445) );
	vdp_slatch g3260 (.Q(w4325), .D(w4323), .C(w3437), .nC(w3439) );
	vdp_slatch g3261 (.Q(w4330), .D(w4328), .C(w3412), .nC(w3440) );
	vdp_slatch g3262 (.Q(w4329), .D(w4327), .C(w3444), .nC(w3443) );
	vdp_slatch g3263 (.Q(w4334), .D(w4332), .C(w3411), .nC(w3445) );
	vdp_slatch g3264 (.Q(w4333), .D(w4331), .C(w3437), .nC(w3439) );
	vdp_slatch g3265 (.Q(w4338), .D(w4336), .C(w3412), .nC(w3440) );
	vdp_slatch g3266 (.Q(w4337), .D(w4335), .C(w3444), .nC(w3443) );
	vdp_slatch g3267 (.Q(w4342), .D(w4340), .C(w3411), .nC(w3445) );
	vdp_slatch g3268 (.Q(w4341), .D(w4339), .C(w3437), .nC(w3439) );
	vdp_slatch g3269 (.Q(w4346), .D(w4344), .C(w3412), .nC(w3440) );
	vdp_slatch g3270 (.Q(w4345), .D(w4343), .C(w3444), .nC(w3443) );
	vdp_slatch g3271 (.Q(w4350), .D(w4348), .C(w3411), .nC(w3445) );
	vdp_slatch g3272 (.Q(w4349), .D(w4347), .C(w3437), .nC(w3439) );
	vdp_slatch g3273 (.Q(w4354), .D(w4352), .C(w3412), .nC(w3440) );
	vdp_slatch g3274 (.Q(w4353), .D(w4351), .C(w3444), .nC(w3443) );
	vdp_slatch g3275 (.Q(w4358), .D(w4356), .C(w3411), .nC(w3445) );
	vdp_slatch g3276 (.Q(w4357), .D(w4355), .C(w3437), .nC(w3439) );
	vdp_slatch g3277 (.Q(w4362), .D(w4360), .C(w3412), .nC(w3440) );
	vdp_slatch g3278 (.Q(w4361), .D(w4359), .C(w3444), .nC(w3443) );
	vdp_slatch g3279 (.Q(w4366), .D(w4364), .C(w3411), .nC(w3445) );
	vdp_slatch g3280 (.Q(w4365), .D(w4363), .C(w3437), .nC(w3439) );
	vdp_slatch g3281 (.Q(w4370), .D(w4368), .C(w3412), .nC(w3440) );
	vdp_slatch g3282 (.Q(w4369), .D(w4367), .C(w3444), .nC(w3443) );
	vdp_slatch g3283 (.Q(w4374), .D(w4372), .C(w3411), .nC(w3445) );
	vdp_slatch g3284 (.Q(w4373), .D(w4371), .C(w3437), .nC(w3439) );
	vdp_slatch g3285 (.Q(w4378), .D(w4376), .C(w3412), .nC(w3440) );
	vdp_slatch g3286 (.Q(w4377), .D(w4375), .C(w3444), .nC(w3443) );
	vdp_slatch g3287 (.Q(w4382), .D(w4380), .C(w3411), .nC(w3445) );
	vdp_slatch g3288 (.Q(w4381), .D(w4379), .C(w3437), .nC(w3439) );
	vdp_slatch g3289 (.Q(w4386), .D(w4384), .C(w3412), .nC(w3440) );
	vdp_slatch g3290 (.Q(w4385), .D(w4383), .C(w3444), .nC(w3443) );
	vdp_slatch g3291 (.Q(w4324), .D(S[3]), .nC(w3438), .C(w3466) );
	vdp_slatch g3292 (.Q(w4323), .D(S[3]), .nC(w3454), .C(w3467) );
	vdp_slatch g3293 (.Q(w4328), .D(S[3]), .nC(w3441), .C(w3465) );
	vdp_slatch g3294 (.Q(w4327), .D(S[3]), .nC(w3442), .C(w3464) );
	vdp_slatch g3295 (.Q(w4332), .D(S[7]), .nC(w3438), .C(w3466) );
	vdp_slatch g3296 (.Q(w4331), .D(S[7]), .nC(w3454), .C(w3467) );
	vdp_slatch g3297 (.Q(w4336), .D(S[7]), .nC(w3441), .C(w3465) );
	vdp_slatch g3298 (.Q(w4335), .D(S[7]), .nC(w3442), .C(w3464) );
	vdp_slatch g3299 (.Q(w4340), .D(S[2]), .nC(w3438), .C(w3466) );
	vdp_slatch g3300 (.Q(w4339), .D(S[2]), .nC(w3454), .C(w3467) );
	vdp_slatch g3301 (.Q(w4344), .D(S[2]), .nC(w3441), .C(w3465) );
	vdp_slatch g3302 (.Q(w4343), .D(S[2]), .nC(w3442), .C(w3464) );
	vdp_slatch g3303 (.Q(w4348), .D(S[6]), .nC(w3438), .C(w3466) );
	vdp_slatch g3304 (.Q(w4347), .D(S[6]), .nC(w3454), .C(w3467) );
	vdp_slatch g3305 (.Q(w4352), .D(S[6]), .nC(w3441), .C(w3465) );
	vdp_slatch g3306 (.Q(w4351), .D(S[6]), .nC(w3442), .C(w3464) );
	vdp_slatch g3307 (.Q(w4356), .D(S[1]), .nC(w3438), .C(w3466) );
	vdp_slatch g3308 (.Q(w4355), .D(S[1]), .nC(w3454), .C(w3467) );
	vdp_slatch g3309 (.Q(w4360), .D(S[1]), .nC(w3441), .C(w3465) );
	vdp_slatch g3310 (.Q(w4359), .D(S[1]), .nC(w3442), .C(w3464) );
	vdp_slatch g3311 (.Q(w4364), .D(S[5]), .nC(w3438), .C(w3466) );
	vdp_slatch g3312 (.Q(w4363), .D(S[5]), .nC(w3454), .C(w3467) );
	vdp_slatch g3313 (.Q(w4368), .D(S[5]), .nC(w3441), .C(w3465) );
	vdp_slatch g3314 (.Q(w4367), .D(S[5]), .nC(w3442), .C(w3464) );
	vdp_slatch g3315 (.Q(w4372), .D(S[0]), .nC(w3438), .C(w3466) );
	vdp_slatch g3316 (.Q(w4371), .D(S[0]), .nC(w3454), .C(w3467) );
	vdp_slatch g3317 (.Q(w4376), .D(S[0]), .nC(w3441), .C(w3465) );
	vdp_slatch g3318 (.Q(w4375), .D(S[0]), .nC(w3442), .C(w3464) );
	vdp_slatch g3319 (.Q(w4380), .D(S[4]), .nC(w3438), .C(w3466) );
	vdp_slatch g3320 (.Q(w4379), .D(S[4]), .nC(w3454), .C(w3467) );
	vdp_slatch g3321 (.Q(w4384), .D(S[4]), .nC(w3441), .C(w3465) );
	vdp_slatch g3322 (.Q(w4383), .D(S[4]), .nC(w3442), .C(w3464) );
	vdp_aon2*8 g3323 (.Z(w4022), .A1(w3183), .B1(w3182), .C1(w3181), .D2(w3180), .A2(w3227), .B2(w3228), .C2(w3233), .D1(w3232), .E2(w3230), .F1(w3231), .E1(w3179), .F2(w3178), .G1(w3177), .H2(w3176), .G2(w3235), .H1(w3225) );
	vdp_aon2*8 g3324 (.Z(w3207), .A1(w3301), .B1(w3228), .C1(w3303), .D2(w3232), .A2(w3227), .B2(w3302), .C2(w3233), .D1(w3304), .E2(w3230), .F1(w3231), .E1(w3305), .F2(w3306), .G1(w3312), .H2(w3313), .G2(w3235), .H1(w3225) );
	vdp_aon2*8 g3325 (.Z(w3210), .A1(w3175), .B1(w3188), .C1(w3192), .D2(w3191), .A2(w3227), .B2(w3228), .C2(w3233), .D1(w3232), .E2(w3230), .F1(w3231), .E1(w3190), .F2(w3186), .G1(w3187), .H2(w3189), .G2(w3235), .H1(w3225) );
	vdp_aon2*8 g3326 (.Z(w3211), .A1(w3314), .B1(w3228), .C1(w3316), .D2(w3232), .A2(w3227), .B2(w3315), .C2(w3233), .D1(w3311), .E2(w3230), .F1(w3231), .E1(w3317), .F2(w3318), .G1(w3319), .H2(w3320), .G2(w3235), .H1(w3225) );
	vdp_aon2*8 g3327 (.Z(w3209), .A1(w3245), .B1(w3228), .C1(w3247), .D2(w3248), .A2(w3227), .B2(w4023), .C2(w3233), .D1(w3232), .E2(w3230), .F1(w3231), .E1(w3321), .F2(w3246), .G1(w3226), .H2(w3249), .G2(w3235), .H1(w3225) );
	vdp_aon2*8 g3328 (.Z(w3212), .A1(w3252), .B1(w3228), .C1(w3259), .D2(w3258), .A2(w3227), .B2(w3260), .C2(w3233), .D1(w3232), .E2(w3230), .F1(w3231), .E1(w3256), .F2(w3250), .G1(w3257), .G2(w3235), .H1(w3225), .H2(w3251) );
	vdp_aon2*8 g3329 (.Z(w3208), .A1(w3193), .B1(w3194), .C1(w3196), .D2(w3195), .A2(w3227), .B2(w3228), .C2(w3233), .D1(w3232), .E2(w3230), .F1(w3231), .E1(w3237), .F2(w3238), .G1(w3234), .H2(w3229), .G2(w3235), .H1(w3225) );
	vdp_aon2*8 g3330 (.Z(w3213), .A1(w3241), .B1(w3240), .C1(w3239), .D2(w3236), .A2(w3227), .B2(w3228), .C2(w3233), .D1(w3232), .E2(w3230), .F1(w3231), .E1(w3222), .F2(w3221), .G1(w3223), .H2(w3224), .G2(w3235), .H1(w3225) );
	vdp_aon2*8 g3331 (.A1(w3367), .B1(w3366), .C1(w3354), .D2(w3352), .A2(w3384), .B2(w3383), .C2(w3382), .D1(w3381), .E2(w3380), .F1(w3379), .E1(w3365), .F2(w3364), .G1(w3363), .H2(w3351), .G2(w3377), .H1(w3378), .Z(w3396) );
	vdp_aon2*8 g3332 (.Z(w3424), .A1(w3362), .B1(w3361), .C1(w3360), .D2(w3359), .A2(w3384), .B2(w3383), .C2(w3382), .D1(w3381), .E2(w3380), .F1(w3379), .E1(w3358), .F2(w3357), .G1(w3356), .H2(w3355), .G2(w3377), .H1(w3378) );
	vdp_aon2*8 g3333 (.Z(w3395), .A1(w3354), .B1(w3363), .C1(w3360), .D2(w3356), .A2(w3379), .B2(w3378), .C2(w3383), .D1(w3381), .E2(w3380), .F1(w3377), .E1(w3348), .F2(w3398), .G1(w3399), .H2(w3353), .G2(w3384), .H1(w3382) );
	vdp_aon2*8 g3334 (.Z(w3427), .A1(w3347), .B1(w3393), .C1(w3348), .D2(w3349), .A2(w3384), .B2(w3383), .C2(w3382), .D1(w3381), .E2(w3380), .F1(w3379), .E1(w3397), .F2(w3406), .G1(w3398), .H2(w3405), .G2(w3377), .H1(w3378) );
	vdp_aon2*8 g3335 (.Z(w3394), .A1(w3404), .B1(w3403), .C1(w3399), .D2(w3402), .A2(w3384), .B2(w3383), .C2(w3382), .D1(w3381), .E2(w3380), .F1(w3379), .E1(w3401), .F2(w3400), .G1(w3353), .H2(w3350), .G2(w3377), .H1(w3378) );
	vdp_aon2*8 g3336 (.Z(w3429), .A1(w3483), .B1(w3383), .C1(w3481), .D2(w3381), .A2(w3384), .B2(w3482), .C2(w3382), .D1(w3480), .E2(w3380), .F1(w3379), .E1(w3479), .F2(w3478), .G1(w3476), .H2(w3477), .G2(w3377), .H1(w3378) );
	vdp_aon2*8 g3337 (.Z(w3430), .A1(w3484), .B1(w3383), .C1(w3486), .D2(w3381), .A2(w3384), .B2(w3485), .C2(w3382), .D1(w3487), .E2(w3380), .F1(w3379), .E1(w3488), .F2(w3489), .G1(w3490), .H2(w3491), .G2(w3377), .H1(w3378) );
	vdp_aon2*8 g3338 (.Z(w3428), .A1(w3352), .B1(w3351), .C1(w3359), .D2(w3355), .A2(w3379), .B2(w3378), .C2(w3383), .D1(w3381), .E2(w3380), .F1(w3377), .E1(w3349), .F2(w3405), .G1(w3402), .H2(w3350), .G2(w3384), .H1(w3382) );
	vdp_aon2*8 g3339 (.Z(w3423), .A1(w3386), .B1(w3378), .C1(w3499), .D2(w3381), .A2(w3379), .B2(w3495), .C2(w3383), .D1(w3390), .E2(w3380), .F1(w3377), .E1(w3487), .F2(w3491), .G1(w3480), .H2(w3477), .G2(w3384), .H1(w3382) );
	vdp_aon2*8 g3340 (.Z(w3426), .A1(w3387), .B1(w3378), .C1(w3492), .D2(w3381), .A2(w3379), .B2(w3496), .C2(w3383), .D1(w3389), .E2(w3380), .F1(w3377), .E1(w3486), .F2(w3490), .G1(w3481), .H2(w3476), .G2(w3384), .H1(w3382) );
	vdp_aon2*8 g3341 (.Z(w3425), .A1(w3388), .B1(w3383), .C1(w3492), .D2(w3381), .A2(w3384), .B2(w3498), .C2(w3382), .D1(w3499), .E2(w3380), .F1(w3379), .E1(w3500), .F2(w3501), .G1(w3389), .H2(w3390), .G2(w3377), .H1(w3378) );
	vdp_aon2*8 g3342 (.A1(w3385), .B1(w3383), .C1(w3387), .D2(w3381), .A2(w3384), .B2(w3494), .C2(w3382), .D1(w3386), .E2(w3380), .F1(w3379), .E1(w3493), .F2(w3497), .G1(w3496), .H2(w3495), .G2(w3377), .H1(w3378), .Z(w3431) );
	vdp_sr_bit g3343 (.Q(w3374), .D(w3529), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3344 (.Q(w3529), .D(w3433), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3345 (.Q(w3434), .D(w3530), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3346 (.Q(w3530), .D(w3436), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3347 (.Q(w3435), .D(w3410), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3348 (.Q(w4053), .D(w3435), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3349 (.Q(w3514), .D(w3432), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3350 (.Q(w3409), .D(w3514), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3351 (.Q(w4055), .D(w3419), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3352 (.Q(w3408), .D(w4055), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3353 (.Q(w3407), .D(w3375), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3354 (.Q(w3375), .D(w3418), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3355 (.Q(w2823), .D(w3420), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3356 (.Q(w3515), .D(w2823), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3357 (.Q(w3199), .D(w3217), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3358 (.Q(w3201), .D(w3199), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3359 (.Q(w3204), .D(w3200), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3360 (.Q(w3200), .D(w3216), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3361 (.Q(w3215), .D(w3197), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3362 (.Q(w3197), .D(w3218), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3363 (.Q(w3198), .D(w3214), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3364 (.Q(w3206), .D(w3198), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3365 (.Q(w3284), .D(w2822), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3366 (.Q(w2822), .D(w3269), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3367 (.Q(w4034), .D(w3219), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3368 (.Q(w3205), .D(w4034), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3369 (.Q(w4033), .D(w3270), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3370 (.Q(w3203), .D(w4033), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3371 (.Q(w3131), .D(VRAMA[1]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3372 (.Q(w3163), .D(VRAMA[2]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3373 (.Q(w3165), .D(VRAMA[3]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3374 (.Q(w3166), .D(VRAMA[4]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3375 (.Q(w3167), .D(VRAMA[5]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3376 (.Q(w3168), .D(VRAMA[6]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3377 (.Q(w4031), .D(w3154), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3378 (.Q(w3516), .D(w4031), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3379 (.Q(w3153), .D(w3517), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3380 (.Q(w3517), .D(w3516), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_dlatch_inv g3381 (.nQ(w3154), .D(w3119), .C(DCLK1), .nC(nDCLK1) );
	vdp_slatch g3382 (.Q(w3278), .D(w4388), .C(w3271), .nC(w3032) );
	vdp_slatch g3383 (.Q(w3277), .D(w4389), .C(w3271), .nC(w3032) );
	vdp_slatch g3384 (.Q(w3276), .D(w4390), .C(w3271), .nC(w3032) );
	vdp_slatch g3385 (.Q(w3275), .D(w4391), .C(w3271), .nC(w3032) );
	vdp_slatch g3386 (.Q(w3274), .D(w4392), .C(w3271), .nC(w3032) );
	vdp_slatch g3387 (.Q(w3273), .D(w4393), .C(w3271), .nC(w3032) );
	vdp_slatch g3388 (.Q(w3272), .D(w4395), .C(w3271), .nC(w3032) );
	vdp_slatch g3389 (.Q(w3033), .D(w4394), .C(w3271), .nC(w3032) );
	vdp_slatch g3390 (.Q(w4388), .D(w3100), .C(w3292), .nC(w3323) );
	vdp_slatch g3391 (.Q(w4389), .D(w3074), .C(w3292), .nC(w3323) );
	vdp_slatch g3392 (.Q(w4390), .D(w3076), .C(w3292), .nC(w3323) );
	vdp_slatch g3393 (.Q(w4391), .D(w3077), .C(w3292), .nC(w3323) );
	vdp_slatch g3394 (.Q(w4392), .D(w3078), .C(w3292), .nC(w3323) );
	vdp_slatch g3395 (.Q(w4393), .D(w3101), .C(w3292), .nC(w3323) );
	vdp_slatch g3396 (.Q(w4395), .D(w3105), .C(w3292), .nC(w3323) );
	vdp_slatch g3397 (.Q(w4394), .D(w3104), .C(w3292), .nC(w3323) );
	vdp_slatch g3398 (.Q(w4396), .D(w3040), .C(w3042), .nC(w3041) );
	vdp_slatch g3399 (.Q(w4397), .D(w3073), .C(w3042), .nC(w3041) );
	vdp_slatch g3400 (.Q(w4398), .D(w3039), .C(w3042), .nC(w3041) );
	vdp_slatch g3401 (.Q(w4399), .D(w4085), .C(w3042), .nC(w3041) );
	vdp_slatch g3402 (.Q(w4400), .D(w3525), .C(w3042), .nC(w3041) );
	vdp_slatch g3403 (.Q(w4401), .D(w3080), .C(w3042), .nC(w3041) );
	vdp_slatch g3404 (.Q(w4402), .D(w3036), .C(w3042), .nC(w3041) );
	vdp_slatch g3405 (.Q(w4403), .D(w3081), .C(w3042), .nC(w3041) );
	vdp_slatch g3406 (.Q(w3332), .D(w4396), .C(w3043), .nC(w3325) );
	vdp_slatch g3407 (.Q(w3331), .D(w4397), .C(w3043), .nC(w3325) );
	vdp_slatch g3408 (.Q(w3330), .D(w4398), .C(w3043), .nC(w3325) );
	vdp_slatch g3409 (.Q(w3329), .D(w4399), .C(w3043), .nC(w3325) );
	vdp_slatch g3410 (.Q(w3328), .D(w4400), .C(w3043), .nC(w3325) );
	vdp_slatch g3411 (.Q(w3327), .D(w4401), .C(w3043), .nC(w3325) );
	vdp_slatch g3412 (.Q(w3326), .D(w4402), .C(w3043), .nC(w3325) );
	vdp_slatch g3413 (.Q(w4429), .D(w4403), .C(w3043), .nC(w3325) );
	vdp_slatch g3414 (.Q(w3468), .D(w3462), .C(w3151), .nC(w3459) );
	vdp_slatch g3415 (.Q(w3461), .D(w3158), .C(w3151), .nC(w3459) );
	vdp_slatch g3416 (.Q(w3864), .D(w3460), .C(w3151), .nC(w3459) );
	vdp_slatch g3417 (.Q(w3455), .D(w3458), .C(w3151), .nC(w3459) );
	vdp_slatch g3418 (.Q(w3040), .D(w3100), .C(w3103), .nC(w3102) );
	vdp_slatch g3419 (.Q(w3073), .D(w3074), .C(w3103), .nC(w3102) );
	vdp_slatch g3420 (.Q(w3039), .D(w3076), .C(w3103), .nC(w3102) );
	vdp_slatch g3421 (.Q(w4085), .D(w3077), .C(w3103), .nC(w3102) );
	vdp_slatch g3422 (.Q(w3525), .D(w3078), .C(w3103), .nC(w3102) );
	vdp_slatch g3423 (.Q(w3080), .D(w3101), .C(w3103), .nC(w3102) );
	vdp_slatch g3424 (.Q(w3036), .D(w3105), .C(w3103), .nC(w3102) );
	vdp_slatch g3425 (.Q(w3081), .D(w3104), .C(w3103), .nC(w3102) );
	vdp_cnt_bit_load g3426 (.D(w3460), .nL(w3123), .L(w3120), .R(1'b0), .Q(w3122), .CI(w3521), .CO(w3522), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3427 (.D(w3158), .nL(w3123), .L(w3120), .R(1'b0), .Q(w4020), .CI(w3522), .CO(w3523), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3428 (.D(w3124), .nL(w3123), .L(w3120), .R(1'b0), .Q(w3108), .CI(w3523), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3429 (.CO(w3521), .CI(1'b1), .D(w3458), .nL(w3123), .L(w3120), .R(1'b0), .Q(w3118), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3430 (.CO(w3520), .CI(1'b1), .D(w3455), .nL(w3457), .L(w3150), .R(1'b0), .Q(w3475), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3431 (.CO(w3519), .CI(w3520), .D(w3864), .nL(w3457), .L(w3150), .R(1'b0), .Q(w3421), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3432 (.CO(w3518), .CI(w3519), .D(w3461), .nL(w3457), .L(w3150), .R(1'b0), .Q(w3463), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g3433 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .CI(w3518), .D(w3468), .nL(w3457), .L(w3150), .R(1'b0), .Q(w3373) );
	vdp_xor g3434 (.Z(w3261), .B(w4020), .A(w3117) );
	vdp_xor g3435 (.B(w3122), .A(w3117), .Z(w3109) );
	vdp_xor g3436 (.Z(w3264), .B(w3118), .A(w3117) );
	vdp_sr_bit g3437 (.Q(w3116), .D(w4029), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3438 (.Q(w4028), .D(w3116), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3439 (.Q(w3283), .D(w4028), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3440 (.Q(w4037), .D(w3524), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3441 (.Q(w3524), .D(w4038), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3442 (.Q(w4038), .D(w4039), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3443 (.Q(w3038), .D(w3037), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3444 (.Q(w3037), .D(w3035), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3445 (.Q(w3035), .D(w3034), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3446 (.Q(w4041), .D(w4042), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3447 (.Q(w4008), .D(w4041), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3448 (.Q(w4040), .D(w4008), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3449 (.Q(w4045), .D(w4044), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3450 (.Q(w4046), .D(w4045), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3451 (.Q(w4043), .D(w4046), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3452 (.Q(w3130), .D(w4043), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3453 (.Q(w4128), .D(w4129), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3454 (.Q(w4129), .D(w4048), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_xor g3455 (.Z(w3335), .A(w3417), .B(w3463) );
	vdp_xor g3456 (.Z(w3340), .A(w3417), .B(w3474) );
	vdp_xor g3457 (.Z(w3334), .A(w3417), .B(w3475) );
	vdp_dlatch_inv g3458 (.nQ(w4027), .D(w4026), .C(HCLK1), .nC(nHCLK1) );
	vdp_dlatch_inv g3459 (.nQ(w3034), .D(w3079), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g3460 (.nQ(w4042), .D(w3030), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g3461 (.nQ(w3473), .D(w4049), .nC(nHCLK1), .C(HCLK1) );
	vdp_xor g3462 (.Z(w3474), .A(w3421), .B(M5) );
	vdp_sr_bit g3463 (.Q(w3527), .D(w3422), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_dlatch_inv g3464 (.nQ(w4044), .D(w3128), .nC(nDCLK1), .C(DCLK1) );
	vdp_comp_strong g3465 (.Z(w3047), .nZ(w3048), .A(w3324) );
	vdp_comp_strong g3466 (.Z(w3055), .nZ(w3050), .A(w3324) );
	vdp_comp_strong g3467 (.Z(w3052), .nZ(w3053), .A(w3324) );
	vdp_comp_strong g3468 (.Z(w3045), .nZ(w3044), .A(w3324) );
	vdp_comp_strong g3469 (.Z(w3046), .nZ(w3086), .A(w3082) );
	vdp_comp_strong g3470 (.Z(w3049), .nZ(w3087), .A(w3082) );
	vdp_comp_strong g3471 (.Z(w3054), .nZ(w3088), .A(w3082) );
	vdp_comp_strong g3472 (.Z(w3051), .nZ(w3056), .A(w3082) );
	vdp_comp_strong g3473 (.Z(w3059), .nZ(w3084), .A(w3083) );
	vdp_comp_strong g3474 (.Z(w3063), .nZ(w3089), .A(w3392) );
	vdp_comp_strong g3475 (.Z(w3064), .nZ(w3090), .A(w3391) );
	vdp_comp_strong g3476 (.Z(w3066), .nZ(w3085), .A(w3075) );
	vdp_comp_strong g3477 (.Z(w3058), .nZ(w3092), .A(w4036) );
	vdp_comp_strong g3478 (.Z(w3062), .nZ(w3096), .A(w3097) );
	vdp_comp_strong g3479 (.Z(w3065), .nZ(w3093), .A(w3099) );
	vdp_comp_strong g3480 (.Z(w3067), .nZ(w3091), .A(w3098) );
	vdp_comp_strong g3481 (.Z(w3291), .nZ(w3285), .A(w3031) );
	vdp_comp_strong g3482 (.Z(w3106), .nZ(w3286), .A(w3031) );
	vdp_comp_strong g3483 (.Z(w3293), .nZ(w3094), .A(w3031) );
	vdp_comp_strong g3484 (.Z(w3294), .nZ(w3095), .A(w3031) );
	vdp_comp_strong g3485 (.Z(w3298), .nZ(w3299), .A(w3107) );
	vdp_comp_strong g3486 (.Z(w3297), .nZ(w3307), .A(w3107) );
	vdp_comp_strong g3487 (.Z(w3296), .nZ(w3308), .A(w3107) );
	vdp_comp_strong g3488 (.Z(w3295), .nZ(w3300), .A(w3107) );
	vdp_comp_strong g3489 (.Z(w3148), .nZ(w3174), .A(w3107) );
	vdp_comp_strong g3490 (.Z(w3127), .nZ(w3184), .A(w3107) );
	vdp_comp_strong g3491 (.Z(w3139), .nZ(w3185), .A(w3107) );
	vdp_comp_strong g3492 (.Z(w3140), .nZ(w3114), .A(w3107) );
	vdp_comp_strong g3493 (.Z(w3126), .nZ(w3143), .A(w3031) );
	vdp_comp_strong g3494 (.Z(w3144), .nZ(w3135), .A(w3031) );
	vdp_comp_strong g3495 (.Z(w3145), .nZ(w3133), .A(w3031) );
	vdp_comp_strong g3496 (.Z(w3141), .nZ(w3142), .A(w3031) );
	vdp_comp_strong g3497 (.Z(w3156), .nZ(w3146), .A(w3157) );
	vdp_comp_strong g3498 (.Z(w3137), .nZ(w3136), .A(w3159) );
	vdp_comp_strong g3499 (.Z(w3138), .nZ(w3134), .A(w3160) );
	vdp_comp_strong g3500 (.Z(w3155), .nZ(w3147), .A(w3161) );
	vdp_comp_strong g3501 (.Z(w3466), .nZ(w3438), .A(w3281) );
	vdp_comp_strong g3502 (.Z(w3467), .nZ(w3454), .A(w3469) );
	vdp_comp_strong g3503 (.Z(w3465), .nZ(w3441), .A(w3470) );
	vdp_comp_strong g3504 (.Z(w3464), .nZ(w3442), .A(w3471) );
	vdp_comp_strong g3505 (.Z(w3411), .nZ(w3445), .A(w3082) );
	vdp_comp_strong g3506 (.Z(w3437), .nZ(w3439), .A(w3082) );
	vdp_comp_strong g3507 (.Z(w3412), .nZ(w3440), .A(w3082) );
	vdp_comp_strong g3508 (.Z(w3444), .nZ(w3443), .A(w3082) );
	vdp_comp_strong g3509 (.Z(w3446), .nZ(w3447), .A(w3324) );
	vdp_comp_strong g3510 (.Z(w3451), .nZ(w3450), .A(w3324) );
	vdp_comp_strong g3511 (.Z(w3448), .nZ(w3449), .A(w3324) );
	vdp_comp_strong g3512 (.Z(w3452), .nZ(w3453), .A(w3324) );
	vdp_not g3513 (.nZ(w3124), .A(w3462) );
	vdp_not g3514 (.nZ(w4029), .A(w3242) );
	vdp_not g3515 (.nZ(w3244), .A(w103) );
	vdp_not g3516 (.nZ(w3243), .A(w440) );
	vdp_not g3517 (.nZ(w3110), .A(w3243) );
	vdp_comp_strong g3518 (.Z(w3271), .nZ(w3032), .A(w3107) );
	vdp_comp_strong g3519 (.Z(w3292), .nZ(w3323), .A(w3031) );
	vdp_comp_strong g3520 (.Z(w3103), .nZ(w3102), .A(w3281) );
	vdp_comp_strong g3521 (.Z(w3043), .nZ(w3325), .A(w3324) );
	vdp_comp_strong g3522 (.Z(w3042), .nZ(w3041), .A(w3082) );
	vdp_comp_strong g3523 (.Z(w3151), .nZ(w3459), .A(w3527) );
	vdp_not g3524 (.nZ(w3341), .A(w3334) );
	vdp_not g3525 (.nZ(w3333), .A(w3340) );
	vdp_not g3526 (.nZ(w3344), .A(w3335) );
	vdp_nand3 g3527 (.Z(w3338), .A(w3344), .B(w3340), .C(w3334) );
	vdp_not g3528 (.nZ(w3383), .A(w3337) );
	vdp_nand3 g3529 (.Z(w3337), .A(w3335), .B(w3333), .C(w3334) );
	vdp_nand3 g3530 (.Z(w3336), .A(w3335), .B(w3340), .C(w3334) );
	vdp_nand3 g3531 (.Z(w3342), .A(w3335), .B(w3340), .C(w3341) );
	vdp_nand3 g3532 (.Z(w3339), .A(w3344), .B(w3333), .C(w3334) );
	vdp_nand3 g3533 (.Z(w3345), .A(w3344), .B(w3340), .C(w3341) );
	vdp_nand3 g3534 (.Z(w3343), .A(w3335), .B(w3333), .C(w3341) );
	vdp_nand3 g3535 (.Z(w3346), .A(w3341), .B(w3344), .C(w3333) );
	vdp_not g3536 (.nZ(w3384), .A(w3336) );
	vdp_not g3537 (.nZ(w3382), .A(w3338) );
	vdp_not g3538 (.nZ(w3381), .A(w3339) );
	vdp_not g3539 (.nZ(w3379), .A(w3343) );
	vdp_not g3540 (.nZ(w3380), .A(w3342) );
	vdp_not g3541 (.nZ(w3378), .A(w3346) );
	vdp_not g3542 (.nZ(w3377), .A(w3345) );
	vdp_not g3543 (.nZ(w3254), .A(w3264) );
	vdp_not g3544 (.nZ(w3262), .A(w3115) );
	vdp_not g3545 (.nZ(w3253), .A(w3261) );
	vdp_nand3 g3546 (.Z(w3266), .A(w3253), .B(w3115), .C(w3264) );
	vdp_not g3547 (.nZ(w3228), .A(w3268) );
	vdp_nand3 g3548 (.Z(w3268), .A(w3261), .B(w3262), .C(w3264) );
	vdp_nand3 g3549 (.Z(w3267), .A(w3261), .B(w3115), .C(w3264) );
	vdp_nand3 g3550 (.Z(w4035), .A(w3261), .B(w3115), .C(w3254) );
	vdp_nand3 g3551 (.Z(w3265), .A(w3253), .B(w3262), .C(w3264) );
	vdp_nand3 g3552 (.Z(w3263), .A(w3261), .B(w3262), .C(w3254) );
	vdp_not g3553 (.nZ(w3227), .A(w3267) );
	vdp_not g3554 (.nZ(w3233), .A(w3266) );
	vdp_not g3555 (.nZ(w3232), .A(w3265) );
	vdp_not g3556 (.nZ(w3231), .A(w3263) );
	vdp_not g3557 (.nZ(w3230), .A(w4035) );
	vdp_aon22 g3558 (.Z(w3269), .A1(w3272), .B1(w3279), .A2(w3280), .B2(w3033) );
	vdp_aon22 g3559 (.Z(w3270), .A1(w3274), .B1(w3279), .A2(w3280), .B2(w3273) );
	vdp_aon22 g3560 (.Z(w3219), .A1(w3276), .B1(w3279), .A2(w3280), .B2(w3275) );
	vdp_aon22 g3561 (.Z(w3117), .A1(w3278), .B1(w3279), .A2(w3280), .B2(w3277) );
	vdp_sr_bit g3562 (.Q(w3113), .D(w4030), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3563 (.Q(w4030), .D(w3112), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_xor g3564 (.Z(1'b1), .A(w3115), .B(w3109) );
	vdp_xor g3565 (.A(HPOS[3]), .B(w3132), .Z(w4084) );
	vdp_aon22 g3566 (.Z(w3170), .A1(w3163), .B1(w3164), .A2(w3162), .B2(w4083) );
	vdp_aon22 g3567 (.Z(w3171), .A1(w3165), .B1(w3164), .A2(w3162), .B2(w4082) );
	vdp_aon22 g3568 (.Z(w3173), .A1(w3166), .B1(w3164), .A2(w3162), .B2(w4081) );
	vdp_aon22 g3569 (.Z(w3172), .A1(w3167), .B1(w3164), .A2(w3162), .B2(w4080) );
	vdp_aon22 g3570 (.Z(w3608), .A1(w3168), .B1(w3164), .A2(w3162), .B2(w4079) );
	vdp_aon22 g3571 (.Z(w3214), .A1(w3310), .B1(w4022), .A2(w3207), .B2(w3309) );
	vdp_aon22 g3572 (.Z(w3218), .A1(w3310), .B1(w3208), .A2(w3209), .B2(w3309) );
	vdp_aon22 g3573 (.Z(w3216), .A1(w3310), .B1(w3213), .A2(w3212), .B2(w3309) );
	vdp_aon22 g3574 (.Z(w3217), .A1(w3310), .B1(w3210), .A2(w3211), .B2(w3309) );
	vdp_aon222 g3575 (.Z(w3433), .A1(w3425), .B1(w3424), .C1(w3423), .A2(w3371), .B2(w3372), .C2(w3370) );
	vdp_aon222 g3576 (.Z(w3436), .A1(w3429), .B1(w3394), .C1(w3428), .A2(w3371), .B2(w3372), .C2(w3370) );
	vdp_aon222 g3577 (.Z(w3410), .A1(w3430), .B1(w3427), .C1(w3395), .A2(w3371), .B2(w3372), .C2(w3370) );
	vdp_aon222 g3578 (.A1(w3431), .B1(w3396), .C1(w3426), .A2(w3371), .B2(w3372), .C2(w3370), .Z(w3432) );
	vdp_and5 g3579 (.Z(w3472), .A(w3422), .B(w3468), .C(w3461), .D(w3864), .E(w3455) );
	vdp_aon22 g3580 (.Z(w3419), .A1(w3328), .B1(w3528), .A2(w3149), .B2(w3327) );
	vdp_aon22 g3581 (.Z(w3418), .A1(w3330), .B1(w3528), .A2(w3149), .B2(w3329) );
	vdp_aon22 g3582 (.Z(w3417), .A1(w3332), .B1(w3528), .A2(w3149), .B2(w3331) );
	vdp_aon22 g3583 (.Z(w3420), .A1(w3326), .B1(w3528), .A2(w3149), .B2(w4429) );
	vdp_aon22 g3584 (.Z(w3129), .A1(w3414), .B1(w3153), .A2(w3130), .B2(M5) );
	vdp_and4 g3585 (.Z(w3415), .A(w3475), .B(w3421), .C(w3463), .D(w3416) );
	vdp_comp_we g3586 (.Z(w3149), .nZ(w3528), .A(w3413) );
	vdp_comp_we g3587 (.Z(w3309), .nZ(w3310), .A(w3108) );
	vdp_comp_we g3588 (.Z(w3280), .nZ(w3279), .A(w3108) );
	vdp_comp_we g3589 (.Z(w3120), .nZ(w3123), .A(w3202) );
	vdp_comp_we g3590 (.Z(w3162), .nZ(w3164), .A(w3698) );
	vdp_comp_we g3591 (.Z(w3150), .nZ(w3457), .A(w3422) );
	vdp_not g3592 (.nZ(w4050), .A(M5) );
	vdp_dlatch_inv g3593 (.nQ(w4039), .D(w3125), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g3594 (.Z(w3289), .A(DCLK2), .B(w3035) );
	vdp_and g3595 (.Z(w3290), .A(DCLK2), .B(w3034) );
	vdp_and g3596 (.Z(w3288), .A(DCLK2), .B(w3037) );
	vdp_and g3597 (.Z(w3287), .A(DCLK2), .B(w3038) );
	vdp_and g3598 (.Z(w3098), .A(w4039), .B(DCLK2) );
	vdp_and g3599 (.Z(w3099), .A(w4038), .B(DCLK2) );
	vdp_and g3600 (.Z(w3097), .A(w3524), .B(DCLK2) );
	vdp_and g3601 (.Z(w4036), .A(w4037), .B(DCLK2) );
	vdp_and g3602 (.Z(w3083), .A(DCLK2), .B(w4040) );
	vdp_and g3603 (.Z(w3392), .A(DCLK2), .B(w4008) );
	vdp_and g3604 (.Z(w3391), .A(DCLK2), .B(w4041) );
	vdp_and g3605 (.Z(w3075), .A(DCLK2), .B(w4042) );
	vdp_and g3606 (.Z(w3107), .A(w4027), .B(HCLK2) );
	vdp_and g3607 (.Z(w3282), .A(w3244), .B(w3116) );
	vdp_and g3608 (.Z(w3324), .A(w3473), .B(HCLK2) );
	vdp_or g3609 (.Z(w3416), .A(w4050), .B(w3373) );
	vdp_and g3610 (.Z(w3082), .A(w3129), .B(DCLK2) );
	vdp_and g3611 (.Z(w3471), .A(DCLK2), .B(w4044) );
	vdp_and g3612 (.Z(w3470), .A(DCLK2), .B(w4045) );
	vdp_and g3613 (.Z(w3469), .A(DCLK2), .B(w4046) );
	vdp_and g3614 (.Z(w3281), .A(DCLK2), .B(w4043) );
	vdp_and g3615 (.Z(w3413), .A(M5), .B(w3373) );
	vdp_and g3616 (.Z(w4080), .A(w44), .B(HPOS[7]) );
	vdp_and g3617 (.Z(w4079), .A(w44), .B(HPOS[8]) );
	vdp_and g3618 (.Z(w3161), .A(DCLK2), .B(w3154) );
	vdp_and g3619 (.Z(w4081), .A(w44), .B(HPOS[6]) );
	vdp_and g3620 (.Z(w3160), .A(DCLK2), .B(w4031) );
	vdp_and g3621 (.Z(w3159), .A(DCLK2), .B(w3516) );
	vdp_and g3622 (.Z(w3157), .A(DCLK2), .B(w3517) );
	vdp_and g3623 (.Z(w4082), .A(w44), .B(HPOS[5]) );
	vdp_and g3624 (.Z(w3031), .A(DCLK2), .B(w3153) );
	vdp_and g3625 (.Z(w4083), .A(w44), .B(HPOS[4]) );
	vdp_aon22 g3626 (.Z(w3169), .A1(w3131), .B1(w3164), .A2(w3162), .B2(w4084) );
	vdp_and g3627 (.nZ(w3132), .A(w44), .B(M5) );
	vdp_or4 g3628 (.Z(w2853), .D(w3197), .C(w3198), .B(w3199), .A(w3200) );
	vdp_or g3629 (.Z(w3202), .A(w92), .B(w15) );
	vdp_or g3630 (.Z(w3422), .A(w10), .B(w90) );
	vdp_or4 g3631 (.Z(w2854), .A(w3530), .B(w3529), .C(w3514), .D(w3435) );
	vdp_not g3632 (.nZ(w4048), .A(w3376) );
	vdp_not g3633 (.nZ(w3112), .A(w3220) );
	vdp_not g3634 (.nZ(w3414), .A(M5) );
	vdp_aoi21 g3635 (.Z(w3376), .A1(w105), .A2(w3110), .B(w17) );
	vdp_aoi21 g3636 (.Z(w3220), .A1(w106), .A2(w3110), .B(w11) );
	vdp_aoi21 g3637 (.Z(w3242), .A1(w103), .A2(w3110), .B(w12) );
	vdp_nand4 g3638 (.D(w3108), .C(w3118), .Z(w4026), .A(w4020), .B(w3122) );
	vdp_nand3 g3639 (.Z(w3255), .A(w3253), .B(w3115), .C(w3254) );
	vdp_not g3640 (.nZ(w3235), .A(w3255) );
	vdp_nand3 g3641 (.Z(w3322), .A(w3254), .B(w3253), .C(w3262) );
	vdp_not g3642 (.nZ(w3225), .A(w3322) );
	vdp_not g3643 (.nZ(w3372), .A(w3368) );
	vdp_not g3644 (.nZ(w3371), .A(w3369) );
	vdp_not g3645 (.nZ(w4025), .A(w3373) );
	vdp_not g3646 (.nZ(w3370), .A(M5) );
	vdp_not g3647 (.nZ(w4054), .A(PLANE_A_PRIO) );
	vdp_not g3648 (.nZ(w4032), .A(PLANE_B_PRIO) );
	vdp_bufif0 g3649 (.Z(COL[5]), .A(w3203), .nE(w4032) );
	vdp_bufif0 g3650 (.Z(COL[6]), .A(w3284), .nE(w4032) );
	vdp_bufif0 g3651 (.Z(COL[4]), .A(w3205), .nE(w4032) );
	vdp_bufif0 g3652 (.Z(COL[3]), .A(w3206), .nE(w4032) );
	vdp_bufif0 g3653 (.Z(COL[2]), .A(w3201), .nE(w4032) );
	vdp_bufif0 g3654 (.Z(COL[1]), .A(w3215), .nE(w4032) );
	vdp_bufif0 g3655 (.Z(COL[0]), .A(w3204), .nE(w4032) );
	vdp_bufif0 g3656 (.Z(COL[5]), .A(w3408), .nE(w4054) );
	vdp_bufif0 g3657 (.Z(COL[6]), .A(w3515), .nE(w4054) );
	vdp_bufif0 g3658 (.Z(COL[4]), .A(w3407), .nE(w4054) );
	vdp_bufif0 g3659 (.Z(COL[3]), .A(w3409), .nE(w4054) );
	vdp_bufif0 g3660 (.Z(COL[2]), .A(w3374), .nE(w4054) );
	vdp_bufif0 g3661 (.Z(COL[1]), .A(w4053), .nE(w4054) );
	vdp_bufif0 g3662 (.Z(COL[0]), .A(w3434), .nE(w4054) );
	vdp_nand g3663 (.Z(w3119), .B(HCLK1), .A(w3113) );
	vdp_nand g3664 (.Z(w3125), .B(HCLK1), .A(w3112) );
	vdp_nand g3665 (.Z(w3079), .A(w3625), .B(HCLK1) );
	vdp_nand g3666 (.Z(w3030), .A(w4048), .B(HCLK1) );
	vdp_nor g3667 (.Z(w4049), .A(w3415), .B(w3472) );
	vdp_nand g3668 (.Z(w3128), .A(w4128), .B(HCLK1) );
	vdp_nand g3669 (.Z(w3369), .A(M5), .B(w3373) );
	vdp_nand g3670 (.Z(w3368), .A(M5), .B(w4025) );
	vdp_xor g3671 (.Z(w3545), .A(w3544), .B(w3543) );
	vdp_aon22 g3672 (.Z(w3543), .A1(w3541), .B1(w3620), .A2(VPOS[3]), .B2(w3542) );
	vdp_xnor g3673 (.Z(w3547), .A(w3544), .B(w3621) );
	vdp_aon22 g3674 (.Z(w3621), .A1(w3541), .B1(w3620), .A2(VPOS[2]), .B2(w3546) );
	vdp_xnor g3675 (.Z(w3549), .A(w3544), .B(w3619) );
	vdp_aon22 g3676 (.Z(w3619), .A1(w3541), .B1(w3620), .A2(VPOS[1]), .B2(w3548) );
	vdp_notif0 g3677 (.nZ(VRAMA[4]), .A(w3547), .nE(w3598) );
	vdp_notif0 g3678 (.nZ(VRAMA[3]), .A(w3549), .nE(w3598) );
	vdp_xnor g3679 (.Z(w3617), .A(w3544), .B(w3618) );
	vdp_aon22 g3680 (.Z(w3618), .A1(w3541), .B1(w3620), .A2(VPOS[0]), .B2(w3550) );
	vdp_notif0 g3681 (.nZ(VRAMA[2]), .A(w3617), .nE(w3598) );
	vdp_notif0 g3682 (.nZ(VRAMA[1]), .A(w3616), .nE(w3598) );
	vdp_notif0 g3683 (.nZ(VRAMA[0]), .A(1'b1), .nE(w3598) );
	vdp_not g3684 (.nZ(w3613), .A(w3624) );
	vdp_not g3685 (.nZ(w3598), .A(w3623) );
	vdp_comp_we g3686 (.Z(w3541), .nZ(w3620), .A(w4122) );
	vdp_comp_we g3687 (.Z(w3551), .nZ(w3615), .A(w1) );
	vdp_notif0 g3688 (.nZ(VRAMA[5]), .A(w3553), .nE(w3613) );
	vdp_aoi22 g3689 (.Z(w3553), .A1(w3545), .B1(w3552), .A2(w3551), .B2(w3615) );
	vdp_notif0 g3690 (.nZ(VRAMA[6]), .A(w3554), .nE(w3613) );
	vdp_aoi22 g3691 (.Z(w3554), .A1(w3552), .B1(w3555), .A2(w3551), .B2(w3615) );
	vdp_notif0 g3692 (.nZ(VRAMA[7]), .A(w3556), .nE(w3613) );
	vdp_aoi22 g3693 (.Z(w3556), .A1(w3555), .B1(w3557), .A2(w3551), .B2(w3615) );
	vdp_notif0 g3694 (.nZ(VRAMA[8]), .A(w3558), .nE(w3613) );
	vdp_aoi22 g3695 (.Z(w3558), .A1(w3557), .B1(w3559), .A2(w3551), .B2(w3615) );
	vdp_notif0 g3696 (.nZ(VRAMA[9]), .A(w4057), .nE(w3613) );
	vdp_aoi22 g3697 (.Z(w4057), .A1(w3559), .B1(w3561), .A2(w3551), .B2(w3615) );
	vdp_notif0 g3698 (.nZ(VRAMA[10]), .A(w3560), .nE(w3613) );
	vdp_aoi22 g3699 (.Z(w3560), .A1(w3561), .B1(w3562), .A2(w3551), .B2(w3615) );
	vdp_notif0 g3700 (.nZ(VRAMA[11]), .A(w4056), .nE(w3613) );
	vdp_aoi22 g3701 (.Z(w4056), .A1(w3562), .B1(w3564), .A2(w3551), .B2(w3615) );
	vdp_notif0 g3702 (.nZ(VRAMA[12]), .A(w3565), .nE(w3613) );
	vdp_aoi22 g3703 (.Z(w3565), .A1(w3564), .B1(w3563), .A2(w3551), .B2(w3615) );
	vdp_notif0 g3704 (.nZ(VRAMA[13]), .A(w3567), .nE(w3613) );
	vdp_aoi22 g3705 (.Z(w3567), .A1(w3563), .B1(w3566), .A2(w3551), .B2(w3615) );
	vdp_not g3706 (.nZ(w3614), .A(w4077) );
	vdp_notif0 g3707 (.nZ(VRAMA[14]), .A(w3569), .nE(w3614) );
	vdp_aoi22 g3708 (.Z(w3569), .A1(w3566), .B1(w3568), .A2(w3551), .B2(w3615) );
	vdp_notif0 g3709 (.nZ(VRAMA[15]), .A(w3571), .nE(w3614) );
	vdp_aoi22 g3710 (.Z(w3571), .A1(w3568), .B1(w3570), .A2(w3551), .B2(w3615) );
	vdp_notif0 g3711 (.nZ(VRAMA[16]), .A(w3573), .nE(w3614) );
	vdp_aoi22 g3712 (.Z(w3573), .A1(w3570), .B1(w3572), .A2(w3551), .B2(w3615) );
	vdp_notif0 g3713 (.nZ(VRAMA[5]), .A(w3576), .nE(w3612) );
	vdp_aoi22 g3714 (.Z(w3576), .A1(w3574), .B1(w3545), .A2(w3575), .B2(w3611) );
	vdp_notif0 g3715 (.nZ(VRAMA[6]), .A(w3578), .nE(w3612) );
	vdp_aoi22 g3716 (.Z(w3578), .A1(w3574), .B1(w3575), .A2(w3577), .B2(w3611) );
	vdp_notif0 g3717 (.nZ(VRAMA[7]), .A(w3579), .nE(w3612) );
	vdp_aoi22 g3718 (.Z(w3579), .A1(w3574), .B1(w3577), .A2(w3597), .B2(w3611) );
	vdp_notif0 g3719 (.nZ(VRAMA[8]), .A(w3580), .nE(w3612) );
	vdp_aoi22 g3720 (.Z(w3580), .A1(w3574), .B1(w3597), .A2(w3581), .B2(w3611) );
	vdp_notif0 g3721 (.nZ(VRAMA[9]), .A(w3582), .nE(w3612) );
	vdp_aoi22 g3722 (.Z(w3582), .A1(w3574), .B1(w3581), .A2(w3583), .B2(w3611) );
	vdp_notif0 g3723 (.nZ(VRAMA[10]), .A(w3585), .nE(w3612) );
	vdp_aoi22 g3724 (.Z(w3585), .A1(w3574), .B1(w3583), .A2(w3584), .B2(w3611) );
	vdp_notif0 g3725 (.nZ(VRAMA[11]), .A(w3587), .nE(w3610) );
	vdp_aoi22 g3726 (.Z(w3587), .A1(w3574), .B1(w3584), .A2(w3586), .B2(w3611) );
	vdp_notif0 g3727 (.nZ(VRAMA[12]), .A(w3589), .nE(w3610) );
	vdp_aoi22 g3728 (.Z(w3589), .A1(w3574), .B1(w3586), .A2(w3588), .B2(w3611) );
	vdp_notif0 g3729 (.nZ(VRAMA[14]), .A(w3592), .nE(w3610) );
	vdp_aoi22 g3730 (.Z(w3592), .A1(w3574), .B1(w3590), .A2(w3593), .B2(w3611) );
	vdp_notif0 g3731 (.nZ(VRAMA[15]), .A(w3595), .nE(w3610) );
	vdp_aoi22 g3732 (.Z(w3595), .A1(w3574), .B1(w3593), .A2(w3594), .B2(w3611) );
	vdp_notif0 g3733 (.nZ(VRAMA[16]), .A(w3596), .nE(w3610) );
	vdp_aoi22 g3734 (.Z(w3596), .A1(w3574), .B1(w3594), .A2(w3572), .B2(w3611) );
	vdp_notif0 g3735 (.nZ(VRAMA[13]), .A(w3591), .nE(w3610) );
	vdp_aoi22 g3736 (.Z(w3591), .A1(w3574), .B1(w3588), .A2(w3590), .B2(w3611) );
	vdp_not g3737 (.nZ(w3612), .A(w3540) );
	vdp_comp_we g3738 (.Z(w3611), .nZ(w3574), .A(w1) );
	vdp_aon22 g3739 (.Z(w3572), .A1(w3535), .B1(w3534), .A2(w3536), .B2(w3607) );
	vdp_not g3740 (.nZ(w3610), .A(w3540) );
	vdp_not g3741 (.nZ(w3536), .A(w3607) );
	vdp_sr_bit g3742 (.Q(w3623), .D(w3638), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3743 (.Q(w3607), .D(HPOS[3]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3744 (.Q(w3616), .D(w3677), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3745 (.Q(w3624), .D(w4130), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3746 (.Q(w3622), .D(w4121), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3747 (.Q(w3642), .D(w4120), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3748 (.Q(w3609), .D(w4119), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3749 (.Q(w4095), .D(w4096), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3750 (.Q(w4097), .D(w4095), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3751 (.Q(w3625), .D(w4097), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3752 (.Q(w3657), .D(w109), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3753 (.Q(w3635), .D(w37), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3754 (.Q(w4098), .D(w38), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3755 (.Q(w3699), .D(w4098), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3756 (.Q(w3700), .D(w3635), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3757 (.Q(w3697), .D(w3657), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3758 (.Q(w3701), .D(w3608), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3759 (.Q(w3702), .D(w3172), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3760 (.Q(w3703), .D(w3173), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3761 (.Q(w3704), .D(w3171), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3762 (.Q(w3732), .D(w3170), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3763 (.Q(w3733), .D(w3169), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g3764 (.Q(w3633), .D(w3631), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3765 (.Q(w3634), .D(w3633), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_sr_bit g3766 (.Q(w4099), .D(w3634), .C1(DCLK2), .C2(DCLK1), .nC2(nDCLK1), .nC1(nDCLK2) );
	vdp_aon22 g3767 (.Z(w3647), .A1(H40), .B1(HPOS[8]), .A2(w3645), .B2(w3644) );
	vdp_aon22 g3768 (.Z(w3729), .A1(w3627), .B1(HPOS[8]), .A2(w3647), .B2(w3637) );
	vdp_aon22 g3769 (.Z(w3692), .A1(w3632), .B1(w3645), .A2(w3647), .B2(w3637) );
	vdp_or3 g3770 (.Z(w3698), .A(w3657), .B(w3635), .C(w4098) );
	vdp_or g3771 (.Z(w3648), .A(M5), .B(w3462) );
	vdp_bufif0 g3772 (.Z(VRAMA[1]), .A(w4094), .nE(w3636) );
	vdp_or g3773 (.Z(w3725), .A(w3647), .B(HPOS[4]) );
	vdp_bufif0 g3774 (.Z(VRAMA[2]), .A(w3650), .nE(w3636) );
	vdp_or g3775 (.Z(w3726), .A(w3647), .B(HPOS[5]) );
	vdp_bufif0 g3776 (.Z(VRAMA[3]), .A(w3651), .nE(w3636) );
	vdp_or g3777 (.Z(w3730), .A(w3647), .B(HPOS[6]) );
	vdp_bufif0 g3778 (.Z(VRAMA[4]), .A(w3652), .nE(w3636) );
	vdp_or g3779 (.Z(w3728), .A(w3647), .B(HPOS[7]) );
	vdp_bufif0 g3780 (.Z(VRAMA[5]), .A(w3653), .nE(w3636) );
	vdp_bufif0 g3781 (.Z(VRAMA[5]), .A(w3626), .nE(w3636) );
	vdp_not g3782 (.nZ(w3641), .A(w3533) );
	vdp_not g3783 (.nZ(w4100), .A(HPOS[3]) );
	vdp_dlatch_inv g3784 (.nQ(w3631), .D(w3630), .C(DCLK1), .nC(nDCLK1) );
	vdp_not g3785 (.nZ(w3645), .A(w4076) );
	vdp_not g3786 (.nZ(w3637), .A(w3647) );
	vdp_not g3787 (.nZ(w3644), .A(H40) );
	vdp_not g3788 (.nZ(w3636), .A(w3643) );
	vdp_bufif0 g3789 (.Z(VRAMA[0]), .A(1'b0), .nE(w3636) );
	vdp_or g3790 (.Z(w3643), .A(w3622), .B(w3642) );
	vdp_or g3791 (.Z(w4096), .A(w3640), .B(w6) );
	vdp_nand3 g3792 (.Z(w3696), .A(M5), .B(w3641), .C(HPOS[3]) );
	vdp_nand3 g3793 (.Z(w3655), .A(M5), .B(w3641), .C(w4100) );
	vdp_and g3794 (.Z(w3656), .A(DCLK2), .B(w4099) );
	vdp_and g3795 (.Z(w3629), .A(w3634), .B(DCLK2) );
	vdp_and g3796 (.Z(w3695), .A(w3633), .B(DCLK2) );
	vdp_and g3797 (.Z(w3628), .A(w3631), .B(DCLK2) );
	vdp_and g3798 (.Z(w4077), .A(M5), .B(w3624) );
	vdp_and g3799 (.Z(w3685), .A(HPOS[3]), .B(w3646) );
	vdp_and g3800 (.Z(w4119), .A(w3533), .B(w6) );
	vdp_and g3801 (.Z(w4120), .A(w3641), .B(w6) );
	vdp_and3 g3802 (.Z(w4121), .A(w3640), .B(M5), .C(w3639) );
	vdp_nor g3803 (.Z(w3646), .A(M5), .B(w3647) );
	vdp_nand g3804 (.Z(w3630), .A(w3283), .B(HCLK1) );
	vdp_oai21 g3805 (.A1(HPOS[6]), .A2(HPOS[7]), .B(HPOS[8]), .Z(w4076) );
	vdp_slatch g3806 (.Q(w3672), .D(REG_BUS[0]), .C(w3720), .nC(w3719) );
	vdp_slatch g3807 (.Q(w3668), .D(S[0]), .C(w3715), .nC(w3714) );
	vdp_slatch g3808 (.Q(w3669), .D(S[0]), .C(w3716), .nC(w3713) );
	vdp_slatch g3809 (.Q(w3670), .D(REG_BUS[1]), .C(w3720), .nC(w3719) );
	vdp_slatch g3810 (.Q(w3666), .D(S[1]), .C(w3715), .nC(w3714) );
	vdp_slatch g3811 (.Q(w3741), .D(S[1]), .C(w3716), .nC(w3713) );
	vdp_slatch g3812 (.Q(w3742), .D(REG_BUS[2]), .C(w3720), .nC(w3719) );
	vdp_slatch g3813 (.Q(w3660), .D(S[2]), .C(w3715), .nC(w3714) );
	vdp_slatch g3814 (.Q(w3743), .D(S[2]), .C(w3716), .nC(w3713) );
	vdp_slatch g3815 (.Q(w3739), .D(REG_BUS[3]), .C(w3720), .nC(w3719) );
	vdp_slatch g3816 (.Q(w3738), .D(S[3]), .C(w3715), .nC(w3714) );
	vdp_slatch g3817 (.Q(w4418), .D(S[3]), .C(w3716), .nC(w3713) );
	vdp_slatch g3818 (.Q(w3684), .D(REG_BUS[4]), .C(w3720), .nC(w3719) );
	vdp_slatch g3819 (.Q(w3737), .D(S[4]), .C(w3715), .nC(w3714) );
	vdp_slatch g3820 (.Q(w3736), .D(S[4]), .C(w3716), .nC(w3713) );
	vdp_slatch g3821 (.Q(w3735), .D(REG_BUS[5]), .C(w3720), .nC(w3719) );
	vdp_slatch g3822 (.Q(w3723), .D(S[5]), .C(w3715), .nC(w3714) );
	vdp_slatch g3823 (.Q(w3722), .D(S[5]), .C(w3716), .nC(w3713) );
	vdp_slatch g3824 (.Q(w3721), .D(REG_BUS[6]), .C(w3720), .nC(w3719) );
	vdp_slatch g3825 (.Q(w3717), .D(S[6]), .C(w3715), .nC(w3714) );
	vdp_slatch g3826 (.Q(w3718), .D(S[6]), .C(w3716), .nC(w3713) );
	vdp_slatch g3827 (.Q(w3712), .D(REG_BUS[7]), .C(w3720), .nC(w3719) );
	vdp_slatch g3828 (.Q(w3711), .D(S[7]), .C(w3715), .nC(w3714) );
	vdp_slatch g3829 (.Q(w3710), .D(S[7]), .C(w3716), .nC(w3713) );
	vdp_slatch g3830 (.Q(w3708), .D(S[0]), .C(w3688), .nC(w3705) );
	vdp_slatch g3831 (.Q(w3690), .D(S[0]), .C(w3689), .nC(w3709) );
	vdp_slatch g3832 (.Q(w3694), .D(S[1]), .C(w3689), .nC(w3709) );
	vdp_slatch g3833 (.Q(w3693), .D(S[1]), .C(w3688), .nC(w3705) );
	vdp_slatch g3834 (.Q(w3686), .D(w3712), .C(w3665), .nC(w3664) );
	vdp_slatch g3835 (.Q(w3680), .D(w3721), .C(w3665), .nC(w3664) );
	vdp_slatch g3836 (.Q(w3683), .D(w3735), .C(w3665), .nC(w3664) );
	vdp_slatch g3837 (.Q(w3745), .D(w3684), .C(w3665), .nC(w3664) );
	vdp_slatch g3838 (.Q(w3658), .D(w3739), .C(w3665), .nC(w3664) );
	vdp_slatch g3839 (.Q(w3659), .D(w3742), .C(w3665), .nC(w3664) );
	vdp_slatch g3840 (.Q(w3667), .D(w3670), .C(w3665), .nC(w3664) );
	vdp_slatch g3841 (.Q(w3671), .D(w3672), .C(w3665), .nC(w3664) );
	vdp_fa g3842 (.CI(w4074), .SUM(w4019), .B(w3692), .A(w3707) );
	vdp_fa g3843 (.CO(w4074), .CI(w3691), .SUM(w3891), .B(w3729), .A(w3734) );
	vdp_fa g3844 (.CO(w3734), .CI(w3687), .SUM(w3653), .B(w3728), .A(w4073) );
	vdp_fa g3845 (.CO(w4073), .CI(w3681), .SUM(w3652), .B(w3730), .A(w3731) );
	vdp_fa g3846 (.CO(w3731), .CI(w3682), .SUM(w3651), .B(w3726), .A(w3727) );
	vdp_fa g3847 (.CO(w3727), .CI(w3787), .SUM(w3650), .B(w3725), .A(w3724) );
	vdp_fa g3848 (.CO(w3724), .CI(w3648), .SUM(w4094), .B(w3685), .A(1'b1) );
	vdp_aon222 g3849 (.A1(w3662), .B1(w3649), .C1(w3661), .A2(w3693), .B2(w3694), .C2(1'b0), .Z(w3707) );
	vdp_aon222 g3850 (.A1(w3662), .B1(w3649), .C1(w3661), .A2(w3708), .B2(w3690), .C2(1'b0), .Z(w3691) );
	vdp_aon222 g3851 (.A1(w3662), .B1(w3649), .C1(w3661), .A2(w3710), .B2(w3711), .C2(w3686), .Z(w3687) );
	vdp_aon222 g3852 (.A1(w3662), .B1(w3649), .C1(w3661), .A2(w3718), .B2(w3717), .C2(w3680), .Z(w3681) );
	vdp_aon222 g3853 (.A1(w3662), .B1(w3649), .C1(w3661), .A2(w3722), .B2(w3723), .C2(w3683), .Z(w3682) );
	vdp_aon222 g3854 (.A1(w3662), .B1(w3649), .C1(w3661), .A2(w3736), .B2(w3737), .C2(w3745), .Z(w3787) );
	vdp_aon222 g3855 (.A1(w3662), .B1(w3649), .C1(w3661), .A2(w4418), .B2(w3738), .C2(w3658), .Z(w3462) );
	vdp_aon222 g3856 (.A1(w3662), .B1(w3649), .C1(w3661), .A2(w3743), .B2(w3660), .C2(w3659), .Z(w3158) );
	vdp_aon222 g3857 (.A1(w3662), .B1(w3649), .A2(w3741), .B2(w3666), .C2(w3667), .Z(w3460), .C1(w3661) );
	vdp_aon222 g3858 (.A1(w3662), .B1(w3649), .C1(w3661), .A2(w3669), .B2(w3668), .C2(w3671), .Z(w3458) );
	vdp_comp_strong g3859 (.Z(w3688), .nZ(w3705), .A(w3656) );
	vdp_comp_strong g3860 (.Z(w3689), .nZ(w3709), .A(w3695) );
	vdp_not g3861 (.nZ(w3649), .A(w3655) );
	vdp_not g3862 (.nZ(w3662), .A(w3696) );
	vdp_not g3863 (.nZ(w3661), .A(w3740) );
	vdp_not g3864 (.nZ(w3675), .A(w96) );
	vdp_not g3865 (.nZ(w3639), .A(w104) );
	vdp_not g3866 (.nZ(w3676), .A(w3677) );
	vdp_not g3867 (.nZ(w3640), .A(w3678) );
	vdp_not g3868 (.nZ(w3679), .A(M5) );
	vdp_comp_strong g3869 (.Z(w3715), .nZ(w3714), .A(w3628) );
	vdp_comp_strong g3870 (.Z(w3716), .nZ(w3713), .A(w3629) );
	vdp_comp_strong g3871 (.Z(w3720), .nZ(w3719), .A(w86) );
	vdp_comp_strong g3872 (.Z(w3665), .nZ(w3664), .A(w3744) );
	vdp_or g3873 (.Z(w3740), .A(w4078), .B(M5) );
	vdp_or g3874 (.Z(w4130), .A(w13), .B(w3676) );
	vdp_or g3875 (.Z(w3638), .A(w13), .B(w14) );
	vdp_or g3876 (.Z(w3744), .A(w4), .B(w103) );
	vdp_or5 g3877 (.E(w3675), .C(w3674), .D(VPOS[5]), .Z(w4078), .A(w3673), .B(VPOS[4]) );
	vdp_aoi21 g3878 (.Z(w3678), .A1(w104), .A2(w3110), .B(w8) );
	vdp_nand g3879 (.Z(w3677), .A(w14), .B(w3679) );
	vdp_slatch g3880 (.Q(w3781), .D(w4408), .C(w3750), .nC(w3751) );
	vdp_slatch g3881 (.Q(w3756), .D(w4409), .C(w3750), .nC(w3751) );
	vdp_slatch g3882 (.Q(w3757), .D(w4410), .C(w3750), .nC(w3751) );
	vdp_slatch g3883 (.Q(w3758), .D(w4407), .C(w3750), .nC(w3751) );
	vdp_slatch g3884 (.Q(w3760), .D(w4406), .C(w3750), .nC(w3751) );
	vdp_slatch g3885 (.Q(w3759), .D(w4405), .C(w3750), .nC(w3751) );
	vdp_slatch g3886 (.nQ(w3765), .D(w4413), .C(w3752), .nC(w3753) );
	vdp_slatch g3887 (.Q(w3776), .D(w4414), .C(w3752), .nC(w3753) );
	vdp_slatch g3888 (.Q(w3764), .D(w4415), .C(w3752), .nC(w3753) );
	vdp_slatch g3889 (.Q(w3763), .D(w4416), .C(w3752), .nC(w3753) );
	vdp_slatch g3890 (.Q(w3762), .D(w4412), .C(w3752), .nC(w3753) );
	vdp_slatch g3891 (.Q(w3761), .D(w4411), .C(w3752), .nC(w3753) );
	vdp_comp_strong g3892 (.Z(w3750), .nZ(w3751), .A(w3770) );
	vdp_comp_strong g3893 (.Z(w3752), .nZ(w3753), .A(w4101) );
	vdp_cgi2a g3894 (.Z(w4018), .A(w3761), .B(HPOS[4]), .C(1'b1) );
	vdp_cgi2a g3895 (.Z(w4013), .A(w3762), .B(HPOS[5]), .C(w4018) );
	vdp_cgi2a g3896 (.Z(w4012), .A(w3763), .B(HPOS[6]), .C(w4013) );
	vdp_cgi2a g3897 (.Z(w4014), .A(w3764), .B(HPOS[7]), .C(w4012) );
	vdp_cgi2a g3898 (.X(w3766), .A(w3776), .B(HPOS[8]), .C(w4014) );
	vdp_cgi2a g3899 (.Z(w3771), .A(w3768), .B(w3756), .C(w4103) );
	vdp_cgi2a g3900 (.Z(w4103), .A(w3769), .B(w3757), .C(w4015) );
	vdp_cgi2a g3901 (.Z(w4015), .A(w3772), .B(w3758), .C(w4016) );
	vdp_cgi2a g3902 (.Z(w4016), .A(w3775), .B(w3760), .C(w4017) );
	vdp_cgi2a g3903 (.Z(w4017), .A(w3774), .B(w3759), .C(1'b0) );
	vdp_slatch g3904 (.Q(w4408), .D(REG_BUS[7]), .C(w3778), .nC(w3755) );
	vdp_slatch g3905 (.Q(w4409), .D(REG_BUS[4]), .C(w3778), .nC(w3755) );
	vdp_slatch g3906 (.Q(w4410), .D(REG_BUS[3]), .C(w3778), .nC(w3755) );
	vdp_slatch g3907 (.Q(w4407), .D(REG_BUS[2]), .C(w3778), .nC(w3755) );
	vdp_slatch g3908 (.Q(w4406), .D(REG_BUS[1]), .C(w3778), .nC(w3755) );
	vdp_slatch g3909 (.Q(w4405), .D(REG_BUS[0]), .C(w3778), .nC(w3755) );
	vdp_comp_strong g3910 (.Z(w3778), .nZ(w3755), .A(w75) );
	vdp_slatch g3911 (.Q(w4413), .D(REG_BUS[7]), .C(w3779), .nC(w3777) );
	vdp_slatch g3912 (.Q(w4414), .D(REG_BUS[4]), .C(w3779), .nC(w3777) );
	vdp_slatch g3913 (.Q(w4415), .D(REG_BUS[3]), .C(w3779), .nC(w3777) );
	vdp_slatch g3914 (.Q(w4416), .D(REG_BUS[2]), .C(w3779), .nC(w3777) );
	vdp_slatch g3915 (.Q(w4412), .D(REG_BUS[1]), .C(w3779), .nC(w3777) );
	vdp_slatch g3916 (.Q(w4411), .D(REG_BUS[0]), .C(w3779), .nC(w3777) );
	vdp_comp_strong g3917 (.Z(w3779), .nZ(w3777), .A(w74) );
	vdp_xor g3918 (.Z(w3780), .A(w3781), .B(w3771) );
	vdp_xor g3919 (.Z(w3767), .A(w3765), .B(w3766) );
	vdp_aon22 g3920 (.Z(w3768), .A1(w3773), .B1(w3784), .A2(VPOS[8]), .B2(VPOS[7]) );
	vdp_aon22 g3921 (.Z(w3769), .A1(w3773), .B1(w3784), .A2(VPOS[7]), .B2(VPOS[6]) );
	vdp_aon22 g3922 (.Z(w3772), .A1(w3773), .B1(w3784), .A2(VPOS[6]), .B2(VPOS[5]) );
	vdp_aon22 g3923 (.Z(w3775), .A1(w3773), .B1(w3784), .A2(VPOS[5]), .B2(VPOS[4]) );
	vdp_aon22 g3924 (.Z(w3774), .A1(w3773), .B1(w3784), .A2(VPOS[4]), .B2(VPOS[3]) );
	vdp_aon22 g3925 (.Z(w3792), .A1(w3773), .B1(w3784), .A2(VPOS[3]), .B2(VPOS[2]) );
	vdp_aon22 g3926 (.Z(w3791), .A1(w3773), .B1(w3784), .A2(VPOS[2]), .B2(VPOS[1]) );
	vdp_aon22 g3927 (.Z(w3790), .A1(w3773), .B1(w3784), .A2(VPOS[1]), .B2(VPOS[0]) );
	vdp_comp_we g3928 (.Z(w3773), .nZ(w3784), .A(w1) );
	vdp_not g3929 (.nZ(w3533), .A(w4102) );
	vdp_not g3930 (.nZ(w3783), .A(HPOS[3]) );
	vdp_not g3931 (.nZ(w4105), .A(w4104) );
	vdp_or g3932 (.Z(w4101), .A(w103), .B(w4) );
	vdp_or g3933 (.Z(w3770), .A(w103), .B(w4105) );
	vdp_oai21 g3934 (.Z(w4104), .A1(w5), .A2(M5), .B(w4) );
	vdp_and g3935 (.Z(w3782), .A(w3767), .B(w3785) );
	vdp_oai211 g3936 (.Z(w4102), .A1(w3783), .A2(M5), .B(w3782), .C(w3780) );
	vdp_slatch g3937 (.nQ(w3825), .D(REG_BUS[4]), .C(w3797), .nC(w3798) );
	vdp_slatch g3938 (.nQ(w3827), .D(REG_BUS[4]), .C(w3795), .nC(w3796) );
	vdp_slatch g3939 (.nQ(w3826), .D(REG_BUS[5]), .C(w3797), .nC(w3798) );
	vdp_slatch g3940 (.nQ(w3828), .D(REG_BUS[5]), .C(w3795), .nC(w3796) );
	vdp_slatch g3941 (.nQ(w3801), .D(REG_BUS[6]), .C(w3797), .nC(w3798) );
	vdp_slatch g3942 (.nQ(w3802), .D(REG_BUS[6]), .C(w3795), .nC(w3796) );
	vdp_slatch g3943 (.nQ(w4404), .D(REG_BUS[1]), .C(w3795), .nC(w3796) );
	vdp_slatch g3944 (.nQ(w3821), .D(REG_BUS[2]), .C(w3797), .nC(w3798) );
	vdp_slatch g3945 (.nQ(w3822), .D(REG_BUS[2]), .C(w3795), .nC(w3796) );
	vdp_slatch g3946 (.nQ(w3823), .D(REG_BUS[3]), .C(w3797), .nC(w3798) );
	vdp_slatch g3947 (.nQ(w3824), .D(REG_BUS[3]), .C(w3795), .nC(w3796) );
	vdp_slatch g3948 (.nQ(w3829), .D(REG_BUS[0]), .C(w3795), .nC(w3796) );
	vdp_slatch g3949 (.nQ(w3799), .D(REG_BUS[1]), .C(w3797), .nC(w3798) );
	vdp_slatch g3950 (.Q(w3535), .D(REG_BUS[0]), .C(w3788), .nC(w3789) );
	vdp_slatch g3951 (.Q(w3534), .D(REG_BUS[4]), .C(w3788), .nC(w3789) );
	vdp_not g3952 (.nZ(w4107), .A(w3799) );
	vdp_aoi22 g3953 (.Z(w3818), .A1(HPOS[8]), .B1(w3774), .A2(w3794), .B2(w3793) );
	vdp_aoi22 g3954 (.Z(w3819), .A1(w3774), .B1(w3775), .A2(w3794), .B2(w3793) );
	vdp_aoi22 g3955 (.Z(w3806), .A1(w3775), .B1(w3772), .A2(w3794), .B2(w3793) );
	vdp_aoi22 g3956 (.Z(w3831), .A1(w3769), .B1(w3768), .A2(w3794), .B2(w3793) );
	vdp_aoi22 g3957 (.Z(w3820), .A1(w3772), .B1(w3769), .A2(w3794), .B2(w3793) );
	vdp_comp_strong g3958 (.Z(w3788), .nZ(w3789), .A(w85) );
	vdp_comp_strong g3959 (.Z(w3797), .nZ(w3798), .A(w71) );
	vdp_comp_strong g3960 (.Z(w3795), .nZ(w3796), .A(w68) );
	vdp_aoi22 g3961 (.Z(w3830), .A1(w3768), .B1(w3793), .A2(w3794), .B2(w4107) );
	vdp_nand g3962 (.Z(w3832), .A(w3768), .B(w93) );
	vdp_nand g3963 (.Z(w3805), .A(w3769), .B(w93) );
	vdp_nand g3964 (.Z(w3833), .A(w3775), .B(w93) );
	vdp_nand g3965 (.Z(w3807), .A(w3772), .B(w93) );
	vdp_nand g3966 (.Z(w3817), .A(w3774), .B(w93) );
	vdp_nand g3967 (.Z(w4106), .A(w3792), .B(w91) );
	vdp_nand g3968 (.Z(w4131), .A(w3791), .B(w91) );
	vdp_nand g3969 (.Z(w3813), .A(w3790), .B(w91) );
	vdp_nand g3970 (.Z(w3785), .A(HPOS[7]), .B(HPOS[8]) );
	vdp_comp_we g3971 (.Z(w3794), .nZ(w3793), .A(H40) );
	vdp_notif0 g3972 (.nZ(VRAMA[16]), .A(w3802), .nE(w3800) );
	vdp_notif0 g3973 (.nZ(VRAMA[16]), .A(w3801), .nE(w3804) );
	vdp_notif0 g3974 (.nZ(VRAMA[15]), .A(w3828), .nE(w3800) );
	vdp_notif0 g3975 (.nZ(VRAMA[15]), .A(w3826), .nE(w3804) );
	vdp_notif0 g3976 (.nZ(VRAMA[14]), .A(w3827), .nE(w3800) );
	vdp_notif0 g3977 (.nZ(VRAMA[14]), .A(w3825), .nE(w3804) );
	vdp_notif0 g3978 (.nZ(VRAMA[13]), .A(w3824), .nE(w3800) );
	vdp_notif0 g3979 (.nZ(VRAMA[13]), .A(w3823), .nE(w3804) );
	vdp_notif0 g3980 (.nZ(VRAMA[12]), .A(w3822), .nE(w3800) );
	vdp_notif0 g3981 (.nZ(VRAMA[12]), .A(w3821), .nE(w3804) );
	vdp_notif0 g3982 (.nZ(VRAMA[11]), .A(w4404), .nE(w3800) );
	vdp_notif0 g3983 (.nZ(VRAMA[11]), .A(w3830), .nE(w3804) );
	vdp_notif0 g3984 (.nZ(VRAMA[10]), .A(w3829), .nE(w3800) );
	vdp_notif0 g3985 (.nZ(VRAMA[10]), .A(w3831), .nE(w3804) );
	vdp_notif0 g3986 (.nZ(VRAMA[9]), .A(w3832), .nE(w3803) );
	vdp_notif0 g3987 (.nZ(VRAMA[9]), .A(w3820), .nE(w3804) );
	vdp_notif0 g3988 (.nZ(VRAMA[6]), .A(w3833), .nE(w3803) );
	vdp_notif0 g3989 (.nZ(VRAMA[6]), .A(w3818), .nE(w3808) );
	vdp_notif0 g3990 (.nZ(VRAMA[5]), .A(w3817), .nE(w3803) );
	vdp_notif0 g3991 (.nZ(VRAMA[5]), .A(w3816), .nE(w3808) );
	vdp_notif0 g3992 (.nZ(VRAMA[4]), .A(w4106), .nE(w3803) );
	vdp_notif0 g3993 (.nZ(VRAMA[4]), .A(w3815), .nE(w3808) );
	vdp_notif0 g3994 (.nZ(VRAMA[3]), .A(w4131), .nE(w3803) );
	vdp_notif0 g3995 (.nZ(VRAMA[3]), .A(w3814), .nE(w3808) );
	vdp_notif0 g3996 (.nZ(VRAMA[2]), .A(w3813), .nE(w3803) );
	vdp_notif0 g3997 (.nZ(VRAMA[2]), .A(w3812), .nE(w3808) );
	vdp_notif0 g3998 (.nZ(VRAMA[1]), .A(1'b1), .nE(w3803) );
	vdp_notif0 g3999 (.nZ(VRAMA[1]), .A(1'b1), .nE(w3808) );
	vdp_notif0 g4000 (.nZ(VRAMA[0]), .A(w3810), .nE(w3803) );
	vdp_notif0 g4001 (.nZ(VRAMA[0]), .A(w3810), .nE(w3808) );
	vdp_notif0 g4002 (.nZ(VRAMA[8]), .A(w3805), .nE(w3803) );
	vdp_notif0 g4003 (.nZ(VRAMA[8]), .A(w3806), .nE(w3808) );
	vdp_notif0 g4004 (.nZ(VRAMA[7]), .A(w3807), .nE(w3803) );
	vdp_notif0 g4005 (.nZ(VRAMA[7]), .A(w3819), .nE(w3808) );
	vdp_not g4006 (.nZ(w3810), .A(1'b0) );
	vdp_not g4007 (.nZ(w3812), .A(HPOS[4]) );
	vdp_not g4008 (.nZ(w3814), .A(HPOS[5]) );
	vdp_not g4009 (.nZ(w3815), .A(HPOS[6]) );
	vdp_not g4010 (.nZ(w3816), .A(HPOS[7]) );
	vdp_not g4011 (.nZ(w3803), .A(w3282) );
	vdp_not g4012 (.nZ(w3800), .A(w3282) );
	vdp_not g4013 (.nZ(w3808), .A(w3609) );
	vdp_not g4014 (.nZ(w3804), .A(w3609) );
	vdp_not g4015 (.nZ(w3842), .A(w4011) );
	vdp_comp_strong g4016 (.Z(w3836), .nZ(w3837), .A(w70) );
	vdp_comp_we g4017 (.Z(w3841), .nZ(w3840), .A(w3622) );
	vdp_comp_strong g4018 (.Z(w3839), .nZ(w3838), .A(w72) );
	vdp_slatch g4019 (.Q(w3862), .D(REG_BUS[6]), .C(w3836), .nC(w3837) );
	vdp_slatch g4020 (.Q(w4116), .D(REG_BUS[3]), .C(w3839), .nC(w3838) );
	vdp_slatch g4021 (.Q(w3861), .D(REG_BUS[5]), .C(w3836), .nC(w3837) );
	vdp_slatch g4022 (.Q(w3859), .D(REG_BUS[2]), .C(w3839), .nC(w3838) );
	vdp_slatch g4023 (.Q(w3845), .D(REG_BUS[4]), .C(w3836), .nC(w3837) );
	vdp_slatch g4024 (.Q(w4419), .D(REG_BUS[1]), .C(w3839), .nC(w3838) );
	vdp_slatch g4025 (.Q(w3848), .D(REG_BUS[3]), .C(w3836), .nC(w3837) );
	vdp_slatch g4026 (.Q(w4117), .D(REG_BUS[0]), .C(w3839), .nC(w3838) );
	vdp_slatch g4027 (.Q(w3856), .D(REG_BUS[1]), .C(w3836), .nC(w3837) );
	vdp_slatch g4028 (.Q(w3853), .D(REG_BUS[2]), .C(w3836), .nC(w3837) );
	vdp_bufif0 g4029 (.Z(VRAMA[11]), .A(w3855), .nE(w3844) );
	vdp_bufif0 g4030 (.Z(VRAMA[10]), .A(w3849), .nE(w3844) );
	vdp_bufif0 g4031 (.Z(VRAMA[13]), .A(w3857), .nE(w3844) );
	vdp_bufif0 g4032 (.Z(VRAMA[9]), .A(w3847), .nE(w3844) );
	vdp_bufif0 g4033 (.Z(VRAMA[8]), .A(w3846), .nE(w3844) );
	vdp_bufif0 g4034 (.Z(VRAMA[14]), .A(w3858), .nE(w3842) );
	vdp_bufif0 g4035 (.Z(VRAMA[7]), .A(w3843), .nE(w3844) );
	vdp_bufif0 g4036 (.Z(VRAMA[15]), .A(w4075), .nE(w3842) );
	vdp_bufif0 g4037 (.Z(VRAMA[16]), .A(w3860), .nE(w3842) );
	vdp_aon22 g4038 (.Z(w3860), .A1(w3840), .B1(w3841), .A2(w3862), .B2(w4116) );
	vdp_aon22 g4039 (.Z(w4075), .A1(w3840), .B1(w3841), .A2(w3861), .B2(w3859) );
	vdp_aon22 g4040 (.Z(w3858), .A1(w3840), .B1(w3841), .A2(w3845), .B2(w4419) );
	vdp_aon22 g4041 (.Z(w3857), .A1(w3840), .B1(w3841), .A2(w3848), .B2(w4117) );
	vdp_aon22 g4042 (.Z(w3855), .A1(w3851), .B1(w3854), .A2(w3856), .B2(w3852) );
	vdp_aon22 g4043 (.Z(w3850), .A1(w3851), .B1(w3865), .A2(w3853), .B2(w3852) );
	vdp_bufif0 g4044 (.Z(VRAMA[12]), .A(w3850), .nE(w3844) );
	vdp_not g4045 (.nZ(w3844), .A(w3643) );
	vdp_and g4046 (.Z(w4011), .A(w3643), .B(M5) );
	vdp_comp_we g4047 (.Z(w3852), .nZ(w3851), .A(M5) );
	vdp_fa g4048 (.CO(w3880), .CI(w4064), .SUM(w3900), .B(VPOS[6]), .A(w4063) );
	vdp_fa g4049 (.CO(w4063), .CI(w4066), .SUM(w3881), .B(VPOS[5]), .A(w4065) );
	vdp_fa g4050 (.CO(w4065), .CI(w4068), .SUM(w3882), .B(VPOS[4]), .A(w4067) );
	vdp_fa g4051 (.CO(w4067), .CI(w3948), .SUM(w3542), .B(VPOS[3]), .A(w4069) );
	vdp_fa g4052 (.CO(w4069), .CI(w4071), .SUM(w3546), .B(VPOS[2]), .A(w4070) );
	vdp_fa g4053 (.CO(w4070), .CI(w4006), .SUM(w3548), .B(VPOS[1]), .A(w4072) );
	vdp_fa g4054 (.CO(w4072), .CI(w3961), .SUM(w3550), .B(VPOS[0]), .A(1'b0) );
	vdp_fa g4055 (.CO(w3899), .CI(w4062), .SUM(w3897), .B(VPOS[7]), .A(w3880) );
	vdp_fa g4056 (.CO(w3879), .CI(w3934), .SUM(w3908), .B(VPOS[8]), .A(w3899) );
	vdp_fa g4057 (.CO(w3907), .CI(w3935), .SUM(w3874), .B(1'b0), .A(w3879) );
	vdp_fa g4058 (.CI(w3919), .SUM(w3875), .B(1'b0), .A(w3907) );
	vdp_aon22 g4059 (.Z(w3919), .A1(w3917), .B1(w3918), .A2(w3878), .B2(w3877) );
	vdp_aon22 g4060 (.Z(w3935), .A1(w4009), .B1(w3922), .A2(w3878), .B2(w3877) );
	vdp_aon22 g4061 (.Z(w3934), .A1(w3923), .B1(w3924), .A2(w3878), .B2(w3877) );
	vdp_aon22 g4062 (.Z(w4062), .A1(w3926), .B1(w3927), .A2(w3878), .B2(w3877) );
	vdp_aon22 g4063 (.Z(w4064), .A1(w3933), .B1(w3930), .A2(w3878), .B2(w3877) );
	vdp_aon22 g4064 (.Z(w4066), .A1(w3938), .B1(w3937), .A2(w3878), .B2(w3877) );
	vdp_aon22 g4065 (.Z(w4068), .A1(w3942), .B1(w3943), .A2(w3878), .B2(w3877) );
	vdp_aon22 g4066 (.Z(w3948), .A1(w3947), .B1(w3946), .A2(w3878), .B2(w3877) );
	vdp_aon22 g4067 (.Z(w4071), .A1(w3949), .B1(w3950), .A2(w3878), .B2(w3877) );
	vdp_aon22 g4068 (.Z(w4006), .A1(w3953), .B1(w4010), .A2(w3878), .B2(w3877) );
	vdp_aon22 g4069 (.Z(w3961), .A1(w3955), .B1(w3954), .A2(w3878), .B2(w3877) );
	vdp_comp_we g4070 (.Z(w3878), .nZ(w3877), .A(w3886) );
	vdp_comp_strong g4071 (.Z(w3888), .nZ(w3883), .A(w69) );
	vdp_sr_bit g4072 (.Q(w3909), .D(RD_DATA[1]), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4073 (.Q(w3884), .D(RD_DATA[2]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4074 (.Q(w3958), .D(w3909), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4075 (.Q(w3976), .D(w3884), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4076 (.Q(w3957), .D(HPOS[3]), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4077 (.Q(w3627), .D(REG_BUS[0]), .C(w3888), .nC(w3883) );
	vdp_slatch g4078 (.Q(w3632), .D(REG_BUS[1]), .C(w3888), .nC(w3883) );
	vdp_slatch g4079 (.Q(w3904), .D(REG_BUS[5]), .C(w3888), .nC(w3883) );
	vdp_slatch g4080 (.Q(w3903), .D(REG_BUS[4]), .C(w3888), .nC(w3883) );
	vdp_slatch g4081 (.Q(w3955), .D(w3959), .C(w3910), .nC(w3914) );
	vdp_slatch g4082 (.Q(w4127), .D(w3960), .C(w3916), .nC(w3911) );
	vdp_slatch g4083 (.Q(w3953), .D(w3952), .C(w3910), .nC(w3914) );
	vdp_slatch g4084 (.Q(w4126), .D(w3951), .C(w3916), .nC(w3911) );
	vdp_slatch g4085 (.Q(w3949), .D(w3978), .C(w3910), .nC(w3914) );
	vdp_slatch g4086 (.Q(w4125), .D(w3945), .C(w3916), .nC(w3911) );
	vdp_slatch g4087 (.Q(w3947), .D(w3944), .C(w3910), .nC(w3914) );
	vdp_slatch g4088 (.Q(w4124), .D(w3941), .C(w3916), .nC(w3911) );
	vdp_slatch g4089 (.Q(w3942), .D(w3940), .C(w3910), .nC(w3914) );
	vdp_slatch g4090 (.Q(w4123), .D(w3939), .C(w3916), .nC(w3911) );
	vdp_slatch g4091 (.Q(w3938), .D(w3932), .C(w3910), .nC(w3914) );
	vdp_slatch g4092 (.Q(w4134), .D(w3931), .C(w3916), .nC(w3911) );
	vdp_slatch g4093 (.Q(w3933), .D(w3928), .C(w3910), .nC(w3914) );
	vdp_slatch g4094 (.Q(w4135), .D(w3929), .C(w3916), .nC(w3911) );
	vdp_slatch g4095 (.Q(w3926), .D(w3925), .C(w3910), .nC(w3914) );
	vdp_slatch g4096 (.Q(w3924), .D(w3936), .C(w3916), .nC(w3911) );
	vdp_slatch g4097 (.Q(w3923), .D(w3983), .C(w3910), .nC(w3914) );
	vdp_slatch g4098 (.Q(w3922), .D(w3921), .C(w3916), .nC(w3911) );
	vdp_slatch g4099 (.Q(w4009), .D(w3920), .C(w3910), .nC(w3914) );
	vdp_slatch g4100 (.Q(w3918), .D(w3998), .C(w3916), .nC(w3911) );
	vdp_slatch g4101 (.Q(w3917), .D(w3915), .C(w3910), .nC(w3914) );
	vdp_slatch g4102 (.Q(w4110), .D(REG_BUS[0]), .C(w3967), .nC(w3966) );
	vdp_aon22 g4103 (.Z(w3956), .A1(w3959), .B1(w3975), .A2(w3977), .B2(w4110) );
	vdp_slatch g4104 (.Q(w3979), .D(REG_BUS[1]), .C(w3967), .nC(w3966) );
	vdp_aon22 g4105 (.Z(w3960), .A1(w3952), .B1(w3975), .A2(w3977), .B2(w3979) );
	vdp_slatch g4106 (.Q(w4109), .D(REG_BUS[2]), .C(w3967), .nC(w3966) );
	vdp_aon22 g4107 (.Z(w3951), .A1(w3978), .B1(w3975), .A2(w3977), .B2(w4109) );
	vdp_slatch g4108 (.Q(w3980), .D(REG_BUS[3]), .C(w3967), .nC(w3966) );
	vdp_aon22 g4109 (.Z(w3945), .A1(w3944), .B1(w3975), .A2(w3977), .B2(w3980) );
	vdp_slatch g4110 (.Q(w3981), .D(REG_BUS[4]), .C(w3967), .nC(w3966) );
	vdp_aon22 g4111 (.Z(w3941), .A1(w3940), .B1(w3975), .A2(w3977), .B2(w3981) );
	vdp_slatch g4112 (.Q(w4007), .D(REG_BUS[5]), .C(w3967), .nC(w3966) );
	vdp_aon22 g4113 (.Z(w3939), .A1(w3932), .B1(w3975), .A2(w3977), .B2(w4007) );
	vdp_slatch g4114 (.Q(w4108), .D(REG_BUS[6]), .C(w3967), .nC(w3966) );
	vdp_aon22 g4115 (.Z(w3931), .A1(w3928), .B1(w3975), .A2(w3977), .B2(w4108) );
	vdp_slatch g4116 (.Q(w3982), .D(REG_BUS[7]), .C(w3967), .nC(w3966) );
	vdp_aon22 g4117 (.Z(w3929), .A1(w3925), .B1(w3975), .A2(w3977), .B2(w3982) );
	vdp_aon22 g4118 (.Z(w3936), .A1(w3983), .B1(w3975), .A2(w3977), .B2(1'b0) );
	vdp_aon22 g4119 (.Z(w3921), .A1(w3920), .B1(w3975), .A2(w3977), .B2(1'b0) );
	vdp_aon22 g4120 (.Z(w3998), .A1(w3915), .B1(w3975), .A2(w3977), .B2(1'b0) );
	vdp_notif0 g4121 (.nZ(RD_DATA[2]), .A(w3999), .nE(w3971) );
	vdp_slatch g4122 (.nQ(w3999), .D(w3915), .C(w3970), .nC(w3969) );
	vdp_notif0 g4123 (.nZ(RD_DATA[1]), .A(w3984), .nE(w3971) );
	vdp_slatch g4124 (.nQ(w3984), .D(w3920), .C(w3970), .nC(w3969) );
	vdp_notif0 g4125 (.nZ(RD_DATA[0]), .A(w4133), .nE(w3971) );
	vdp_slatch g4126 (.nQ(w4133), .D(w3983), .C(w3970), .nC(w3969) );
	vdp_notif0 g4127 (.nZ(AD_DATA[7]), .A(w4428), .nE(w3971) );
	vdp_slatch g4128 (.nQ(w4428), .D(w3925), .C(w3970), .nC(w3969) );
	vdp_notif0 g4129 (.nZ(AD_DATA[6]), .A(w3985), .nE(w3971) );
	vdp_slatch g4130 (.nQ(w3985), .D(w3928), .C(w3970), .nC(w3969) );
	vdp_notif0 g4131 (.nZ(AD_DATA[5]), .A(w3986), .nE(w3971) );
	vdp_slatch g4132 (.nQ(w3986), .D(w3932), .C(w3970), .nC(w3969) );
	vdp_notif0 g4133 (.nZ(AD_DATA[4]), .A(w3987), .nE(w3971) );
	vdp_slatch g4134 (.nQ(w3987), .D(w3940), .C(w3970), .nC(w3969) );
	vdp_notif0 g4135 (.nZ(AD_DATA[3]), .A(w3996), .nE(w3971) );
	vdp_slatch g4136 (.nQ(w3996), .D(w3944), .C(w3970), .nC(w3969) );
	vdp_notif0 g4137 (.nZ(AD_DATA[2]), .A(w3994), .nE(w3971) );
	vdp_slatch g4138 (.nQ(w3994), .D(w3978), .C(w3970), .nC(w3969) );
	vdp_notif0 g4139 (.nZ(AD_DATA[1]), .A(w3989), .nE(w3971) );
	vdp_slatch g4140 (.nQ(w3989), .D(w3952), .C(w3970), .nC(w3969) );
	vdp_notif0 g4141 (.nZ(AD_DATA[0]), .A(w3993), .nE(w3971) );
	vdp_slatch g4142 (.nQ(w3993), .D(w3959), .C(w3970), .nC(w3969) );
	vdp_sr_bit g4143 (.Q(w3992), .D(w3697), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4144 (.Q(w4000), .D(w4004), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4145 (.Q(w4004), .D(RD_DATA[0]), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4146 (.Q(w4132), .D(w3956), .C(w3916), .nC(w3911) );
	vdp_comp_strong g4147 (.Z(w3916), .nZ(w3911), .A(w3974) );
	vdp_comp_strong g4148 (.Z(w3910), .nZ(w3914), .A(w3972) );
	vdp_comp_strong g4149 (.Z(w3967), .nZ(w3966), .A(w87) );
	vdp_sr_bit g4150 (.Q(w3912), .D(w4113), .nC1(nHCLK1), .nC2(nHCLK2), .C2(HCLK2), .C1(HCLK1) );
	vdp_comp_strong g4151 (.Z(w3970), .nZ(w3969), .A(w3991) );
	vdp_not g4152 (.nZ(w3971), .A(w3992) );
	vdp_and g4153 (.Z(w3991), .A(w3697), .B(HCLK1) );
	vdp_and g4154 (.Z(w3927), .A(w4135), .B(w3912) );
	vdp_and g4155 (.Z(w3930), .A(w4134), .B(w3912) );
	vdp_and g4156 (.Z(w3937), .A(w4123), .B(w3912) );
	vdp_and g4157 (.Z(w3943), .A(w4124), .B(w3912) );
	vdp_and g4158 (.Z(w3946), .A(w4125), .B(w3912) );
	vdp_and g4159 (.Z(w3950), .A(w4126), .B(w3912) );
	vdp_and g4160 (.Z(w4010), .A(w4127), .B(w3912) );
	vdp_and g4161 (.Z(w3954), .A(w4132), .B(w3912) );
	vdp_not g4162 (.nZ(w4112), .A(w4111) );
	vdp_not g4163 (.nZ(w3972), .A(w3973) );
	vdp_not g4164 (.nZ(w3886), .A(w3885) );
	vdp_not g4165 (.nZ(w3890), .A(w3627) );
	vdp_not g4166 (.nZ(w3889), .A(w3632) );
	vdp_not g4167 (.nZ(w3867), .A(w4114) );
	vdp_not g4168 (.nZ(w3866), .A(w4115) );
	vdp_not g4169 (.nZ(w3868), .A(w4118) );
	vdp_not g4170 (.nZ(w4061), .A(M5) );
	vdp_not g4171 (.nZ(w3906), .A(w4060) );
	vdp_aon22 g4172 (.Z(w3894), .A1(w3873), .B1(w3881), .A2(w3900), .B2(w3876) );
	vdp_aon22 g4173 (.Z(w3898), .A1(w3873), .B1(w3900), .A2(w3897), .B2(w3876) );
	vdp_ha g4174 (.CO(w3902), .SUM(w3872), .B(w3901), .A(w3898) );
	vdp_aon222 g4175 (.A1(w3868), .B1(w3866), .C1(w3867), .A2(w3896), .B2(w3895), .C2(w3872), .Z(w3847) );
	vdp_aon22 g4176 (.Z(w4059), .A1(w3873), .B1(w3897), .A2(w3908), .B2(w3876) );
	vdp_ha g4177 (.SUM(w3871), .B(w3902), .A(w4059) );
	vdp_aon222 g4178 (.A1(w3868), .B1(w3866), .C1(w3867), .A2(w3895), .B2(w3872), .C2(w3871), .Z(w3849) );
	vdp_ha g4179 (.CO(w3901), .SUM(w3895), .B(w3894), .A(w3905) );
	vdp_aon222 g4180 (.A1(w3868), .B1(w3866), .C1(w3867), .A2(w3892), .B2(w3896), .C2(w3895), .Z(w3846) );
	vdp_aon22 g4181 (.Z(w3896), .A1(w3873), .B1(w3882), .A2(w3881), .B2(w3876) );
	vdp_aon222 g4182 (.A1(w3868), .B1(w3866), .C1(w3867), .A2(w4019), .B2(w3892), .C2(w3896), .Z(w3843) );
	vdp_aon222 g4183 (.A1(w3868), .B1(w3866), .C1(w3867), .A2(w3891), .B2(w3891), .C2(w3892), .Z(w3626) );
	vdp_aon22 g4184 (.Z(w3892), .A1(w3873), .B1(w3542), .A2(w3882), .B2(w3876) );
	vdp_comp_we g4185 (.Z(w3977), .nZ(w3975), .A(M5) );
	vdp_comp_we g4186 (.Z(w3873), .nZ(w3876), .A(w1) );
	vdp_and g4187 (.Z(w3905), .A(w3906), .B(w4061) );
	vdp_aon222 g4188 (.A1(w3868), .B1(w3866), .C1(w3867), .A2(w3872), .B2(w3871), .C2(w3869), .Z(w3854) );
	vdp_aon222 g4189 (.A1(w3868), .B1(w3866), .C1(w3867), .A2(w3871), .B2(w3869), .C2(w4058), .Z(w3865) );
	vdp_aon22 g4190 (.Z(w3870), .A1(w3873), .B1(w3874), .A2(w3875), .B2(w3876) );
	vdp_aon22 g4191 (.Z(w3893), .A1(w3873), .B1(w3908), .A2(w3874), .B2(w3876) );
	vdp_and g4192 (.Z(w3869), .B(w3893), .A(w3903) );
	vdp_and g4193 (.Z(w4058), .B(w3870), .A(w3904) );
	vdp_oai21 g4194 (.Z(w3885), .A1(w44), .A2(w3957), .B(M5) );
	vdp_aoi21 g4195 (.Z(w3973), .A1(HCLK1), .A2(w16), .B(w103) );
	vdp_oai211 g4196 (.Z(w4111), .A1(HCLK1), .A2(w4), .B(w5), .C(M5) );
	vdp_or g4197 (.Z(w3974), .A(w103), .B(w4112) );
	vdp_nand3 g4198 (.Z(w4113), .A(w95), .B(HPOS[6]), .C(HPOS[7]) );
	vdp_nand g4199 (.Z(w4118), .A(w3632), .B(w3627) );
	vdp_nand g4200 (.Z(w4115), .A(w3627), .B(w3889) );
	vdp_nand g4201 (.Z(w4114), .A(w3889), .B(w3890) );
	vdp_aoi31 g4202 (.Z(w4060), .B3(w4059), .B2(w3898), .B1(w3894), .A(w3893) );
	vdp_slatch g4203 (.Q(w3575), .D(S[0]), .C(w3537), .nC(w3152) );
	vdp_slatch g4204 (.Q(w3577), .D(S[1]), .C(w3537), .nC(w3152) );
	vdp_slatch g4205 (.Q(w3597), .D(S[2]), .C(w3537), .nC(w3152) );
	vdp_slatch g4206 (.Q(w3581), .D(S[3]), .C(w3537), .nC(w3152) );
	vdp_slatch g4207 (.Q(w3583), .D(S[4]), .C(w3537), .nC(w3152) );
	vdp_slatch g4208 (.Q(w3584), .D(S[5]), .C(w3537), .nC(w3152) );
	vdp_slatch g4209 (.Q(w3586), .D(S[6]), .C(w3537), .nC(w3152) );
	vdp_slatch g4210 (.Q(w3588), .D(S[7]), .C(w3537), .nC(w3152) );
	vdp_slatch g4211 (.Q(w3590), .D(S[0]), .C(w3532), .nC(w3531) );
	vdp_slatch g4212 (.Q(w3593), .D(S[1]), .C(w3532), .nC(w3531) );
	vdp_slatch g4213 (.Q(w3594), .D(S[2]), .C(w3532), .nC(w3531) );
	vdp_slatch g4214 (.Q(w3100), .D(S[3]), .C(w3532), .nC(w3531) );
	vdp_slatch g4215 (.Q(w3601), .D(S[4]), .C(w3532), .nC(w3531) );
	vdp_slatch g4216 (.Q(w3076), .D(S[5]), .C(w3532), .nC(w3531) );
	vdp_slatch g4217 (.Q(w3078), .D(S[6]), .C(w3532), .nC(w3531) );
	vdp_slatch g4218 (.Q(w3105), .D(S[7]), .C(w3532), .nC(w3531) );
	vdp_comp_strong g4219 (.Z(w3532), .nZ(w3531), .A(w3287) );
	vdp_comp_strong g4220 (.Z(w3537), .nZ(w3152), .A(w3288) );
	vdp_comp_strong g4221 (.Z(w3538), .nZ(w3599), .A(w3289) );
	vdp_slatch g4222 (.Q(w4093), .D(S[7]), .C(w3538), .nC(w3599) );
	vdp_slatch g4223 (.Q(w4092), .D(S[6]), .C(w3538), .nC(w3599) );
	vdp_slatch g4224 (.Q(w4091), .D(S[5]), .C(w3538), .nC(w3599) );
	vdp_slatch g4225 (.Q(w3604), .D(S[4]), .C(w3538), .nC(w3599) );
	vdp_slatch g4226 (.Q(w3605), .D(S[3]), .C(w3538), .nC(w3599) );
	vdp_slatch g4227 (.Q(w3570), .D(S[2]), .C(w3538), .nC(w3599) );
	vdp_slatch g4228 (.Q(w3568), .D(S[1]), .C(w3538), .nC(w3599) );
	vdp_slatch g4229 (.Q(w3566), .D(S[0]), .C(w3538), .nC(w3599) );
	vdp_slatch g4230 (.Q(w3563), .D(S[7]), .C(w3539), .nC(w3600) );
	vdp_slatch g4231 (.Q(w3564), .D(S[6]), .C(w3539), .nC(w3600) );
	vdp_slatch g4232 (.Q(w3562), .D(S[5]), .C(w3539), .nC(w3600) );
	vdp_slatch g4233 (.Q(w3561), .D(S[4]), .C(w3539), .nC(w3600) );
	vdp_slatch g4234 (.Q(w3559), .D(S[3]), .C(w3539), .nC(w3600) );
	vdp_slatch g4235 (.Q(w3557), .D(S[2]), .C(w3539), .nC(w3600) );
	vdp_slatch g4236 (.Q(w3555), .D(S[1]), .C(w3539), .nC(w3600) );
	vdp_slatch g4237 (.Q(w3552), .D(S[0]), .C(w3539), .nC(w3600) );
	vdp_sr_bit g4238 (.Q(w4122), .D(w3533), .C1(HCLK2), .C2(HCLK1), .nC2(nHCLK1), .nC1(nHCLK2) );
	vdp_sr_bit g4239 (.Q(w3540), .D(w4090), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_and g4240 (.Z(w4090), .A(w14), .B(M5) );
	vdp_not g4241 (.nZ(w4088), .A(w3540) );
	vdp_aon22 g4242 (.Z(w3104), .A1(w4093), .B1(w3604), .A2(w3603), .B2(w4051) );
	vdp_aon22 g4243 (.Z(w3101), .A1(w4092), .B1(1'b0), .A2(w3603), .B2(w4051) );
	vdp_aon22 g4244 (.Z(w3602), .A1(w3604), .B1(w3570), .A2(w3603), .B2(w4051) );
	vdp_aon22 g4245 (.Z(w3074), .A1(w3605), .B1(w3568), .A2(w3603), .B2(w4051) );
	vdp_aon22 g4246 (.Z(w3077), .A1(w4091), .B1(w3605), .A2(w3603), .B2(w4051) );
	vdp_comp_strong g4247 (.Z(w3539), .nZ(w3600), .A(w3290) );
	vdp_comp_we g4248 (.Z(w3603), .nZ(w4051), .A(M5) );
	vdp_aon22 g4249 (.Z(w3544), .A1(w3601), .B1(w3602), .A2(w3540), .B2(w4088) );
	vdp_sr_bit g4250 (.Q(w4001), .D(FIFOo[0]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4251 (.Q(w4005), .D(FIFOo[1]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4252 (.Q(w4003), .D(FIFOo[2]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4253 (.Q(w4002), .D(FIFOo[3]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4254 (.Q(w3990), .D(FIFOo[4]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4255 (.Q(w3988), .D(FIFOo[5]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4256 (.Q(w3995), .D(FIFOo[6]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_sr_bit g4257 (.Q(w3997), .D(FIFOo[7]), .C1(HCLK1), .C2(HCLK2), .nC2(nHCLK2), .nC1(nHCLK1) );
	vdp_aon22 g4258 (.Z(w1409), .B1(w4471), .A1(w1437), .B2(w4489), .A2(w43) );
	vdp_not g4259 (.nZ(w4489), .A(w43) );
	vdp_not g4260 (.nZ(w4461), .A(w4448) );
	vdp_not g4261 (.nZ(w4460), .A(w4461) );
	vdp_not g4262 (.nZ(w4459), .A(w4460) );
	vdp_not g4263 (.nZ(w4458), .A(w4459) );
	vdp_and g4264 (.Z(w4471), .B(w4462), .A(w4466) );
	vdp_not g4265 (.nZ(w4462), .A(w4465) );
	vdp_not g4266 (.nZ(w4465), .A(w4464) );
	vdp_not g4267 (.nZ(w4464), .A(w4463) );
	vdp_not g4268 (.nZ(w4463), .A(w4466) );
	vdp_or g4269 (.Z(w4466), .B(w4446), .A(w4445) );
	vdp_dff g4270 (.Q(w4446), .R(w4435), .D(w4445), .C(w4444) );
	vdp_not g4271 (.nZ(w4444), .A(w4467) );
	vdp_nor g4272 (.Z(w4443), .B(w4468), .A(w4445) );
	vdp_dff g4273 (.Q(w4445), .R(w4435), .D(w4468), .C(w4467) );
	vdp_dff g4274 (.Q(w4468), .R(w4435), .D(w4443), .C(w4467) );
	vdp_not g4275 (.nZ(w4467), .A(w4454) );
	vdp_not g4276 (.nZ(w4441), .A(w4454) );
	vdp_dff g4277 (.Q(w4438), .R(w4435), .D(w4469), .C(w4437) );
	vdp_dff g4278 (.Q(w4469), .R(w4435), .D(w4436), .C(w4434) );
	vdp_not g4279 (.nZ(w4434), .A(w4477) );
	vdp_dff g4280 (.Q(w4436), .R(w4435), .D(w4455), .C(w4434) );
	vdp_not g4281 (.nZ(w4437), .A(w4434) );
	vdp_nor g4282 (.Z(w4496), .B(w4472), .A(w4473) );
	vdp_nor g4283 (.Z(w4474), .B(w4472), .A(H40) );
	vdp_not g4284 (.nZ(w4473), .A(H40) );
	vdp_not g4285 (.nZ(w4449), .A(PAL) );
	vdp_AOI222 g4286 (.Z(w4442), .B1(w4476), .A1(w4475), .B2(w4496), .A2(w4472), .C1(w4441), .C2(w4474) );
	vdp_not g4287 (.nZ(EDCLK_O), .A(w4442) );
	vdp_or g4288 (.Z(w4470), .B(w4438), .A(w4469) );
	vdp_nor g4289 (.Z(w4455), .B(w4436), .A(w4469) );
	vdp_not g4290 (.nZ(w4431), .A(w4495) );
	vdp_nand g4291 (.Z(w4450), .B(w4431), .A(w4430) );
	vdp_SR_bit g4292 (.Q(w4495), .D(w4430), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_not g4293 (.nZ(w4494), .A(w4480) );
	vdp_not g4294 (.nZ(w1167), .A(w4493) );
	vdp_not g4295 (.nZ(SYSRES), .A(w4494) );
	vdp_comp_DFF g4296 (.Q(w4430), .D(w4480), .C1(DCLK1), .C2(DCLK2), .nC1(nDCLK1), .nC2(nDCLK2) );
	vdp_not g4297 (.nZ(w4490), .A(w4491) );
	vdp_not g4298 (.nZ(w4435), .A(w4492) );
	vdp_not g4299 (.nZ(w4479), .A(w4478) );
	vdp_nand g4300 (.Z(w4492), .B(w4479), .A(w4433) );
	vdp_not g4301 (.nZ(w4477), .A(w4481) );
	vdp_nand g4302 (.Z(w4484), .B(w4483), .A(w4482) );
	vdp_not g4303 (.nZ(w4454), .A(w4439) );
	vdp_nand g4304 (.Z(w4487), .B(w4486), .A(w4485) );
	vdp_not g4305 (.nZ(w4448), .A(w4453) );
	vdp_not g4306 (.nZ(RES), .A(w4450) );
	vdp_dff g4307 (.Q(w4433), .R(1'b0), .D(w4480), .C(w4451) );
	vdp_dff g4308 (.Q(w4478), .R(1'b0), .D(w4433), .C(w4451) );
	vdp_dff g4309 (.Q(w4491), .R(w4435), .D(w4481), .C(w4451) );
	vdp_dff g4310 (.Q(w4481), .R(w4435), .D(w4490), .C(w4451) );
	vdp_dff g4311 (.Q(w4482), .R(w4435), .D(w4439), .C(w4451) );
	vdp_dff g4312 (.Q(w4483), .R(w4435), .D(w4482), .C(w4451) );
	vdp_dff g4313 (.Q(w4439), .R(w4435), .D(w4484), .C(w4451) );
	vdp_dff g4314 (.Q(w4485), .R(w4435), .D(w4453), .C(w4451) );
	vdp_dff g4315 (.Q(w4486), .R(w4435), .D(w4485), .C(w4451) );
	vdp_dff g4316 (.Q(w4488), .R(w4435), .D(w4487), .C(w4451) );
	vdp_dff g4317 (.Q(w4453), .R(w4435), .D(w4488), .C(w4451) );
	vdp_not g4318 (.nZ(w4476), .A(w4477) );
	vdp_nand g4319 (.Z(w4480), .B(w1438), .A(w4493) );
	vdp_not g4320 (.nZ(68K CPU CLOCK), .A(w4447) );
	vdp_or g4321 (.Z(w4472), .B(w43), .A(w1148) );
	vdp_aon22 g4322 (.Z(w4440), .B1(w4470), .A1(w4471), .B2(PAL), .A2(w4449) );
	vdp_or g4323 (.Z(w4447), .B(w4458), .A(w4448) );
	vdp_comp_we g4324 (.A(w2634), .nZ(nHCLK2), .Z(HCLK2) );
	vdp_comp_we g4325 (.A(w2633), .nZ(nHCLK1), .Z(HCLK1) );
	vdp_comp_we g4326 (.A(w4504), .nZ(nDCLK2), .Z(DCLK2) );
	vdp_comp_we g4327 (.A(EDCLK_O), .nZ(nDCLK1), .Z(DCLK1) );
	vdp_not g4328 (.nZ(w4504), .A(EDCLK_O) );
	vdp_sr_bit g4329 (.Q(w4602), .D(w4601), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4330 (.Q(w4620), .D(w4597), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4331 (.Q(w4597), .D(w4582), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4332 (.Q(w4582), .D(w4574), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4333 (.Q(w4577), .D(w6552), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4334 (.Q(w6552), .D(w6553), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4335 (.Q(w6553), .D(w6555), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4336 (.Q(w6555), .D(w6554), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4337 (.Q(w6554), .D(w6556), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4338 (.Q(w6556), .D(w6557), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4339 (.Q(w6557), .D(w6559), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4340 (.Q(w6559), .D(w6558), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4341 (.Q(w6558), .D(w6385), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4342 (.Q(w6385), .D(w4520), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4343 (.Q(w4558), .D(w4559), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4344 (.Q(w4559), .D(w24), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4345 (.Q(w4556), .D(w6560), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4346 (.Q(w4525), .D(w4555), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4347 (.Q(w4524), .D(w6548), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4348 (.Q(w6248), .D(w4604), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4349 (.Q(w4603), .D(w6561), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4350 (.Q(w4605), .D(w4595), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4351 (.Q(w6550), .D(w4), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4352 (.Q(w4545), .D(w4567), .nC(w4570), .C(w4571) );
	vdp_slatch g4353 (.Q(w4549), .D(w4568), .nC(w4570), .C(w4571) );
	vdp_slatch g4354 (.Q(w4537), .D(w4569), .nC(w4570), .C(w4571) );
	vdp_slatch g4355 (.Q(w4528), .D(w4575), .nC(w4570), .C(w4571) );
	vdp_slatch g4356 (.Q(w4527), .D(w4566), .nC(w4570), .C(w4571) );
	vdp_slatch g4357 (.Q(w4526), .D(w4565), .nC(w4570), .C(w4571) );
	vdp_slatch g4358 (.Q(w4579), .D(w4564), .nC(w4570), .C(w4571) );
	vdp_slatch g4359 (.Q(w4529), .D(w4562), .nC(w4570), .C(w4571) );
	vdp_slatch g4360 (.Q(w4533), .D(w4563), .nC(w4570), .C(w4571) );
	vdp_slatch g4361 (.Q(w4534), .D(w4561), .nC(w4570), .C(w4571) );
	vdp_comp_str g4362 (.nZ(w4570), .A(w4576), .Z(w4571) );
	vdp_sr_bit g4363 (.Q(w4598), .D(w4621), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4364 (.Q(w6234), .D(w7), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_xor g4365 (.Z(w4543), .B(w4535), .A(w4546) );
	vdp_xor g4366 (.Z(w4538), .B(w4536), .A(w4544) );
	vdp_xor g4367 (.Z(w4540), .B(w4522), .A(w4537) );
	vdp_xor g4368 (.Z(w6337), .B(w4522), .A(w4528) );
	vdp_xor g4369 (.Z(w6338), .B(w4522), .A(w4527) );
	vdp_xor g4370 (.Z(w6333), .B(w4522), .A(w4526) );
	vdp_aon22 g4371 (.Z(w6334), .B2(w4550), .B1(w4545), .A1(w4543), .A2(w4539) );
	vdp_aon22 g4372 (.Z(w6335), .B2(w4550), .B1(w4543), .A1(w4538), .A2(w4539) );
	vdp_aon22 g4373 (.Z(w6336), .B2(w4550), .B1(w4538), .A1(w4540), .A2(w4539) );
	vdp_aon22 g4374 (.Z(w4541), .B2(w4532), .B1(w4537), .A1(w4549), .A2(w4542) );
	vdp_aon22 g4375 (.Z(w4547), .B2(w4532), .B1(w4549), .A1(w4545), .A2(w4542) );
	vdp_aon22 g4376 (.Z(w4613), .B2(w4606), .B1(w4609), .A1(w4610), .A2(w80) );
	vdp_aon22 g4377 (.Z(w4614), .B2(w4608), .B1(w4609), .A1(w4610), .A2(w79) );
	vdp_aon22 g4378 (.Z(w4615), .B2(w4607), .B1(w4609), .A1(w4610), .A2(w78) );
	vdp_aon22 g4379 (.Z(w4616), .B2(w4611), .B1(w4609), .A1(w4610), .A2(w77) );
	vdp_aon22 g4380 (.Z(w4617), .B2(w4612), .B1(w4609), .A1(w4610), .A2(w76) );
	vdp_not g4381 (.nZ(w4583), .A(w4520) );
	vdp_not g4382 (.nZ(w4553), .A(w4587) );
	vdp_not g4383 (.nZ(w4586), .A(w125) );
	vdp_not g4384 (.nZ(w4591), .A(w4589) );
	vdp_not g4385 (.nZ(w4578), .A(M5) );
	vdp_not g4386 (.nZ(w4619), .A(w81) );
	vdp_not g4387 (.nZ(w4618), .A(w82) );
	vdp_not g4388 (.nZ(w4593), .A(1'b0) );
	vdp_not g4389 (.nZ(w4594), .A(M5) );
	vdp_not g4390 (.nZ(w4519), .A(w4520) );
	vdp_not g4391 (.nZ(w4523), .A(w4554) );
	vdp_not g4392 (.nZ(w4530), .A(w4534) );
	vdp_not g4393 (.nZ(w4536), .A(w4573) );
	vdp_and g4394 (.Z(w4574), .B(w4583), .A(w4584) );
	vdp_and g4395 (.Z(w4588), .B(w4586), .A(w4597) );
	vdp_or g4396 (.Z(w4585), .B(w4588), .A(w4600) );
	vdp_or g4397 (.Z(w4581), .B(w4623), .A(w4588) );
	vdp_and g4398 (.Z(w4599), .B(w4592), .A(1'b0) );
	vdp_and g4399 (.Z(w4622), .B(w4592), .A(w4593) );
	vdp_or g4400 (.Z(w4621), .B(w7), .A(w27) );
	vdp_and g4401 (.Z(w127), .B(w6709), .A(w4) );
	vdp_and g4402 (.Z(w6548), .B(w4519), .A(w4521) );
	vdp_or g4403 (.Z(w4572), .B(w4525), .A(w4524) );
	vdp_and g4404 (.Z(w4535), .B(w4529), .A(w4522) );
	vdp_comp_we g4405 (.nZ(w4532), .A(w1), .Z(w4542) );
	vdp_comp_we g4406 (.nZ(w4550), .A(w1), .Z(w4539) );
	vdp_comp_we g4407 (.nZ(w4609), .A(w125), .Z(w4610) );
	vdp_not g4408 (.nZ(w4631), .A(w4601) );
	vdp_rs_FF g4409 (.Q(w6549), .R(w6550), .S(w4572) );
	vdp_rs_FF g4410 (.Q(w6709), .R(w6550), .S(w4524) );
	vdp_ha g4411 (.SUM(w4546), .B(w4547), .A(w4548) );
	vdp_ha g4412 (.SUM(w4544), .B(w4541), .A(w4531), .CO(w4548) );
	vdp_not g4413 (.nZ(w4557), .A(w4518) );
	vdp_and g4414 (.Z(w4560), .B(w4520), .A(w4521) );
	vdp_and3 g4415 (.Z(w4531), .B(w4529), .A(w4522), .C(w4530) );
	vdp_and3 g4416 (.Z(w4604), .B(w4602), .A(M5), .C(w4631) );
	vdp_and3 g4417 (.Z(w6561), .B(w4607), .A(w4606), .C(w4605) );
	vdp_and3 g4418 (.Z(w4623), .B(w82), .A(w4619), .C(w118) );
	vdp_and3 g4419 (.Z(w6551), .B(w81), .A(w4618), .C(w118) );
	vdp_and3 g4420 (.Z(w4600), .B(w4619), .A(w4618), .C(w118) );
	vdp_or3 g4421 (.Z(w4580), .B(w6551), .A(w4588), .C(w4591) );
	vdp_and3 g4422 (.Z(w4576), .B(HCLK1), .A(w4558), .C(DCLK1) );
	vdp_or3 g4423 (.Z(w4592), .B(w4595), .A(w4620), .C(w4594) );
	vdp_oai21 g4424 (.Z(w4573), .B(w4522), .A1(w4529), .A2(w4534) );
	vdp_nor g4425 (.Z(w4518), .B(w4560), .A(w4559) );
	vdp_nor g4426 (.Z(w6560), .B(w4523), .A(w6549) );
	vdp_nand g4427 (.Z(w4596), .B(w4578), .A(w4577) );
	vdp_nand g4428 (.Z(w4552), .B(w4619), .A(w4618) );
	vdp_nand g4429 (.Z(w4587), .B(w81), .A(w4618) );
	vdp_nand g4430 (.Z(w4551), .B(w82), .A(w4619) );
	vdp_nor g4431 (.Z(w4601), .B(w4603), .A(w4516) );
	vdp_cnt_bit_rev g4432 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4606), .CI(w4635), .B(w4598), .A(w4599) );
	vdp_cnt_bit_rev g4433 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4608), .CI(w4634), .B(w4598), .A(w4599), .CO(w4635) );
	vdp_cnt_bit_rev g4434 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4607), .CI(w4633), .B(w4598), .A(w4599), .CO(w4634) );
	vdp_cnt_bit_rev g4435 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4611), .CI(w4632), .B(w4598), .A(w4599), .CO(w4633) );
	vdp_cnt_bit_rev g4436 (.nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .Q(w4612), .CI(w4622), .B(w4598), .A(w4599), .CO(w4632) );
	vdp_cnt_bit_load g4437 (.Q(w4642), .D(w4682), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4644), .CI(w6612), .L(w4683), .nL(w4648) );
	vdp_cnt_bit_load g4438 (.Q(w4645), .D(w4687), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4644), .CI(w6611), .L(w4683), .nL(w4648), .CO(w6612) );
	vdp_cnt_bit_load g4439 (.Q(w4647), .D(w4688), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4644), .CI(w6610), .L(w4683), .nL(w4648), .CO(w6611) );
	vdp_cnt_bit_load g4440 (.Q(w4649), .D(w4712), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4644), .CI(w6609), .L(w4683), .nL(w4648), .CO(w6610) );
	vdp_cnt_bit_load g4441 (.Q(w4653), .D(w4713), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4644), .CI(w6608), .L(w4683), .nL(w4648), .CO(w6609) );
	vdp_cnt_bit_load g4442 (.Q(w4650), .D(w4714), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4644), .CI(w6607), .L(w4683), .nL(w4648), .CO(w6608) );
	vdp_cnt_bit_load g4443 (.Q(w4646), .D(w4715), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w4644), .CI(w4643), .L(w4683), .nL(w4648), .CO(w6607) );
	vdp_fa g4444 (.SUM(w4790), .CO(w6622), .CI(1'b1), .A(w4844), .B(w4793) );
	vdp_fa g4445 (.SUM(w4792), .CO(w6623), .CI(w6622), .A(w4843), .B(w4797) );
	vdp_fa g4446 (.SUM(w4798), .CO(w6624), .CI(w6623), .A(w4842), .B(w4801) );
	vdp_fa g4447 (.SUM(w4800), .CO(w6625), .CI(w6624), .A(w4841), .B(w4803) );
	vdp_fa g4448 (.SUM(w4805), .CO(w6626), .CI(w6625), .A(w4840), .B(w4807) );
	vdp_fa g4449 (.SUM(w4811), .CO(w6627), .CI(w6626), .A(w4839), .B(w4835) );
	vdp_fa g4450 (.SUM(w4814), .CO(w6628), .CI(w6627), .A(w4837), .B(w4813) );
	vdp_fa g4451 (.SUM(w4818), .CO(w6629), .CI(w6628), .A(w4849), .B(w4817) );
	vdp_fa g4452 (.SUM(w4820), .CO(w6630), .CI(w6629), .A(w4850), .B(w4819) );
	vdp_fa g4453 (.SUM(w4833), .CI(w6630), .A(w4854), .B(w4832) );
	vdp_fa g4454 (.SUM(w4844), .CO(w6613), .CI(1'b0), .A(VPOS[0]), .B(w4845) );
	vdp_fa g4455 (.SUM(w4843), .CO(w6614), .CI(w6613), .A(VPOS[1]), .B(w1) );
	vdp_fa g4456 (.SUM(w4842), .CO(w6615), .CI(w6614), .A(VPOS[2]), .B(1'b0) );
	vdp_fa g4457 (.SUM(w4841), .CO(w6616), .CI(w6615), .A(VPOS[3]), .B(1'b0) );
	vdp_fa g4458 (.SUM(w4840), .CO(w6617), .CI(w6616), .A(VPOS[4]), .B(1'b0) );
	vdp_fa g4459 (.SUM(w4839), .CO(w6618), .CI(w6617), .A(VPOS[5]), .B(1'b0) );
	vdp_fa g4460 (.SUM(w4837), .CO(w6619), .CI(w6618), .A(VPOS[6]), .B(1'b0) );
	vdp_fa g4461 (.SUM(w4849), .CO(w6620), .CI(w6619), .A(VPOS[7]), .B(w4845) );
	vdp_fa g4462 (.SUM(w4850), .CO(w6621), .CI(w6620), .A(VPOS[8]), .B(w1) );
	vdp_fa g4463 (.SUM(w4854), .CI(w6621), .A(VPOS[9]), .B(1'b0) );
	vdp_slatch g4464 (.nC(w4738), .C(w4737), .Q(w4784), .D(S[0]) );
	vdp_dlatch_inv g4465 (.nQ(w4783), .D(w4751), .nC(nHCLK2), .C(HCLK2) );
	vdp_slatch g4466 (.nC(w4723), .C(w4722), .Q(w4751), .D(w4740) );
	vdp_slatch g4467 (.nC(w4738), .C(w4737), .Q(w4781), .D(S[1]) );
	vdp_slatch g4468 (.nC(w4723), .C(w4722), .Q(w6652), .D(w4742) );
	vdp_slatch g4469 (.nC(w4738), .C(w4737), .Q(w4779), .D(S[2]) );
	vdp_slatch g4470 (.nC(w4723), .C(w4722), .Q(w6653), .D(w4733) );
	vdp_slatch g4471 (.nC(w4738), .C(w4737), .Q(w4777), .D(S[3]) );
	vdp_slatch g4472 (.nC(w4723), .C(w4722), .Q(w6654), .D(w4729) );
	vdp_slatch g4473 (.nC(w4738), .C(w4737), .Q(w4773), .D(S[4]) );
	vdp_slatch g4474 (.nC(w4723), .C(w4722), .Q(w6655), .D(w4725) );
	vdp_slatch g4475 (.nC(w4738), .C(w4737), .Q(w4772), .D(S[5]) );
	vdp_slatch g4476 (.nC(w4723), .C(w4722), .Q(w6656), .D(w4721) );
	vdp_slatch g4477 (.nC(w4738), .C(w4737), .Q(w4769), .D(S[6]) );
	vdp_slatch g4478 (.nC(w4723), .C(w4722), .Q(w6657), .D(w6599) );
	vdp_slatch g4479 (.nC(w4738), .C(w4737), .Q(w6658), .D(S[7]) );
	vdp_slatch g4480 (.nC(w4723), .C(w4722), .Q(w6659), .D(w4753) );
	vdp_slatch g4481 (.nC(w4723), .C(w4722), .Q(w4754), .D(w4755) );
	vdp_slatch g4482 (.nC(w4723), .C(w4722), .Q(w6660), .D(w4757) );
	vdp_dlatch_inv g4483 (.nQ(w4780), .D(w6652), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4484 (.nQ(w4778), .D(w6653), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4485 (.nQ(w4775), .D(w6654), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4486 (.nQ(w4774), .D(w6655), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4487 (.nQ(w4771), .D(w6656), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4488 (.nQ(w4768), .D(w6657), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4489 (.nQ(w4767), .D(w6659), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4490 (.nQ(w4766), .D(w4754), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4491 (.nQ(w4756), .D(w6660), .nC(nHCLK2), .C(HCLK2) );
	vdp_sr_bit g4492 (.Q(w4708), .D(w4639), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4493 (.Z(w4554), .B2(w4704), .B1(w4710), .A1(M5), .A2(w4709) );
	vdp_sr_bit g4494 (.Q(w4639), .D(w4705), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4495 (.Q(w6598), .D(w4706), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4496 (.Q(w4706), .D(w4684), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4497 (.Q(w4745), .D(w4747), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4498 (.Q(w4736), .D(w4750), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4499 (.Q(w4732), .D(w4743), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4500 (.Q(w4728), .D(w4744), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4501 (.Q(w4724), .D(w4726), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4502 (.Q(w4720), .D(w4718), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4503 (.Q(w4752), .D(w4719), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4504 (.Q(w6661), .D(w4717), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4505 (.Q(w4666), .D(w4716), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4506 (.Q(w4673), .D(w4711), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4507 (.Q(w4707), .D(w4640), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4508 (.Q(w4640), .D(w4662), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4509 (.Q(w4890), .D(w131), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4510 (.Q(w4892), .D(VRAMA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4511 (.Q(w4662), .D(w9), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4512 (.Q(w4893), .D(w6606), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4513 (.Q(w6606), .D(w4890), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4514 (.Q(w6650), .D(w4876), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4515 (.Q(w6648), .D(w4879), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4516 (.Q(w6646), .D(w4894), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4517 (.Q(w6644), .D(w4856), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4518 (.Q(w6642), .D(w4682), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4519 (.Q(w6640), .D(w4687), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4520 (.Q(w6638), .D(w4688), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4521 (.Q(w6636), .D(w4712), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4522 (.Q(w6634), .D(w4713), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4523 (.Q(w6632), .D(w4714), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4524 (.Q(w4874), .D(w4715), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_slatch g4525 (.Q(w4866), .D(w6631), .nC(w4865), .C(w4857) );
	vdp_dlatch_inv g4526 (.nQ(w6631), .D(w4874), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4527 (.Q(w4867), .D(w6633), .nC(w4865), .C(w4857) );
	vdp_dlatch_inv g4528 (.nQ(w6633), .D(w6632), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4529 (.Q(w4868), .D(w6635), .nC(w4865), .C(w4857) );
	vdp_dlatch_inv g4530 (.nQ(w6635), .D(w6634), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4531 (.Q(w4869), .D(w6637), .nC(w4865), .C(w4857) );
	vdp_dlatch_inv g4532 (.nQ(w6637), .D(w6636), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4533 (.Q(w4870), .D(w6639), .nC(w4865), .C(w4857) );
	vdp_dlatch_inv g4534 (.nQ(w6639), .D(w6638), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4535 (.Q(w6605), .D(w6641), .nC(w4865), .C(w4857) );
	vdp_dlatch_inv g4536 (.nQ(w6641), .D(w6640), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4537 (.Q(w4871), .D(w6643), .nC(w4865), .C(w4857) );
	vdp_dlatch_inv g4538 (.nQ(w6643), .D(w6642), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4539 (.Q(w4861), .D(w6645), .nC(w4865), .C(w4857) );
	vdp_dlatch_inv g4540 (.nQ(w6645), .D(w6644), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4541 (.Q(w4864), .D(w6647), .nC(w4865), .C(w4857) );
	vdp_dlatch_inv g4542 (.nQ(w6647), .D(w6646), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4543 (.Q(w4862), .D(w6649), .nC(w4865), .C(w4857) );
	vdp_dlatch_inv g4544 (.nQ(w6649), .D(w6648), .nC(nHCLK1), .C(HCLK1) );
	vdp_slatch g4545 (.Q(w4863), .D(w6651), .nC(w4865), .C(w4857) );
	vdp_dlatch_inv g4546 (.nQ(w6651), .D(w6650), .nC(nHCLK1), .C(HCLK1) );
	vdp_aon22 g4547 (.Z(w6404), .B2(w4692), .B1(w4642), .A1(w4641), .A2(w6383) );
	vdp_aon22 g4548 (.Z(w6405), .B2(w4692), .B1(w4645), .A1(w4641), .A2(w4697) );
	vdp_aon22 g4549 (.Z(w6406), .B2(w4692), .B1(w4647), .A1(w4641), .A2(w4696) );
	vdp_aon22 g4550 (.Z(w6407), .B2(w4692), .B1(w4649), .A1(w4641), .A2(w4695) );
	vdp_aon22 g4551 (.Z(w6408), .B2(w4692), .B1(w4653), .A1(w4641), .A2(w4694) );
	vdp_aon22 g4552 (.Z(w6410), .B2(w4692), .B1(w4650), .A1(w4641), .A2(w4693) );
	vdp_aon22 g4553 (.Z(w6409), .B2(w4692), .B1(w4646), .A1(w4641), .A2(w4691) );
	vdp_aon22 g4554 (.Z(w4915), .B2(w4655), .B1(w3), .A1(w4651), .A2(w4646) );
	vdp_aon22 g4555 (.Z(w4804), .B2(w4764), .B1(w4773), .A1(w4774), .A2(w4788) );
	vdp_2x_sr_bit g4556 (.Q(w4703), .D(w4646), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4557 (.Z(w6384), .B2(w4655), .B1(w4703), .A1(w4651), .A2(w4650) );
	vdp_2x_sr_bit g4558 (.Q(w4652), .D(w4650), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4559 (.Z(w4972), .B2(w4655), .B1(w4652), .A1(w4651), .A2(w4653) );
	vdp_2x_sr_bit g4560 (.Q(w4690), .D(w4653), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4561 (.Z(w4978), .B2(w4655), .B1(w4690), .A1(w4651), .A2(w4649) );
	vdp_2x_sr_bit g4562 (.Q(w4654), .D(w4649), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4563 (.Z(w5028), .B2(w4655), .B1(w4654), .A1(w4651), .A2(w4647) );
	vdp_2x_sr_bit g4564 (.Q(w4657), .D(w4647), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .nC4(nHCLK2), .nC3(nHCLK1), .C4(HCLK2), .C3(HCLK1) );
	vdp_aon22 g4565 (.Z(w5080), .B2(w4655), .B1(w4657), .A1(w4651), .A2(w4645) );
	vdp_aon22 g4566 (.Z(w5095), .B2(w4655), .B1(1'b1), .A1(w4651), .A2(w4642) );
	vdp_aon22 g4567 (.Z(w4740), .B2(w4665), .B1(w4741), .A1(w4668), .A2(w4739) );
	vdp_dlatch_inv g4568 (.nQ(w4739), .D(w4745), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4569 (.nZ(w4741), .A(S[0]) );
	vdp_aon22 g4570 (.Z(w4742), .B2(w4665), .B1(w4735), .A1(w4668), .A2(w4734) );
	vdp_dlatch_inv g4571 (.nQ(w4734), .D(w4736), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4572 (.nZ(w4735), .A(S[1]) );
	vdp_aon22 g4573 (.Z(w4733), .B2(w4665), .B1(w4731), .A1(w4668), .A2(w4730) );
	vdp_dlatch_inv g4574 (.nQ(w4730), .D(w4732), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4575 (.nZ(w4731), .A(S[2]) );
	vdp_aon22 g4576 (.Z(w4729), .B2(w4665), .B1(w4689), .A1(w4668), .A2(w4727) );
	vdp_dlatch_inv g4577 (.nQ(w4727), .D(w4728), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4578 (.nZ(w4689), .A(S[3]) );
	vdp_aon22 g4579 (.Z(w4725), .B2(w4665), .B1(w4685), .A1(w4668), .A2(w4686) );
	vdp_dlatch_inv g4580 (.nQ(w4686), .D(w4724), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4581 (.nZ(w4685), .A(S[4]) );
	vdp_aon22 g4582 (.Z(w4721), .B2(w4665), .B1(w4681), .A1(w4668), .A2(w4680) );
	vdp_dlatch_inv g4583 (.nQ(w4680), .D(w4720), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4584 (.nZ(w4681), .A(S[5]) );
	vdp_aon22 g4585 (.Z(w6599), .B2(w4665), .B1(w4676), .A1(w4668), .A2(w4675) );
	vdp_dlatch_inv g4586 (.nQ(w4675), .D(w4752), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4587 (.nZ(w4676), .A(S[6]) );
	vdp_aon22 g4588 (.Z(w4753), .B2(w4665), .B1(w4669), .A1(w4668), .A2(w4667) );
	vdp_dlatch_inv g4589 (.nQ(w4667), .D(w6661), .nC(nHCLK1), .C(HCLK1) );
	vdp_not g4590 (.nZ(w4669), .A(S[7]) );
	vdp_aon22 g4591 (.Z(w4755), .B2(w4665), .B1(w4910), .A1(w4668), .A2(1'b1) );
	vdp_dlatch_inv g4592 (.nQ(w4910), .D(w4666), .nC(nHCLK1), .C(HCLK1) );
	vdp_aon22 g4593 (.Z(w4757), .B2(w4665), .B1(1'b1), .A1(w4668), .A2(w4674) );
	vdp_dlatch_inv g4594 (.nQ(w4674), .D(w4673), .nC(nHCLK1), .C(HCLK1) );
	vdp_sr_bit g4595 (.Q(w4644), .D(w6578), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4596 (.Q(w4656), .D(w30), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4597 (.Q(w4677), .D(w4656), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4598 (.Q(w4661), .D(w5), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4599 (.Q(w4671), .D(w4661), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4600 (.Q(w4684), .D(w6577), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_not g4601 (.nZ(w4679), .A(w4678) );
	vdp_not g4602 (.nZ(w4672), .A(M5) );
	vdp_not g4603 (.nZ(w6578), .A(w4670) );
	vdp_not g4604 (.nZ(w4660), .A(w4671) );
	vdp_not g4605 (.nZ(w6577), .A(w4663) );
	vdp_not g4606 (.nZ(w4658), .A(w4643) );
	vdp_aon22 g4607 (.Z(w4763), .B2(w4759), .B1(w4569), .A1(w4758), .A2(w4568) );
	vdp_aon22 g4608 (.Z(w4762), .B2(w4759), .B1(w4568), .A1(w4758), .A2(w4567) );
	vdp_aon22 g4609 (.Z(w4761), .B2(w4759), .B1(w4567), .A1(w4758), .A2(1'b0) );
	vdp_slatch g4610 (.nQ(w6670), .D(w4889), .nC(w4873), .C(w4878) );
	vdp_aon22 g4611 (.Z(w4889), .B2(w4872), .B1(w4747), .A1(w4877), .A2(w4715) );
	vdp_notif0 g4612 (.A(w6670), .nZ(AD_DATA[0]), .nE(w4883) );
	vdp_slatch g4613 (.nQ(w6669), .D(w4888), .nC(w4873), .C(w4878) );
	vdp_aon22 g4614 (.Z(w4888), .B2(w4872), .B1(w4750), .A1(w4877), .A2(w4714) );
	vdp_notif0 g4615 (.A(w6669), .nZ(AD_DATA[1]), .nE(w4883) );
	vdp_slatch g4616 (.nQ(w6668), .D(w4887), .nC(w4873), .C(w4878) );
	vdp_aon22 g4617 (.Z(w4887), .B2(w4872), .B1(w4743), .A1(w4877), .A2(w4713) );
	vdp_notif0 g4618 (.A(w6668), .nZ(AD_DATA[2]), .nE(w4883) );
	vdp_slatch g4619 (.nQ(w6667), .D(w6603), .nC(w4873), .C(w4878) );
	vdp_aon22 g4620 (.Z(w6603), .B2(w4872), .B1(w4744), .A1(w4877), .A2(w4712) );
	vdp_notif0 g4621 (.A(w6667), .nZ(AD_DATA[3]), .nE(w4883) );
	vdp_slatch g4622 (.nQ(w6666), .D(w6602), .nC(w4873), .C(w4878) );
	vdp_aon22 g4623 (.Z(w6602), .B2(w4872), .B1(w4726), .A1(w4877), .A2(w4688) );
	vdp_notif0 g4624 (.A(w6666), .nZ(AD_DATA[4]), .nE(w4883) );
	vdp_slatch g4625 (.nQ(w6665), .D(w6601), .nC(w4873), .C(w4878) );
	vdp_aon22 g4626 (.Z(w6601), .B2(w4872), .B1(w4718), .A1(w4877), .A2(w4687) );
	vdp_notif0 g4627 (.A(w6665), .nZ(AD_DATA[5]), .nE(w4883) );
	vdp_slatch g4628 (.nQ(w6664), .D(w4886), .nC(w4873), .C(w4878) );
	vdp_aon22 g4629 (.Z(w4886), .B2(w4872), .B1(w4719), .A1(w4877), .A2(w4682) );
	vdp_notif0 g4630 (.A(w6664), .nZ(AD_DATA[6]), .nE(w4883) );
	vdp_slatch g4631 (.nQ(w6663), .D(w4895), .nC(w4873), .C(w4878) );
	vdp_aon22 g4632 (.Z(w4895), .B2(w4872), .B1(w4717), .A1(w4877), .A2(w4856) );
	vdp_notif0 g4633 (.A(w6663), .nZ(AD_DATA[7]), .nE(w4883) );
	vdp_slatch g4634 (.nQ(w4885), .D(w4884), .nC(w4873), .C(w4878) );
	vdp_aon22 g4635 (.Z(w4884), .B2(w4872), .B1(w4716), .A1(w4877), .A2(w4894) );
	vdp_notif0 g4636 (.A(w4885), .nZ(RD_DATA[0]), .nE(w4883) );
	vdp_slatch g4637 (.nQ(w4882), .D(w4881), .nC(w4873), .C(w4878) );
	vdp_aon22 g4638 (.Z(w4881), .B2(w4872), .B1(w4711), .A1(w4877), .A2(w4879) );
	vdp_notif0 g4639 (.A(w4882), .nZ(RD_DATA[1]), .nE(w4883) );
	vdp_slatch g4640 (.nQ(w4880), .D(w4875), .nC(w4873), .C(w4878) );
	vdp_aon22 g4641 (.Z(w4875), .B2(w4872), .B1(1'b0), .A1(w4877), .A2(w4876) );
	vdp_notif0 g4642 (.A(w4880), .nZ(RD_DATA[2]), .nE(w4883) );
	vdp_not g4643 (.nZ(w4883), .A(w4893) );
	vdp_sr_bit g4644 (.Q(w4562), .D(w6674), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4645 (.Q(w4563), .D(w4852), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4646 (.Q(w4848), .D(w4846), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_dlatch_inv g4647 (.nQ(w4847), .D(w4749), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4648 (.nQ(w4846), .D(w4787), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g4649 (.nQ(w4793), .D(w4789), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4650 (.nQ(w6600), .D(w4790), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4651 (.nQ(w4797), .D(w4791), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4652 (.nQ(w4795), .D(w4792), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4653 (.nQ(w4801), .D(w4796), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4654 (.nQ(w4799), .D(w4798), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4655 (.nQ(w4803), .D(w4802), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4656 (.nQ(w4812), .D(w4800), .nC(nHCLK2), .C(HCLK2) );
	vdp_aon22 g4657 (.Z(w4802), .B2(w4764), .B1(w4777), .A1(w4775), .A2(w4788) );
	vdp_aon22 g4658 (.Z(w4796), .B2(w4764), .B1(w4779), .A1(w4778), .A2(w4788) );
	vdp_aon22 g4659 (.Z(w4791), .B2(w4764), .B1(w4781), .A1(w4780), .A2(w4788) );
	vdp_aon22 g4660 (.Z(w4789), .B2(w4764), .B1(w4784), .A1(w4783), .A2(w4788) );
	vdp_not g4661 (.nZ(w4786), .A(w4749) );
	vdp_not g4662 (.nZ(w4565), .A(w6600) );
	vdp_not g4663 (.nZ(w4566), .A(w4795) );
	vdp_not g4664 (.nZ(w4575), .A(w4799) );
	vdp_not g4665 (.nZ(w4569), .A(w4812) );
	vdp_not g4666 (.nZ(w4808), .A(w4804) );
	vdp_not g4667 (.nZ(w4568), .A(w4806) );
	vdp_dlatch_inv g4668 (.nQ(w4807), .D(w4804), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4669 (.nQ(w4806), .D(w4805), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g4670 (.nZ(w4567), .A(w4815) );
	vdp_dlatch_inv g4671 (.nQ(w4835), .D(w4770), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4672 (.nQ(w4815), .D(w4811), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g4673 (.nZ(w4816), .A(w4836) );
	vdp_dlatch_inv g4674 (.nQ(w4813), .D(w4836), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4675 (.nQ(w4825), .D(w4814), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g4676 (.nZ(w4810), .A(w4821) );
	vdp_dlatch_inv g4677 (.nQ(w4817), .D(w4821), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4678 (.nQ(w4826), .D(w4818), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4679 (.nQ(w4819), .D(w4809), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4680 (.nQ(w4823), .D(w4820), .nC(nHCLK2), .C(HCLK2) );
	vdp_dlatch_inv g4681 (.nQ(w4832), .D(w4822), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g4682 (.nQ(w4834), .D(w4833), .nC(nHCLK2), .C(HCLK2) );
	vdp_sr_bit g4683 (.Q(w4561), .D(w6662), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4684 (.Z(w4822), .B2(w4764), .B1(1'b0), .A1(w4756), .A2(w4788) );
	vdp_aon22 g4685 (.Z(w4809), .B2(w4764), .B1(1'b0), .A1(w4766), .A2(w4788) );
	vdp_aon22 g4686 (.Z(w6662), .B2(w4860), .B1(M5), .A1(w132), .A2(w4906) );
	vdp_not g4687 (.nZ(w4851), .A(w1) );
	vdp_not g4688 (.nZ(w4909), .A(w4863) );
	vdp_not g4689 (.nZ(w4852), .A(w4862) );
	vdp_not g4690 (.nZ(w4907), .A(w4864) );
	vdp_not g4691 (.nZ(w4860), .A(w4861) );
	vdp_not g4692 (.nZ(w4906), .A(M5) );
	vdp_not g4693 (.nZ(w4555), .A(w4858) );
	vdp_not g4694 (.nZ(w4853), .A(w4561) );
	vdp_not g4695 (.nZ(w6671), .A(w4562) );
	vdp_not g4696 (.nZ(w4908), .A(M5) );
	vdp_not g4697 (.nZ(w4824), .A(w1) );
	vdp_not g4698 (.nZ(w4828), .A(w4761) );
	vdp_bufif0 g4699 (.A(1'b0), .Z(VRAMA[0]), .nE(w4658) );
	vdp_bufif0 g4700 (.A(w4646), .Z(VRAMA[1]), .nE(w4658) );
	vdp_bufif0 g4701 (.A(w4650), .Z(VRAMA[2]), .nE(w4658) );
	vdp_bufif0 g4702 (.A(w4653), .Z(VRAMA[3]), .nE(w4658) );
	vdp_bufif0 g4703 (.A(w4649), .Z(VRAMA[4]), .nE(w4658) );
	vdp_bufif0 g4704 (.A(w4647), .Z(VRAMA[5]), .nE(w4658) );
	vdp_bufif0 g4705 (.A(1'b0), .Z(VRAMA[6]), .nE(w4658) );
	vdp_bufif0 g4706 (.A(1'b0), .Z(VRAMA[7]), .nE(w4658) );
	vdp_aon22 g4707 (.Z(w4821), .B2(w4764), .B1(w6658), .A1(w4767), .A2(w4788) );
	vdp_aon22 g4708 (.Z(w4836), .B2(w4764), .B1(w4769), .A1(w4768), .A2(w4788) );
	vdp_aon22 g4709 (.Z(w4770), .B2(w4764), .B1(w4772), .A1(w4771), .A2(w4788) );
	vdp_comp_str g4710 (.A(w4785), .nZ(w4723), .Z(w4722) );
	vdp_and g4711 (.Z(w4748), .B(w4708), .A(w4704) );
	vdp_comp_we g4712 (.A(w4748), .nZ(w4788), .Z(w4764) );
	vdp_comp_str g4713 (.A(w4782), .nZ(w4738), .Z(w4737) );
	vdp_not g4714 (.nZ(w4704), .A(M5) );
	vdp_comp_str g4715 (.A(w4855), .nZ(w4865), .Z(w4857) );
	vdp_comp_str g4716 (.A(w4891), .nZ(w4873), .Z(w4878) );
	vdp_comp_we g4717 (.A(M5), .nZ(w4665), .Z(w4668) );
	vdp_comp_we g4718 (.A(w4700), .nZ(w4692), .Z(w4641) );
	vdp_comp_we g4719 (.A(w4679), .nZ(w4648), .Z(w4683) );
	vdp_comp_we g4720 (.A(M5), .nZ(w4655), .Z(w4651) );
	vdp_comp_we g4721 (.A(w1), .nZ(w4759), .Z(w4758) );
	vdp_comp_we g4722 (.nZ(w4872), .A(w4892), .Z(w4877) );
	vdp_and g4723 (.Z(w4785), .B(w4846), .A(DCLK2) );
	vdp_and g4724 (.Z(w4782), .B(w4848), .A(DCLK2) );
	vdp_and g4725 (.Z(w4845), .B(M5), .A(w4851) );
	vdp_and g4726 (.Z(w6674), .B(w4907), .A(M5) );
	vdp_and g4727 (.Z(w6673), .B(w4853), .A(w4562) );
	vdp_and g4728 (.Z(w4891), .B(w4890), .A(HCLK1) );
	vdp_or g4729 (.Z(w4827), .B(w4824), .A(w4834) );
	vdp_or g4730 (.Z(w6675), .B(w4908), .A(w4823) );
	vdp_and g4731 (.Z(w4643), .B(w4672), .A(w4656) );
	vdp_and g4732 (.Z(w4701), .B(w4637), .A(w4699) );
	vdp_and g4733 (.Z(w6401), .B(w4699), .A(w4638) );
	vdp_and g4734 (.Z(w6402), .B(w4636), .A(w4638) );
	vdp_and g4735 (.Z(w6403), .B(w4637), .A(w4636) );
	vdp_and g4736 (.Z(w6377), .B(H40), .A(VRAMA[9]) );
	vdp_or g4737 (.Z(w4710), .B(w4639), .A(w4708) );
	vdp_or g4738 (.Z(w4709), .B(w4639), .A(w4705) );
	vdp_not g4739 (.nZ(w4636), .A(w4699) );
	vdp_oai21 g4740 (.Z(w4663), .B(w30), .A1(w31), .A2(w5) );
	vdp_oai21 g4741 (.Z(w4858), .B(w4554), .A1(w4776), .A2(w4859) );
	vdp_aoi22 g4742 (.Z(w4749), .B2(w4704), .B1(w4705), .A1(M5), .A2(w4746) );
	vdp_or3 g4743 (.Z(w4746), .B(w6598), .A(w4706), .C(w4707) );
	vdp_and3 g4744 (.Z(w4855), .B(DCLK1), .A(HCLK2), .C(w4847) );
	vdp_oai21 g4745 (.Z(w4678), .B(M5), .A1(w4656), .A2(w4677) );
	vdp_2a3oi g4746 (.Z(w4670), .B(w4661), .A1(w4660), .A2(w4), .C(SYSRES) );
	vdp_or8 g4747 (.Z(w4859), .B(w4871), .A(M5), .C(w6605), .D(w4870), .F(w4868), .E(w4869), .G(w4867), .H(w4866) );
	vdp_and9 g4748 (.Z(w4521), .B(w4829), .A(w4831), .C(w4830), .D(w4828), .F(w4826), .E(w4827), .G(w4825), .H(w4556), .I(w6675) );
	vdp_nor12 g4749 (.Z(w4776), .B(w4770), .A(1'b0), .C(w4810), .D(M5), .F(w4822), .E(w4809), .G(w4816), .H(w4808), .J(w4791), .I(w4796), .K(w4789), .L(w4802) );
	vdp_or4 g4750 (.Z(w4700), .B(w4638), .A(w4637), .C(w4698), .D(w4640) );
	vdp_nand g4751 (.Z(w4787), .B(w4786), .A(HCLK1) );
	vdp_nand g4752 (.Z(w4831), .B(w4763), .A(w6672) );
	vdp_nand g4753 (.Z(w4830), .B(w4762), .A(w6671) );
	vdp_nor g4754 (.Z(w6672), .B(w4561), .A(w4562) );
	vdp_nand3 g4755 (.Z(w4829), .B(w4762), .A(w6673), .C(w4763) );
	vdp_sr_bit g4756 (.Q(w4564), .D(w4909), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4757 (.Q(w4917), .D(w4918), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4758 (.Q(w4584), .D(w6579), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4759 (.Q(w4916), .D(w6563), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4760 (.Q(w6563), .D(w6564), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4761 (.Q(w6564), .D(w4915), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4762 (.Z(w4921), .B2(w4916), .B1(w5282), .A1(DB[4]), .A2(w5283) );
	vdp_noif0 g4763 (.A(HPOS[1]), .nZ(VRAMA[1]), .nE(w5139) );
	vdp_aon22 g4764 (.Z(w6579), .B2(w4914), .B1(w4917), .A1(M5), .A2(w4918) );
	vdp_not g4765 (.nZ(w4914), .A(M5) );
	vdp_lfsr_bit g4766 (.Q(w4922), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6596), .A1(w4921), .A2(w6595) );
	vdp_lfsr_bit g4767 (.Q(w4925), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5284), .A1(w4922), .A2(w6594) );
	vdp_lfsr_bit g4768 (.Q(w4927), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5285), .A1(w4925), .A2(w6593) );
	vdp_lfsr_bit g4769 (.Q(w4928), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5286), .A1(w4927), .A2(w6592) );
	vdp_lfsr_bit g4770 (.Q(w4932), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5287), .A1(w4928), .A2(w6591) );
	vdp_lfsr_bit g4771 (.Q(w4930), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5288), .A1(w4932), .A2(w6590) );
	vdp_lfsr_bit g4772 (.Q(w4934), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5289), .A1(w4930), .A2(w6589) );
	vdp_lfsr_bit g4773 (.Q(w4913), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5290), .A1(w4934), .A2(w6588) );
	vdp_lfsr_bit g4774 (.Q(w4938), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5119), .A1(w4913), .A2(w6587) );
	vdp_lfsr_bit g4775 (.Q(w4940), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5293), .A1(w4938), .A2(w5294) );
	vdp_lfsr_bit g4776 (.Q(w4944), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5167), .A1(w4940), .A2(w5168) );
	vdp_lfsr_bit g4777 (.Q(w4941), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5164), .A1(w4944), .A2(w5165) );
	vdp_lfsr_bit g4778 (.Q(w4943), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5162), .A1(w4941), .A2(w5163) );
	vdp_lfsr_bit g4779 (.Q(w4947), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6586), .A1(w4943), .A2(w5161) );
	vdp_lfsr_bit g4780 (.Q(w4948), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5158), .A1(w4947), .A2(w5159) );
	vdp_lfsr_bit g4781 (.Q(w4952), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6584), .A1(w4948), .A2(w6585) );
	vdp_lfsr_bit g4782 (.Q(w4951), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6583), .A1(w4952), .A2(w6582) );
	vdp_lfsr_bit g4783 (.Q(w4956), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5155), .A1(w4951), .A2(w5156) );
	vdp_lfsr_bit g4784 (.Q(w4958), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5154), .A1(w4956), .A2(w5153) );
	vdp_lfsr_bit g4785 (.Q(w4912), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5151), .A1(w4958), .A2(w5152) );
	vdp_bufif0 g4786 (.A(w4913), .Z(VRAMA[1]), .nE(w6581) );
	vdp_bufif0 g4787 (.A(1'b0), .Z(VRAMA[1]), .nE(w5175) );
	vdp_noif0 g4788 (.A(w4912), .nZ(DB[4]), .nE(w5295) );
	vdp_sr_bit g4789 (.Q(w4965), .D(w6566), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4790 (.Q(w6566), .D(w6565), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4791 (.Q(w6565), .D(w6384), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4792 (.Z(w4920), .B2(w4965), .B1(w5282), .A1(DB[5]), .A2(w5283) );
	vdp_noif0 g4793 (.A(w4974), .nZ(VRAMA[2]), .nE(w5139) );
	vdp_lfsr_bit g4794 (.Q(w4923), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6596), .A1(w4920), .A2(w6595) );
	vdp_lfsr_bit g4795 (.Q(w4924), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5284), .A1(w4923), .A2(w6594) );
	vdp_lfsr_bit g4796 (.Q(w4926), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5285), .A1(w4924), .A2(w6593) );
	vdp_lfsr_bit g4797 (.Q(w4929), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5286), .A1(w4926), .A2(w6592) );
	vdp_lfsr_bit g4798 (.Q(w4933), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5287), .A1(w4929), .A2(w6591) );
	vdp_lfsr_bit g4799 (.Q(w4931), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5288), .A1(w4933), .A2(w6590) );
	vdp_lfsr_bit g4800 (.Q(w4935), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5289), .A1(w4931), .A2(w6589) );
	vdp_lfsr_bit g4801 (.Q(w4936), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5290), .A1(w4935), .A2(w6588) );
	vdp_lfsr_bit g4802 (.Q(w4939), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5119), .A1(w4936), .A2(w6587) );
	vdp_lfsr_bit g4803 (.Q(w4937), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5293), .A1(w4939), .A2(w5294) );
	vdp_lfsr_bit g4804 (.Q(w4945), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5167), .A1(w4937), .A2(w5168) );
	vdp_lfsr_bit g4805 (.Q(w4942), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5164), .A1(w4945), .A2(w5165) );
	vdp_lfsr_bit g4806 (.Q(w4946), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5162), .A1(w4942), .A2(w5163) );
	vdp_lfsr_bit g4807 (.Q(w4950), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6586), .A1(w4946), .A2(w5161) );
	vdp_lfsr_bit g4808 (.Q(w4949), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5158), .A1(w4950), .A2(w5159) );
	vdp_lfsr_bit g4809 (.Q(w4953), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6584), .A1(w4949), .A2(w6585) );
	vdp_lfsr_bit g4810 (.Q(w4954), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6583), .A1(w4953), .A2(w6582) );
	vdp_lfsr_bit g4811 (.Q(w4955), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5155), .A1(w4954), .A2(w5156) );
	vdp_lfsr_bit g4812 (.Q(w4959), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5154), .A1(w4955), .A2(w5153) );
	vdp_lfsr_bit g4813 (.Q(w4963), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5151), .A1(w4959), .A2(w5152) );
	vdp_bufif0 g4814 (.A(w4936), .Z(VRAMA[2]), .nE(w6581) );
	vdp_bufif0 g4815 (.A(1'b1), .Z(VRAMA[2]), .nE(w5175) );
	vdp_noif0 g4816 (.A(w4963), .nZ(DB[5]), .nE(w5295) );
	vdp_aon22 g4817 (.Z(w4962), .B2(w4952), .B1(w5148), .A1(w5147), .A2(w4912) );
	vdp_dlatch_inv g4818 (.nQ(w4975), .D(w4968), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g4819 (.nQ(w4970), .D(w4919), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g4820 (.Z(w4969), .B(w4970), .A(DCLK2) );
	vdp_nand g4821 (.Z(w4968), .B(HCLK1), .A(w4584) );
	vdp_nand g4822 (.Z(w4919), .B(HCLK1), .A(w4918) );
	vdp_sr_bit g4823 (.Q(w4967), .D(w6568), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4824 (.Q(w6568), .D(w6567), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4825 (.Q(w6567), .D(w4972), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4826 (.Z(w4983), .B2(w4967), .B1(w5282), .A1(w4966), .A2(w5283) );
	vdp_noif0 g4827 (.A(w4981), .nZ(VRAMA[3]), .nE(w5139) );
	vdp_lfsr_bit g4828 (.Q(w4985), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6596), .A1(w4983), .A2(w6595) );
	vdp_lfsr_bit g4829 (.Q(w4986), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5284), .A1(w4985), .A2(w6594) );
	vdp_lfsr_bit g4830 (.Q(w4989), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5285), .A1(w4986), .A2(w6593) );
	vdp_lfsr_bit g4831 (.Q(w4990), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5286), .A1(w4989), .A2(w6592) );
	vdp_lfsr_bit g4832 (.Q(w4995), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5287), .A1(w4990), .A2(w6591) );
	vdp_lfsr_bit g4833 (.Q(w4994), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5288), .A1(w4995), .A2(w6590) );
	vdp_lfsr_bit g4834 (.Q(w4997), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5289), .A1(w4994), .A2(w6589) );
	vdp_lfsr_bit g4835 (.Q(w4999), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5290), .A1(w4997), .A2(w6588) );
	vdp_lfsr_bit g4836 (.Q(w5001), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5119), .A1(w4999), .A2(w6587) );
	vdp_lfsr_bit g4837 (.Q(w5003), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5293), .A1(w5001), .A2(w5294) );
	vdp_lfsr_bit g4838 (.Q(w5005), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5167), .A1(w5003), .A2(w5168) );
	vdp_lfsr_bit g4839 (.Q(w5007), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5164), .A1(w5005), .A2(w5165) );
	vdp_lfsr_bit g4840 (.Q(w5009), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5162), .A1(w5007), .A2(w5163) );
	vdp_lfsr_bit g4841 (.Q(w5012), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6586), .A1(w5009), .A2(w5161) );
	vdp_lfsr_bit g4842 (.Q(w5013), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5158), .A1(w5012), .A2(w5159) );
	vdp_lfsr_bit g4843 (.Q(w5014), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6584), .A1(w5013), .A2(w6585) );
	vdp_lfsr_bit g4844 (.Q(w5019), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6583), .A1(w5014), .A2(w6582) );
	vdp_lfsr_bit g4845 (.Q(w5018), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5155), .A1(w5019), .A2(w5156) );
	vdp_lfsr_bit g4846 (.Q(w5021), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5154), .A1(w5018), .A2(w5153) );
	vdp_lfsr_bit g4847 (.Q(w4964), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5151), .A1(w5021), .A2(w5152) );
	vdp_bufif0 g4848 (.A(w4999), .Z(VRAMA[3]), .nE(w6581) );
	vdp_bufif0 g4849 (.A(w4962), .Z(VRAMA[3]), .nE(w5175) );
	vdp_noif0 g4850 (.A(w4964), .nZ(w4966), .nE(w5295) );
	vdp_aon22 g4851 (.Z(w5022), .B2(w4953), .B1(w5148), .A1(w5147), .A2(w4963) );
	vdp_sr_bit g4852 (.Q(w4977), .D(w4975), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g4853 (.Q(w4971), .D(w4970), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_and g4854 (.Z(w4973), .B(w4975), .A(DCLK2) );
	vdp_and g4855 (.Z(w4979), .B(DCLK2), .A(w4977) );
	vdp_and g4856 (.Z(w4976), .B(w4971), .A(DCLK2) );
	vdp_sr_bit g4857 (.Q(w5035), .D(w6569), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4858 (.Q(w6569), .D(w6570), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4859 (.Q(w6570), .D(w4978), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4860 (.Z(w4982), .B2(w5035), .B1(w5282), .A1(DB[7]), .A2(w5283) );
	vdp_noif0 g4861 (.A(w5033), .nZ(VRAMA[4]), .nE(w5139) );
	vdp_lfsr_bit g4862 (.Q(w4984), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6596), .A1(w4982), .A2(w6595) );
	vdp_lfsr_bit g4863 (.Q(w4987), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5284), .A1(w4984), .A2(w6594) );
	vdp_lfsr_bit g4864 (.Q(w4988), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5285), .A1(w4987), .A2(w6593) );
	vdp_lfsr_bit g4865 (.Q(w4991), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5286), .A1(w4988), .A2(w6592) );
	vdp_lfsr_bit g4866 (.Q(w4992), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5287), .A1(w4991), .A2(w6591) );
	vdp_lfsr_bit g4867 (.Q(w4993), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5288), .A1(w4992), .A2(w6590) );
	vdp_lfsr_bit g4868 (.Q(w4996), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5289), .A1(w4993), .A2(w6589) );
	vdp_lfsr_bit g4869 (.Q(w4998), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5290), .A1(w4996), .A2(w6588) );
	vdp_lfsr_bit g4870 (.Q(w5000), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5119), .A1(w4998), .A2(w6587) );
	vdp_lfsr_bit g4871 (.Q(w5002), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5293), .A1(w5000), .A2(w5294) );
	vdp_lfsr_bit g4872 (.Q(w5004), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5167), .A1(w5002), .A2(w5168) );
	vdp_lfsr_bit g4873 (.Q(w5006), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5164), .A1(w5004), .A2(w5165) );
	vdp_lfsr_bit g4874 (.Q(w5008), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5162), .A1(w5006), .A2(w5163) );
	vdp_lfsr_bit g4875 (.Q(w5011), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6586), .A1(w5008), .A2(w5161) );
	vdp_lfsr_bit g4876 (.Q(w5010), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5158), .A1(w5011), .A2(w5159) );
	vdp_lfsr_bit g4877 (.Q(w5015), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6584), .A1(w5010), .A2(w6585) );
	vdp_lfsr_bit g4878 (.Q(w5016), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6583), .A1(w5015), .A2(w6582) );
	vdp_lfsr_bit g4879 (.Q(w5017), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5155), .A1(w5016), .A2(w5156) );
	vdp_lfsr_bit g4880 (.Q(w5020), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5154), .A1(w5017), .A2(w5153) );
	vdp_lfsr_bit g4881 (.Q(w5037), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5151), .A1(w5020), .A2(w5152) );
	vdp_bufif0 g4882 (.A(w4998), .Z(VRAMA[4]), .nE(w6581) );
	vdp_bufif0 g4883 (.A(w5022), .Z(VRAMA[4]), .nE(w5175) );
	vdp_noif0 g4884 (.A(w5037), .nZ(DB[7]), .nE(w5295) );
	vdp_aon22 g4885 (.Z(w5038), .B2(w5014), .B1(w5148), .A1(w5147), .A2(w4964) );
	vdp_aon22 g4886 (.Z(w5032), .B2(w5025), .B1(w132), .A1(w4980), .A2(w5031) );
	vdp_not g4887 (.nZ(w4980), .A(w132) );
	vdp_comp_str g4888 (.nZ(w5026), .A(w4976), .Z(w5027) );
	vdp_comp_str g4889 (.nZ(w5030), .A(w4979), .Z(w5029) );
	vdp_sr_bit g4890 (.Q(w5034), .D(w6572), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4891 (.Q(w6572), .D(w6571), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4892 (.Q(w6571), .D(w5028), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4893 (.Z(w5079), .B2(w5034), .B1(w5282), .A1(DB[8]), .A2(w5283) );
	vdp_noif0 g4894 (.A(w5032), .nZ(VRAMA[5]), .nE(w5139) );
	vdp_lfsr_bit g4895 (.Q(w5077), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6596), .A1(w5079), .A2(w6595) );
	vdp_lfsr_bit g4896 (.Q(w5074), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5284), .A1(w5077), .A2(w6594) );
	vdp_lfsr_bit g4897 (.Q(w5073), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5285), .A1(w5074), .A2(w6593) );
	vdp_lfsr_bit g4898 (.Q(w5070), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5286), .A1(w5073), .A2(w6592) );
	vdp_lfsr_bit g4899 (.Q(w5069), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5287), .A1(w5070), .A2(w6591) );
	vdp_lfsr_bit g4900 (.Q(w5066), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5288), .A1(w5069), .A2(w6590) );
	vdp_lfsr_bit g4901 (.Q(w5065), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5289), .A1(w5066), .A2(w6589) );
	vdp_lfsr_bit g4902 (.Q(w5043), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5290), .A1(w5065), .A2(w6588) );
	vdp_lfsr_bit g4903 (.Q(w5062), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5119), .A1(w5043), .A2(w6587) );
	vdp_lfsr_bit g4904 (.Q(w5036), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5293), .A1(w5062), .A2(w5294) );
	vdp_lfsr_bit g4905 (.Q(w5059), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5167), .A1(w5036), .A2(w5168) );
	vdp_lfsr_bit g4906 (.Q(w5058), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5164), .A1(w5059), .A2(w5165) );
	vdp_lfsr_bit g4907 (.Q(w5055), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5162), .A1(w5058), .A2(w5163) );
	vdp_lfsr_bit g4908 (.Q(w5053), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6586), .A1(w5055), .A2(w5161) );
	vdp_lfsr_bit g4909 (.Q(w5052), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5158), .A1(w5053), .A2(w5159) );
	vdp_lfsr_bit g4910 (.Q(w5041), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6584), .A1(w5052), .A2(w6585) );
	vdp_lfsr_bit g4911 (.Q(w5048), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6583), .A1(w5041), .A2(w6582) );
	vdp_lfsr_bit g4912 (.Q(w5046), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5155), .A1(w5048), .A2(w5156) );
	vdp_lfsr_bit g4913 (.Q(w5044), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5154), .A1(w5046), .A2(w5153) );
	vdp_lfsr_bit g4914 (.Q(w5061), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5151), .A1(w5044), .A2(w5152) );
	vdp_bufif0 g4915 (.A(w5043), .Z(VRAMA[5]), .nE(w6581) );
	vdp_bufif0 g4916 (.A(w5038), .Z(VRAMA[5]), .nE(w5175) );
	vdp_noif0 g4917 (.A(w5061), .nZ(DB[8]), .nE(w5295) );
	vdp_aon22 g4918 (.Z(w5040), .B2(w5015), .B1(w5148), .A1(w5147), .A2(w5037) );
	vdp_slatch g4919 (.D(S[0]), .nC(w5030), .C(w5029), .Q(w5084) );
	vdp_slatch g4920 (.D(S[0]), .nC(w5026), .C(w5027), .Q(w5024) );
	vdp_aoi22 g4921 (.Z(w5031), .B2(w5083), .B1(w5084), .A1(w5082), .A2(w5024) );
	vdp_sr_bit g4922 (.Q(w5092), .D(w6574), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4923 (.Q(w6574), .D(w6573), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4924 (.Q(w6573), .D(w5080), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4925 (.Z(w5078), .B2(w5092), .B1(w5282), .A1(DB[9]), .A2(w5283) );
	vdp_noif0 g4926 (.A(w5081), .nZ(VRAMA[6]), .nE(w5139) );
	vdp_lfsr_bit g4927 (.Q(w5076), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w6596), .A1(w5078), .A2(w6595) );
	vdp_lfsr_bit g4928 (.Q(w5075), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w5284), .A1(w5076), .A2(w6594) );
	vdp_lfsr_bit g4929 (.Q(w5072), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w5285), .A1(w5075), .A2(w6593) );
	vdp_lfsr_bit g4930 (.Q(w5071), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w5286), .A1(w5072), .A2(w6592) );
	vdp_lfsr_bit g4931 (.Q(w5068), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w5287), .A1(w5071), .A2(w6591) );
	vdp_lfsr_bit g4932 (.Q(w5067), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w5288), .A1(w5068), .A2(w6590) );
	vdp_lfsr_bit g4933 (.Q(w5064), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w5289), .A1(w5067), .A2(w6589) );
	vdp_lfsr_bit g4934 (.Q(w5042), .C2(nHCLK2), .C1(nHCLK1), .nC2(HCLK2), .nC1(HCLK1), .B(w5290), .A1(w5064), .A2(w6588) );
	vdp_lfsr_bit g4935 (.Q(w5063), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5119), .A1(w5042), .A2(w6587) );
	vdp_lfsr_bit g4936 (.Q(w5090), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5293), .A1(w5063), .A2(w5294) );
	vdp_lfsr_bit g4937 (.Q(w5060), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5167), .A1(w5090), .A2(w5168) );
	vdp_lfsr_bit g4938 (.Q(w5057), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5164), .A1(w5060), .A2(w5165) );
	vdp_lfsr_bit g4939 (.Q(w5056), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5162), .A1(w5057), .A2(w5163) );
	vdp_lfsr_bit g4940 (.Q(w5054), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6586), .A1(w5056), .A2(w5161) );
	vdp_lfsr_bit g4941 (.Q(w5051), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5158), .A1(w5054), .A2(w5159) );
	vdp_lfsr_bit g4942 (.Q(w5050), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6584), .A1(w5051), .A2(w6585) );
	vdp_lfsr_bit g4943 (.Q(w5049), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6583), .A1(w5050), .A2(w6582) );
	vdp_lfsr_bit g4944 (.Q(w5047), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5155), .A1(w5049), .A2(w5156) );
	vdp_lfsr_bit g4945 (.Q(w5045), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5154), .A1(w5047), .A2(w5153) );
	vdp_lfsr_bit g4946 (.Q(w5087), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5151), .A1(w5045), .A2(w5152) );
	vdp_bufif0 g4947 (.A(w5042), .Z(VRAMA[6]), .nE(w6581) );
	vdp_bufif0 g4948 (.A(w5040), .Z(VRAMA[6]), .nE(w5175) );
	vdp_noif0 g4949 (.A(w5087), .nZ(DB[9]), .nE(w5295) );
	vdp_aon22 g4950 (.Z(w5089), .B2(w5041), .B1(w5148), .A1(w5147), .A2(w5061) );
	vdp_aoi22 g4951 (.Z(w5081), .B2(w5083), .B1(w5094), .A1(w5082), .A2(w5085) );
	vdp_slatch g4952 (.D(S[1]), .nC(w5030), .C(w5029), .Q(w5094) );
	vdp_slatch g4953 (.D(S[1]), .nC(w5026), .C(w5027), .Q(w5085) );
	vdp_sr_bit g4954 (.Q(w5091), .D(w6576), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4955 (.Q(w6576), .D(w6575), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4956 (.Q(w6575), .D(w5095), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4957 (.Z(w5138), .B2(w5091), .B1(w5282), .A1(DB[10]), .A2(w5283) );
	vdp_noif0 g4958 (.A(w5141), .nZ(VRAMA[7]), .nE(w5142) );
	vdp_lfsr_bit g4959 (.Q(w5137), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6596), .A1(w5138), .A2(w6595) );
	vdp_lfsr_bit g4960 (.Q(w5132), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5284), .A1(w5137), .A2(w6594) );
	vdp_lfsr_bit g4961 (.Q(w5133), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5285), .A1(w5132), .A2(w6593) );
	vdp_lfsr_bit g4962 (.Q(w5127), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5286), .A1(w5133), .A2(w6592) );
	vdp_lfsr_bit g4963 (.Q(w5128), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5287), .A1(w5127), .A2(w6591) );
	vdp_lfsr_bit g4964 (.Q(w5125), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5288), .A1(w5128), .A2(w6590) );
	vdp_lfsr_bit g4965 (.Q(w5123), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5289), .A1(w5125), .A2(w6589) );
	vdp_lfsr_bit g4966 (.Q(w5088), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5290), .A1(w5123), .A2(w6588) );
	vdp_lfsr_bit g4967 (.Q(w5120), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5119), .A1(w5088), .A2(w6587) );
	vdp_lfsr_bit g4968 (.Q(w5115), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5293), .A1(w5120), .A2(w5294) );
	vdp_lfsr_bit g4969 (.Q(w5117), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5167), .A1(w5115), .A2(w5168) );
	vdp_lfsr_bit g4970 (.Q(w5114), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5164), .A1(w5117), .A2(w5165) );
	vdp_lfsr_bit g4971 (.Q(w5113), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5162), .A1(w5114), .A2(w5163) );
	vdp_lfsr_bit g4972 (.Q(w5110), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6586), .A1(w5113), .A2(w5161) );
	vdp_lfsr_bit g4973 (.Q(w5108), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5158), .A1(w5110), .A2(w5159) );
	vdp_lfsr_bit g4974 (.Q(w5106), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6584), .A1(w5108), .A2(w6585) );
	vdp_lfsr_bit g4975 (.Q(w5104), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6583), .A1(w5106), .A2(w6582) );
	vdp_lfsr_bit g4976 (.Q(w5102), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5155), .A1(w5104), .A2(w5156) );
	vdp_lfsr_bit g4977 (.Q(w5100), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5154), .A1(w5102), .A2(w5153) );
	vdp_lfsr_bit g4978 (.Q(w5098), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5151), .A1(w5100), .A2(w5152) );
	vdp_bufif0 g4979 (.A(w5088), .Z(VRAMA[7]), .nE(w6581) );
	vdp_bufif0 g4980 (.A(w5089), .Z(VRAMA[7]), .nE(w5175) );
	vdp_noif0 g4981 (.A(w5098), .nZ(DB[10]), .nE(w5295) );
	vdp_aon22 g4982 (.Z(w5097), .B2(w5050), .B1(w5148), .A1(w5147), .A2(w5087) );
	vdp_aoi22 g4983 (.Z(w5141), .B2(w5083), .B1(w5143), .A1(w5082), .A2(w5093) );
	vdp_slatch g4984 (.D(S[2]), .nC(w5030), .C(w5029), .Q(w5143) );
	vdp_slatch g4985 (.D(S[2]), .nC(w5026), .C(w5027), .Q(w5093) );
	vdp_sr_bit g4986 (.Q(w5170), .D(w29), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g4987 (.Q(w5169), .D(w22), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g4988 (.Z(w5135), .B2(w4559), .B1(w5282), .A1(DB[11]), .A2(w5283) );
	vdp_noif0 g4989 (.A(w5140), .nZ(VRAMA[8]), .nE(w5142) );
	vdp_lfsr_bit g4990 (.Q(w5136), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6596), .A1(w5135), .A2(w6595) );
	vdp_lfsr_bit g4991 (.Q(w5131), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5284), .A1(w5136), .A2(w6594) );
	vdp_lfsr_bit g4992 (.Q(w5134), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5285), .A1(w5131), .A2(w6593) );
	vdp_lfsr_bit g4993 (.Q(w5130), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5286), .A1(w5134), .A2(w6592) );
	vdp_lfsr_bit g4994 (.Q(w5129), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5287), .A1(w5130), .A2(w6591) );
	vdp_lfsr_bit g4995 (.Q(w5126), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5288), .A1(w5129), .A2(w6590) );
	vdp_lfsr_bit g4996 (.Q(w5124), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5289), .A1(w5126), .A2(w6589) );
	vdp_lfsr_bit g4997 (.Q(w5122), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5290), .A1(w5124), .A2(w6588) );
	vdp_lfsr_bit g4998 (.Q(w5121), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5119), .A1(w5122), .A2(w6587) );
	vdp_lfsr_bit g4999 (.Q(w5118), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5293), .A1(w5121), .A2(w5294) );
	vdp_lfsr_bit g5000 (.Q(w5116), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5167), .A1(w5118), .A2(w5168) );
	vdp_lfsr_bit g5001 (.Q(w5112), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5164), .A1(w5116), .A2(w5165) );
	vdp_lfsr_bit g5002 (.Q(w5111), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5162), .A1(w5112), .A2(w5163) );
	vdp_lfsr_bit g5003 (.Q(w5109), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6586), .A1(w5111), .A2(w5161) );
	vdp_lfsr_bit g5004 (.Q(w5107), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5158), .A1(w5109), .A2(w5159) );
	vdp_lfsr_bit g5005 (.Q(w5105), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6584), .A1(w5107), .A2(w6585) );
	vdp_lfsr_bit g5006 (.Q(w5103), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6583), .A1(w5105), .A2(w6582) );
	vdp_lfsr_bit g5007 (.Q(w5101), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5155), .A1(w5103), .A2(w5156) );
	vdp_lfsr_bit g5008 (.Q(w5099), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5154), .A1(w5101), .A2(w5153) );
	vdp_lfsr_bit g5009 (.Q(w5166), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5151), .A1(w5099), .A2(w5152) );
	vdp_bufif0 g5010 (.A(1'b0), .Z(VRAMA[0]), .nE(w6581) );
	vdp_bufif0 g5011 (.A(w5097), .Z(VRAMA[8]), .nE(w5175) );
	vdp_noif0 g5012 (.A(w5166), .nZ(DB[11]), .nE(w5295) );
	vdp_aon22 g5013 (.Z(w5176), .B2(w5149), .B1(w5148), .A1(w5147), .A2(w5098) );
	vdp_aoi22 g5014 (.Z(w5140), .B2(w5083), .B1(w5144), .A1(w5082), .A2(w5145) );
	vdp_slatch g5015 (.D(S[3]), .nC(w5030), .C(w5029), .Q(w5144) );
	vdp_slatch g5016 (.D(S[3]), .nC(w5026), .C(w5027), .Q(w5145) );
	vdp_bufif0 g5017 (.A(1'b0), .Z(VRAMA[0]), .nE(w5175) );
	vdp_bufif0 g5018 (.A(w5179), .Z(VRAMA[8]), .nE(w5183) );
	vdp_aon22 g5019 (.Z(w5206), .B2(w4569), .B1(w5282), .A1(DB[3]), .A2(w5283) );
	vdp_lfsr_bit g5020 (.Q(w5204), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6596), .A1(w5206), .A2(w6595) );
	vdp_lfsr_bit g5021 (.Q(w5202), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5284), .A1(w5204), .A2(w6594) );
	vdp_lfsr_bit g5022 (.Q(w5200), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5285), .A1(w5202), .A2(w6593) );
	vdp_lfsr_bit g5023 (.Q(w5198), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5286), .A1(w5200), .A2(w6592) );
	vdp_lfsr_bit g5024 (.Q(w5195), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5287), .A1(w5198), .A2(w6591) );
	vdp_lfsr_bit g5025 (.Q(w5194), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5288), .A1(w5195), .A2(w6590) );
	vdp_lfsr_bit g5026 (.Q(w5192), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5289), .A1(w5194), .A2(w6589) );
	vdp_lfsr_bit g5027 (.Q(w5190), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5290), .A1(w5192), .A2(w6588) );
	vdp_lfsr_bit g5028 (.Q(w5174), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5119), .A1(w5190), .A2(w6587) );
	vdp_lfsr_bit g5029 (.Q(w5172), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5293), .A1(w5174), .A2(w5294) );
	vdp_noif0 g5030 (.A(w5172), .nZ(DB[3]), .nE(w5295) );
	vdp_not g5031 (.nZ(w5160), .A(M5) );
	vdp_not g5032 (.nZ(w5171), .A(H40) );
	vdp_noif0 g5033 (.A(1'b1), .nZ(VRAMA[0]), .nE(w5139) );
	vdp_aoi22 g5034 (.Z(w5025), .B2(w5211), .B1(w5174), .A1(w5082), .A2(w5172) );
	vdp_not g5035 (.nZ(w5208), .A(M5) );
	vdp_or g5036 (.Z(w5209), .B(w5170), .A(w5169) );
	vdp_sr_bit g5037 (.Q(w5180), .D(w9), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5038 (.Q(w5186), .D(w30), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_comp_we g5039 (.nZ(w5151), .A(w5178), .Z(w5152) );
	vdp_comp_we g5040 (.nZ(w5154), .A(w5178), .Z(w5153) );
	vdp_comp_we g5041 (.nZ(w5155), .A(w5178), .Z(w5156) );
	vdp_comp_we g5042 (.nZ(w6583), .A(w5178), .Z(w6582) );
	vdp_comp_we g5043 (.nZ(w6584), .A(w5178), .Z(w6585) );
	vdp_comp_we g5044 (.nZ(w5148), .A(H40), .Z(w5147) );
	vdp_comp_we g5045 (.nZ(w5158), .A(w5178), .Z(w5159) );
	vdp_comp_we g5046 (.nZ(w6586), .A(w5178), .Z(w5161) );
	vdp_comp_we g5047 (.nZ(w5162), .A(w5178), .Z(w5163) );
	vdp_comp_we g5048 (.nZ(w5164), .A(w5178), .Z(w5165) );
	vdp_comp_we g5049 (.nZ(w5167), .A(w5178), .Z(w5168) );
	vdp_comp_we g5050 (.nZ(w5083), .A(w5169), .Z(w5082) );
	vdp_not g5051 (.nZ(w5142), .A(w5173) );
	vdp_not g5052 (.nZ(w5139), .A(w5173) );
	vdp_not g5053 (.nZ(w5175), .A(w5182) );
	vdp_not g5054 (.nZ(w6581), .A(w5157) );
	vdp_and g5055 (.Z(w5157), .B(w5180), .A(w5160) );
	vdp_oai21 g5056 (.Z(w5185), .B(w5160), .A1(w5186), .A2(w5180) );
	vdp_aon333 g5057 (.Z(w4520), .B1(M5), .A1(1'b1), .C1(M5), .A2(w5160), .A3(w5122), .B2(w5105), .B3(w5171), .C2(H40), .C3(w5166) );
	vdp_aon22 g5058 (.Z(w5205), .B2(w4575), .B1(w5282), .A1(DB[2]), .A2(w5283) );
	vdp_lfsr_bit g5059 (.Q(w5203), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6596), .A1(w5205), .A2(w6595) );
	vdp_lfsr_bit g5060 (.Q(w5201), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5284), .A1(w5203), .A2(w6594) );
	vdp_lfsr_bit g5061 (.Q(w5199), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5285), .A1(w5201), .A2(w6593) );
	vdp_lfsr_bit g5062 (.Q(w5197), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5286), .A1(w5199), .A2(w6592) );
	vdp_lfsr_bit g5063 (.Q(w5196), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5287), .A1(w5197), .A2(w6591) );
	vdp_lfsr_bit g5064 (.Q(w5193), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5288), .A1(w5196), .A2(w6590) );
	vdp_lfsr_bit g5065 (.Q(w5191), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5289), .A1(w5193), .A2(w6589) );
	vdp_lfsr_bit g5066 (.Q(w5189), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5290), .A1(w5191), .A2(w6588) );
	vdp_lfsr_bit g5067 (.Q(w5188), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5119), .A1(w5189), .A2(w6587) );
	vdp_lfsr_bit g5068 (.Q(w5187), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5293), .A1(w5188), .A2(w5294) );
	vdp_noif0 g5069 (.A(w5187), .nZ(DB[2]), .nE(w5295) );
	vdp_aoi22 g5070 (.Z(w5033), .B2(w5211), .B1(w5188), .A1(w5082), .A2(w5187) );
	vdp_aoi22 g5071 (.Z(w5224), .B2(w5211), .B1(w5225), .A1(w5082), .A2(w4522) );
	vdp_noif0 g5072 (.A(w5224), .nZ(VRAMA[9]), .nE(w5142) );
	vdp_slatch g5074 (.D(S[4]), .nC(w5027), .C(w5026), .Q(w4522) );
	vdp_and g5075 (.Z(w5173), .B(w5208), .A(w5209) );
	vdp_slatch g5076 (.D(REG_BUS[0]), .nC(w5292), .C(w5291), .Q(w5149) );
	vdp_slatch g5077 (.D(REG_BUS[7]), .nC(w5292), .C(w5291), .Q(w5181) );
	vdp_bufif0 g5078 (.A(w5176), .Z(VRAMA[9]), .nE(w5214) );
	vdp_bufif0 g5079 (.A(w5181), .Z(VRAMA[16]), .nE(w5214) );
	vdp_and g5080 (.Z(w5182), .B(w5180), .A(M5) );
	vdp_not g5081 (.nZ(w5214), .A(w5182) );
	vdp_not g5082 (.nZ(w5183), .A(w5184) );
	vdp_not g5083 (.nZ(w5184), .A(w5185) );
	vdp_xor g5084 (.Z(w5213), .B(w5181), .A(VRAMA[16]) );
	vdp_xor g5085 (.Z(w5217), .B(w5219), .A(w5218) );
	vdp_and3 g5086 (.Z(w5210), .B(w5223), .A(w5220), .C(M5) );
	vdp_nor g5087 (.Z(w5219), .B(H40), .A(w5149) );
	vdp_nor g5088 (.Z(w5218), .B(H40), .A(VRAMA[9]) );
	vdp_aon22 g5089 (.Z(w5244), .B2(w4566), .B1(w5282), .A1(DB[1]), .A2(w5283) );
	vdp_lfsr_bit g5090 (.Q(w5243), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w6596), .A1(w5244), .A2(w6595) );
	vdp_lfsr_bit g5091 (.Q(w5242), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5284), .A1(w5243), .A2(w6594) );
	vdp_lfsr_bit g5092 (.Q(w5241), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5285), .A1(w5242), .A2(w6593) );
	vdp_lfsr_bit g5093 (.Q(w5240), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5286), .A1(w5241), .A2(w6592) );
	vdp_lfsr_bit g5094 (.Q(w5239), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5287), .A1(w5240), .A2(w6591) );
	vdp_lfsr_bit g5095 (.Q(w5238), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5288), .A1(w5239), .A2(w6590) );
	vdp_lfsr_bit g5096 (.Q(w5237), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5289), .A1(w5238), .A2(w6589) );
	vdp_lfsr_bit g5097 (.Q(w5236), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5290), .A1(w5237), .A2(w6588) );
	vdp_lfsr_bit g5098 (.Q(w5222), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5119), .A1(w5236), .A2(w6587) );
	vdp_lfsr_bit g5099 (.Q(w5234), .C2(HCLK2), .C1(HCLK1), .nC2(nHCLK2), .nC1(nHCLK1), .B(w5293), .A1(w5222), .A2(w5294) );
	vdp_noif0 g5100 (.A(w5234), .nZ(DB[1]), .nE(w5295) );
	vdp_slatch g5101 (.D(REG_BUS[1]), .nC(w5292), .C(w5291), .Q(w5179) );
	vdp_slatch g5102 (.D(REG_BUS[6]), .nC(w5292), .C(w5291), .Q(w5233) );
	vdp_xor g5103 (.Z(w5216), .B(w5233), .A(VRAMA[15]) );
	vdp_xor g5104 (.Z(w5215), .B(w5179), .A(VRAMA[10]) );
	vdp_aon22 g5105 (.Z(w5253), .B2(w4565), .B1(w5282), .A1(DB[0]), .A2(w5283) );
	vdp_lfsr_bit g5106 (.Q(w5254), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w6596), .A1(w5253), .A2(w6595) );
	vdp_lfsr_bit g5107 (.Q(w5255), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5284), .A1(w5254), .A2(w6594) );
	vdp_lfsr_bit g5108 (.Q(w5256), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5285), .A1(w5255), .A2(w6593) );
	vdp_lfsr_bit g5109 (.Q(w5258), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5286), .A1(w5256), .A2(w6592) );
	vdp_lfsr_bit g5110 (.Q(w5257), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5287), .A1(w5258), .A2(w6591) );
	vdp_lfsr_bit g5111 (.Q(w5260), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5288), .A1(w5257), .A2(w6590) );
	vdp_lfsr_bit g5112 (.Q(w5259), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5289), .A1(w5260), .A2(w6589) );
	vdp_lfsr_bit g5113 (.Q(w5261), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5290), .A1(w5259), .A2(w6588) );
	vdp_lfsr_bit g5114 (.Q(w5235), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5119), .A1(w5261), .A2(w6587) );
	vdp_lfsr_bit g5115 (.Q(w6580), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .B(w5293), .A1(w5235), .A2(w5294) );
	vdp_noif0 g5116 (.A(w6580), .nZ(DB[0]), .nE(w5295) );
	vdp_slatch g5117 (.D(REG_BUS[2]), .nC(w5292), .C(w5291), .Q(w5232) );
	vdp_slatch g5118 (.D(REG_BUS[5]), .nC(w5292), .C(w5291), .Q(w5276) );
	vdp_xor g5119 (.Z(w5229), .B(w5276), .A(VRAMA[14]) );
	vdp_xor g5120 (.Z(w5228), .B(w5232), .A(VRAMA[11]) );
	vdp_slatch g5121 (.D(S[5]), .nC(w5029), .C(w5030), .Q(w5247) );
	vdp_slatch g5122 (.D(S[5]), .nC(w5027), .C(w5026), .Q(w5226) );
	vdp_slatch g5123 (.D(S[6]), .nC(w5029), .C(w5030), .Q(w5248) );
	vdp_slatch g5124 (.D(S[6]), .nC(w5027), .C(w5026), .Q(w5246) );
	vdp_slatch g5125 (.D(S[7]), .nC(w5029), .C(w5030), .Q(w5281) );
	vdp_slatch g5126 (.D(S[7]), .nC(w5027), .C(w5026), .Q(w5211) );
	vdp_slatch g5127 (.D(REG_BUS[2]), .nC(w5251), .C(w5252), .Q(w5249) );
	vdp_slatch g5128 (.D(REG_BUS[5]), .nC(w5251), .C(w5252), .Q(w5245) );
	vdp_bufif0 g5129 (.A(w5232), .Z(VRAMA[9]), .nE(w5183) );
	vdp_bufif0 g5130 (.A(w5179), .Z(VRAMA[10]), .nE(w5214) );
	vdp_bufif0 g5131 (.A(w5270), .Z(VRAMA[10]), .nE(w5183) );
	vdp_bufif0 g5132 (.A(w5233), .Z(VRAMA[13]), .nE(w5183) );
	vdp_bufif0 g5133 (.A(w5276), .Z(VRAMA[14]), .nE(w5214) );
	vdp_bufif0 g5134 (.A(w5232), .Z(VRAMA[11]), .nE(w5214) );
	vdp_bufif0 g5135 (.A(w5269), .Z(VRAMA[13]), .nE(w5214) );
	vdp_bufif0 g5136 (.A(w5270), .Z(VRAMA[12]), .nE(w5214) );
	vdp_bufif0 g5137 (.A(w5269), .Z(VRAMA[11]), .nE(w5183) );
	vdp_bufif0 g5138 (.A(w5276), .Z(VRAMA[12]), .nE(w5183) );
	vdp_bufif0 g5139 (.A(w5233), .Z(VRAMA[15]), .nE(w5214) );
	vdp_slatch g5140 (.D(REG_BUS[3]), .nC(w5292), .C(w5291), .Q(w5270) );
	vdp_slatch g5141 (.D(REG_BUS[4]), .nC(w5292), .C(w5291), .Q(w5269) );
	vdp_xor g5142 (.Z(w5231), .B(w5269), .A(VRAMA[13]) );
	vdp_xor g5143 (.Z(w5230), .B(w5270), .A(VRAMA[12]) );
	vdp_dlatch_inv g5144 (.nQ(w5268), .D(w5273), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5145 (.nQ(w5267), .D(w5274), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5146 (.nQ(w5266), .D(w6702), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5147 (.nQ(w5265), .D(w6704), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5148 (.nQ(w5264), .D(w5275), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5149 (.nQ(w5263), .D(w5272), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5150 (.nQ(w5262), .D(w6703), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5151 (.nQ(w6378), .D(w5271), .nC(nDCLK1), .C(DCLK1) );
	vdp_comp_we g5152 (.nZ(w5293), .A(w5178), .Z(w5294) );
	vdp_comp_we g5153 (.nZ(w5119), .A(w5178), .Z(w6587) );
	vdp_comp_we g5154 (.nZ(w5290), .A(w5178), .Z(w6588) );
	vdp_comp_we g5155 (.nZ(w5289), .A(w5178), .Z(w6589) );
	vdp_comp_we g5156 (.nZ(w5288), .A(w5178), .Z(w6590) );
	vdp_comp_we g5157 (.nZ(w5287), .A(w5178), .Z(w6591) );
	vdp_comp_we g5158 (.nZ(w5286), .A(w5178), .Z(w6592) );
	vdp_comp_we g5159 (.nZ(w5285), .A(w5178), .Z(w6593) );
	vdp_comp_we g5160 (.nZ(w5284), .A(w5178), .Z(w6594) );
	vdp_comp_we g5161 (.nZ(w6596), .A(w5178), .Z(w6595) );
	vdp_comp_we g5162 (.nZ(w5282), .A(w119), .Z(w5283) );
	vdp_noif0 g5163 (.A(w5221), .nZ(VRAMA[10]), .nE(w5142) );
	vdp_noif0 g5164 (.A(w5250), .nZ(VRAMA[13]), .nE(w5142) );
	vdp_noif0 g5165 (.A(w5280), .nZ(VRAMA[11]), .nE(w5142) );
	vdp_noif0 g5166 (.A(w5279), .nZ(VRAMA[12]), .nE(w5142) );
	vdp_not g5167 (.nZ(w5223), .A(VRAMA[2]) );
	vdp_not g5168 (.nZ(w5250), .A(w5249) );
	vdp_not g5169 (.nZ(w5278), .A(w124) );
	vdp_aoi22 g5170 (.Z(w4981), .B2(w5211), .B1(w5222), .A1(w5082), .A2(w5234) );
	vdp_aoi22 g5171 (.Z(w5221), .B2(w5211), .B1(w5247), .A1(w5082), .A2(w5226) );
	vdp_aoi22 g5172 (.Z(w4974), .B2(w5211), .B1(w5235), .A1(w5082), .A2(w6580) );
	vdp_aoi22 g5173 (.Z(w5280), .B2(w5211), .B1(w5248), .A1(w5082), .A2(w5246) );
	vdp_aoi22 g5174 (.Z(w5279), .B2(w5211), .B1(w5281), .A1(w5082), .A2(w5211) );
	vdp_and g5175 (.Z(w5277), .B(w5278), .A(w4557) );
	vdp_nor8 g5176 (.Z(w5220), .B(w5230), .A(w5231), .C(w5229), .D(w5228), .F(w5217), .E(w5213), .G(w5215), .H(w5216) );
	vdp_not g5177 (.nZ(w5295), .A(w123) );
	vdp_comp_str g5178 (.nZ(w5292), .A(w142), .Z(w5291) );
	vdp_comp_str g5179 (.nZ(w5252), .A(w143), .Z(w5251) );
	vdp_or3 g5180 (.Z(w5178), .B(w119), .A(w123), .C(w5277) );
	vdp_not g5181 (.nZ(S[7]), .A(w5268) );
	vdp_not g5182 (.nZ(S[6]), .A(w5267) );
	vdp_not g5183 (.nZ(S[5]), .A(w5266) );
	vdp_not g5184 (.nZ(S[4]), .A(w5265) );
	vdp_not g5185 (.nZ(S[3]), .A(w5264) );
	vdp_not g5186 (.nZ(S[2]), .A(w5263) );
	vdp_not g5187 (.nZ(S[1]), .A(w5262) );
	vdp_not g5188 (.nZ(S[0]), .A(w6378) );
	vdp_aon21_sr g5189 (.Q(w5371), .A1(w5370), .A2(w6481), .B(w6488), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5190 (.Q(w6488), .A1(w5338), .A2(w6481), .B(w6487), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5191 (.Q(w6487), .A1(w5337), .A2(w6481), .B(w6486), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5192 (.Q(w6486), .A1(w5336), .A2(w6481), .B(w6485), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5193 (.Q(w6485), .A1(w5335), .A2(w6481), .B(w6484), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5194 (.Q(w6484), .A1(w5334), .A2(w6481), .B(w6483), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5195 (.Q(w6483), .A1(w5333), .A2(w6481), .B(w6482), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5196 (.Q(w6482), .A1(w5332), .A2(w6481), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5197 (.Q(w6490), .A1(w5327), .A2(w6489), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5198 (.Q(w6491), .A1(w5326), .A2(w6489), .B(w6490), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5199 (.Q(w6492), .A1(w5325), .A2(w6489), .B(w6491), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5200 (.Q(w6493), .A1(w5324), .A2(w6489), .B(w6492), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5201 (.Q(w6494), .A1(w5323), .A2(w6489), .B(w6493), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5202 (.Q(w6495), .A1(w5322), .A2(w6489), .B(w6494), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5203 (.Q(w6496), .A1(w5321), .A2(w6489), .B(w6495), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5204 (.Q(w5352), .A1(w5341), .A2(w6489), .B(w6496), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5205 (.Q(w5479), .A1(w5316), .A2(w6473), .B(w6474), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5206 (.Q(w6474), .A1(w5315), .A2(w6473), .B(w6475), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5207 (.Q(w6475), .A1(w5314), .A2(w6473), .B(w6476), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5208 (.Q(w6476), .A1(w5313), .A2(w6473), .B(w6477), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5209 (.Q(w6477), .A1(w5312), .A2(w6473), .B(w6478), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5210 (.Q(w6478), .A1(w5311), .A2(w6473), .B(w6479), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5211 (.Q(w6479), .A1(w5310), .A2(w6473), .B(w6480), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5212 (.Q(w6480), .A1(w5309), .A2(w6473), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5213 (.Q(w6466), .A1(w5304), .A2(w6465), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5214 (.Q(w6467), .A1(w5303), .A2(w6465), .B(w6466), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5215 (.Q(w6468), .A1(w5302), .A2(w6465), .B(w6467), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5216 (.Q(w6469), .A1(w5301), .A2(w6465), .B(w6468), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5217 (.Q(w6471), .A1(w5379), .A2(w6465), .B(w6469), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5218 (.Q(w6470), .A1(w5384), .A2(w6465), .B(w6471), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5219 (.Q(w6472), .A1(w5378), .A2(w6465), .B(w6470), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5220 (.Q(w5300), .A1(w5299), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .A2(w6465), .B(w6472) );
	vdp_not g5221 (.nZ(w6473), .A(w5364) );
	vdp_not g5222 (.nZ(w6465), .A(w5364) );
	vdp_not g5223 (.nZ(w6489), .A(w5364) );
	vdp_not g5224 (.nZ(w6481), .A(w5364) );
	vdp_or4 g5225 (.Z(w5369), .B(w5330), .A(w5387), .D(w5365), .C(w5331) );
	vdp_or4 g5226 (.Z(w5356), .B(w5328), .A(w5359), .D(w5363), .C(w5329) );
	vdp_or4 g5227 (.Z(w5372), .B(w5340), .A(w5299), .D(w5718), .C(w5339) );
	vdp_or4 g5228 (.Z(w5355), .B(w5320), .A(w5714), .D(w5378), .C(w5319) );
	vdp_or4 g5229 (.Z(w5351), .B(w5318), .A(w5713), .D(w5384), .C(w5317) );
	vdp_or4 g5230 (.Z(w5375), .B(w5306), .A(w5305), .D(w6379), .C(w5307) );
	vdp_or4 g5231 (.Z(w5346), .B(w5344), .A(w5345), .D(w5308), .C(w5343) );
	vdp_slatch g5232 (.Q(w5365), .D(w5424), .nC(w5360), .C(w5361) );
	vdp_comp_str g5233 (.nZ(w5360), .A(w5395), .Z(w5361) );
	vdp_slatch g5234 (.Q(w5331), .D(w5422), .nC(w5360), .C(w5361) );
	vdp_slatch g5235 (.Q(w5330), .D(w5421), .nC(w5360), .C(w5361) );
	vdp_slatch g5236 (.Q(w5387), .D(w5420), .nC(w5360), .C(w5361) );
	vdp_slatch g5237 (.Q(w5363), .D(w5419), .nC(w5360), .C(w5361) );
	vdp_slatch g5238 (.Q(w5329), .D(w5418), .nC(w5360), .C(w5361) );
	vdp_slatch g5239 (.Q(w5328), .D(w5416), .nC(w5360), .C(w5361) );
	vdp_slatch g5240 (.Q(w5359), .D(w5412), .nC(w5360), .C(w5361) );
	vdp_slatch g5241 (.Q(w5308), .D(w6462), .nC(w5342), .C(w5377) );
	vdp_slatch g5242 (.Q(w5343), .D(w6463), .nC(w5342), .C(w5377) );
	vdp_slatch g5243 (.Q(w5344), .D(w6464), .nC(w5342), .C(w5377) );
	vdp_slatch g5244 (.Q(w5345), .D(w5401), .nC(w5342), .C(w5377) );
	vdp_slatch g5245 (.Q(w6379), .D(w5399), .nC(w5342), .C(w5377) );
	vdp_slatch g5246 (.Q(w5307), .D(w5398), .nC(w5342), .C(w5377) );
	vdp_slatch g5247 (.Q(w5306), .D(w5397), .nC(w5342), .C(w5377) );
	vdp_slatch g5248 (.Q(w5305), .D(w5394), .nC(w5342), .C(w5377) );
	vdp_aon22 g5249 (.Z(w5432), .B2(w5348), .B1(w5382), .A1(w5375), .A2(w5354) );
	vdp_comp_we g5250 (.nZ(w5348), .A(w5381), .Z(w5354) );
	vdp_notif0 g5251 (.A(w5376), .nZ(DB[11]), .nE(w5393) );
	vdp_notif0 g5252 (.A(w5380), .nZ(DB[3]), .nE(w5393) );
	vdp_notif0 g5253 (.A(w5349), .nZ(DB[10]), .nE(w5404) );
	vdp_notif0 g5254 (.A(w5350), .nZ(DB[2]), .nE(w5404) );
	vdp_notif0 g5255 (.A(w5358), .nZ(DB[1]), .nE(w5404) );
	vdp_notif0 g5256 (.A(w5385), .nZ(DB[9]), .nE(w5404) );
	vdp_notif0 g5257 (.A(w5367), .nZ(DB[8]), .nE(w5404) );
	vdp_notif0 g5258 (.A(w5368), .nZ(DB[0]), .nE(w5404) );
	vdp_not g5259 (.nZ(w5373), .A(w5372) );
	vdp_aon22 g5260 (.Z(w5405), .B2(w5348), .B1(w5353), .A1(w5346), .A2(w5354) );
	vdp_aon22 g5261 (.Z(w5410), .B2(w5348), .B1(w5357), .A1(w5356), .A2(w5354) );
	vdp_aon22 g5262 (.Z(w5427), .B2(w5348), .B1(w5373), .A1(w5369), .A2(w5354) );
	vdp_comp_str g5263 (.nZ(w5342), .A(w5395), .Z(w5377) );
	vdp_not g5264 (.nZ(w5382), .A(w5383) );
	vdp_not g5265 (.nZ(w5353), .A(w5351) );
	vdp_not g5266 (.nZ(w5357), .A(w5355) );
	vdp_and3 g5267 (.Z(w5814), .B(w5408), .A(w5356), .C(w5355) );
	vdp_and3 g5268 (.Z(w5414), .B(w5428), .A(w5369), .C(w5372) );
	vdp_and3 g5269 (.Z(w5430), .B(w5406), .A(w5346), .C(w5351) );
	vdp_and3 g5270 (.Z(w5771), .B(w5375), .A(w5388), .C(w5383) );
	vdp_aon2222 g5271 (.Z(w5380), .B2(w5301), .B1(w5391), .A1(w5392), .A2(w5303), .D2(w5299), .D1(w5389), .C1(w5390), .C2(w5384) );
	vdp_aon2222 g5272 (.Z(w5376), .B2(w5302), .B1(w5391), .A1(w5392), .A2(w5304), .D2(w5378), .D1(w5389), .C1(w5390), .C2(w5379) );
	vdp_aon2222 g5273 (.Z(w5349), .B2(w5311), .B1(w5391), .A1(w5392), .A2(w5309), .D2(w5315), .D1(w5389), .C1(w5390), .C2(w5313) );
	vdp_aon2222 g5274 (.Z(w5350), .B2(w5312), .B1(w5391), .A1(w5392), .A2(w5310), .D2(w5316), .D1(w5389), .C1(w5390), .C2(w5314) );
	vdp_aon2222 g5275 (.Z(w5358), .B2(w5324), .B1(w5391), .A1(w5392), .A2(w5326), .D2(w5341), .D1(w5389), .C1(w5390), .C2(w5322) );
	vdp_aon2222 g5276 (.Z(w5385), .B2(w5325), .B1(w5391), .A1(w5392), .A2(w5327), .D2(w5321), .D1(w5389), .C1(w5390), .C2(w5323) );
	vdp_aon2222 g5277 (.Z(w5367), .B2(w5334), .B1(w5391), .A1(w5392), .A2(w5332), .D2(w5338), .D1(w5389), .C1(w5390), .C2(w5336) );
	vdp_aon2222 g5278 (.Z(w5368), .B2(w5335), .B1(w5391), .A1(w5392), .A2(w5333), .D2(w5370), .D1(w5389), .C1(w5390), .C2(w5337) );
	vdp_slatch g5279 (.Q(w5424), .D(w5445), .nC(w5444), .C(w5423) );
	vdp_comp_str g5280 (.nZ(w5444), .A(w5443), .Z(w5423) );
	vdp_slatch g5281 (.Q(w5422), .D(w5449), .nC(w5444), .C(w5423) );
	vdp_slatch g5282 (.Q(w5421), .D(w5450), .nC(w5444), .C(w5423) );
	vdp_slatch g5283 (.Q(w5420), .D(w5453), .nC(w5444), .C(w5423) );
	vdp_slatch g5284 (.Q(w5419), .D(w5458), .nC(w5459), .C(w5417) );
	vdp_comp_str g5285 (.nZ(w5459), .A(w5454), .Z(w5417) );
	vdp_slatch g5286 (.Q(w5418), .D(w5461), .nC(w5459), .C(w5417) );
	vdp_slatch g5287 (.Q(w5416), .D(w5462), .nC(w5459), .C(w5417) );
	vdp_slatch g5288 (.Q(w5412), .D(w5464), .nC(w5459), .C(w5417) );
	vdp_sr_bit g5289 (.Q(w5466), .D(w5352), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5290 (.nQ(w5411), .D(w5469), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5291 (.nQ(w5471), .D(w5409), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5292 (.nQ(w5407), .D(w5478), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5293 (.nQ(w5484), .D(w6420), .nC(nDCLK2), .C(DCLK2) );
	vdp_slatch g5294 (.Q(w5401), .D(w5445), .nC(w5486), .C(w5403) );
	vdp_slatch g5295 (.Q(w6462), .D(w5449), .nC(w5486), .C(w5403) );
	vdp_slatch g5296 (.Q(w6463), .D(w5450), .nC(w5486), .C(w5403) );
	vdp_slatch g5297 (.Q(w6464), .D(w5453), .nC(w5486), .C(w5403) );
	vdp_comp_str g5298 (.nZ(w5486), .A(w5485), .Z(w5403) );
	vdp_slatch g5299 (.Q(w5399), .D(w5458), .nC(w5497), .C(w5396) );
	vdp_slatch g5300 (.Q(w5398), .D(w5461), .nC(w5497), .C(w5396) );
	vdp_slatch g5301 (.Q(w5397), .D(w5462), .nC(w5497), .C(w5396) );
	vdp_slatch g5302 (.Q(w5394), .D(w5464), .nC(w5497), .C(w5396) );
	vdp_comp_str g5303 (.nZ(w5497), .A(w5502), .Z(w5396) );
	vdp_dlatch_inv g5304 (.nQ(w5495), .D(w5494), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5305 (.nQ(w5498), .D(w6419), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5306 (.nQ(w5431), .D(w5501), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5307 (.Z(w5500), .B(w5431), .A(w5436) );
	vdp_xor g5308 (.Z(w6458), .B(w5407), .A(w5436) );
	vdp_xor g5309 (.Z(w5467), .B(w5411), .A(w5436) );
	vdp_xor g5310 (.Z(w6387), .B(w6386), .A(w5436) );
	vdp_sr_bit g5311 (.Q(w6461), .D(w5371), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5312 (.nQ(w6386), .D(w5434), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5313 (.nQ(w6388), .D(w5426), .nC(nDCLK2), .C(DCLK2) );
	vdp_and g5314 (.Z(w5428), .B(w6387), .A(w5437) );
	vdp_and g5315 (.Z(w5429), .B(w6388), .A(DCLK1) );
	vdp_and g5316 (.Z(w5413), .B(w5471), .A(DCLK1) );
	vdp_and g5317 (.Z(w5408), .B(w5467), .A(w5437) );
	vdp_and g5318 (.Z(w5389), .B(w5473), .A(w5472) );
	vdp_and g5319 (.Z(w5390), .B(w82), .A(w5473) );
	vdp_and g5320 (.Z(w5391), .B(w83), .A(w5472) );
	vdp_and g5321 (.Z(w5392), .B(w82), .A(w83) );
	vdp_and g5322 (.Z(w5406), .B(w6458), .A(w83) );
	vdp_and g5323 (.Z(w5425), .B(w5484), .A(DCLK1) );
	vdp_and g5324 (.Z(w5415), .B(w5498), .A(DCLK1) );
	vdp_and g5325 (.Z(w5388), .B(w5500), .A(w5437) );
	vdp_sr_bit g5326 (.Q(w5476), .D(w5479), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5327 (.Q(w5487), .D(w5456), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_not g5328 (.nZ(w5395), .A(w5402) );
	vdp_not g5329 (.nZ(w5400), .A(w4505) );
	vdp_not g5330 (.nZ(w5472), .A(w82) );
	vdp_not g5331 (.nZ(w5473), .A(w83) );
	vdp_aoi21 g5332 (.Z(w5426), .B(w5440), .A1(w5427), .A2(w5428) );
	vdp_aoi21 g5333 (.Z(w5409), .B(w5468), .A1(w5410), .A2(w5408) );
	vdp_aoi21 g5334 (.Z(w6420), .B(w5483), .A1(w5405), .A2(w5406) );
	vdp_oai21 g5335 (.Z(w5402), .B(DCLK2), .A1(w5488), .A2(w5487) );
	vdp_aoi21 g5336 (.Z(w6419), .B(w5483), .A1(w5388), .A2(w5432) );
	vdp_not g5337 (.nZ(w5393), .A(w121) );
	vdp_nand g5338 (.Z(w5456), .B(w5495), .A(w5400) );
	vdp_sr_bit g5339 (.Q(w5447), .D(w5504), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5340 (.Q(w5452), .D(w6389), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5341 (.Q(w5463), .D(w6460), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5342 (.Q(w5448), .D(w5465), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5343 (.Q(w5470), .D(w2706), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5344 (.Q(w5474), .D(w5475), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5345 (.Q(w6430), .D(w5491), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5346 (.Q(w5491), .D(w5503), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5347 (.Q(w5506), .D(w5300), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon22 g5348 (.Z(w5503), .B2(w5300), .B1(w5510), .A1(w5509), .A2(w5506) );
	vdp_aon22 g5349 (.Z(w5475), .B2(w5479), .B1(w5510), .A1(w5509), .A2(w5476) );
	vdp_aon22 g5350 (.Z(w5465), .B2(w5352), .B1(w5510), .A1(w5509), .A2(w5466) );
	vdp_aon22 g5351 (.Z(w5504), .B2(w5371), .B1(w5510), .A1(w5509), .A2(w6461) );
	vdp_not g5352 (.nZ(w5446), .A(w5501) );
	vdp_not g5353 (.nZ(w5438), .A(w83) );
	vdp_not g5354 (.nZ(w5443), .A(w5522) );
	vdp_not g5355 (.nZ(w5451), .A(M5) );
	vdp_not g5356 (.nZ(w5454), .A(w5455) );
	vdp_not g5357 (.nZ(w5441), .A(w5515) );
	vdp_not g5358 (.nZ(w5435), .A(w5513) );
	vdp_not g5359 (.nZ(w5485), .A(w5482) );
	vdp_not g5360 (.nZ(w5502), .A(w5490) );
	vdp_not g5361 (.nZ(w5496), .A(w5491) );
	vdp_comp_we g5362 (.nZ(w5510), .A(M5), .Z(w5509) );
	vdp_and g5363 (.Z(w2824), .B(w5448), .A(w5447) );
	vdp_or g5364 (.Z(w6389), .B(w5447), .A(w5451) );
	vdp_or g5365 (.Z(w5457), .B(w5460), .A(w5456) );
	vdp_and g5366 (.Z(w6460), .B(w5448), .A(M5) );
	vdp_and g5367 (.Z(w2706), .B(w5474), .A(M5) );
	vdp_or g5368 (.Z(w5499), .B(w5456), .A(w5489) );
	vdp_not g5369 (.nZ(w5521), .A(SPR_PRIO) );
	vdp_bufif0 g5370 (.A(w6430), .Z(COL[0]), .nE(w5521) );
	vdp_oai21 g5371 (.Z(w5482), .B(DCLK2), .A1(w5457), .A2(w5481) );
	vdp_bufif0 g5372 (.A(w5470), .Z(COL[6]), .nE(w5521) );
	vdp_bufif0 g5373 (.A(w5463), .Z(COL[5]), .nE(w5521) );
	vdp_bufif0 g5374 (.A(w5452), .Z(COL[4]), .nE(w5521) );
	vdp_oai21 g5375 (.Z(w5455), .B(DCLK2), .A1(w5457), .A2(w5442) );
	vdp_oai21 g5376 (.Z(w5522), .B(DCLK2), .A1(w5516), .A2(w5442) );
	vdp_and3 g5377 (.Z(w5442), .B(w5520), .A(w5441), .C(w5519) );
	vdp_and3 g5378 (.Z(w5460), .B(w5520), .A(w5441), .C(w5507) );
	vdp_and3 g5379 (.Z(w5481), .B(w5519), .A(w5508), .C(w5441) );
	vdp_and3 g5380 (.Z(w5489), .B(w5507), .A(w5508), .C(w5441) );
	vdp_or4 g5381 (.Z(w2705), .B(w5512), .A(w5493), .D(w5491), .C(w5492) );
	vdp_and4 g5382 (.Z(w2765), .B(w5492), .A(w5512), .D(w5496), .C(w5493) );
	vdp_and4 g5383 (.Z(w2764), .B(w5492), .A(w5512), .D(w5491), .C(w5493) );
	vdp_oai21 g5384 (.Z(w5490), .B(DCLK2), .A1(w5481), .A2(w5499) );
	vdp_nand3 g5385 (.Z(w5434), .B(w5435), .A(w5446), .C(w5518) );
	vdp_nand3 g5386 (.Z(w5439), .B(w5517), .A(w120), .C(w5438) );
	vdp_nand3 g5387 (.Z(w5480), .B(w82), .A(w120), .C(w5438) );
	vdp_nand g5388 (.Z(w5483), .B(w5480), .A(w5511) );
	vdp_nand g5389 (.Z(w5477), .B(w5514), .A(w5513) );
	vdp_nand g5390 (.Z(w5478), .B(w5446), .A(w5477) );
	vdp_nand g5391 (.Z(w5469), .B(w5435), .A(w5446) );
	vdp_nand g5392 (.Z(w5440), .B(w5439), .A(w5511) );
	vdp_sr_bit g5393 (.Q(w6392), .D(w6391), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5394 (.Q(w6393), .D(w6392), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5395 (.Q(w5589), .D(w6393), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5396 (.Q(w5596), .D(w5589), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5397 (.Q(w5587), .D(w6394), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5398 (.Q(w6459), .D(nDCLK2), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5399 (.Q(w5598), .D(w6497), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5400 (.Q(w5579), .D(w6390), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_dlatch_inv g5401 (.nQ(w5545), .D(w5537), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5402 (.nQ(w5550), .D(w5536), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5403 (.nQ(w5556), .D(w5535), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5404 (.nQ(w5561), .D(w5534), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5405 (.nQ(w5562), .D(w5533), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5406 (.nQ(w5565), .D(w5532), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5407 (.nQ(w5566), .D(w5531), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5408 (.nQ(w5569), .D(w5529), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5409 (.nQ(w5593), .D(w5594), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5410 (.nQ(w5591), .D(w5574), .nC(nDCLK1), .C(DCLK1) );
	vdp_cnt_bit_load g5411 (.Q(w5594), .D(w5595), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1), .R(1'b0), .CI(w6499), .L(w5526), .nL(w5571) );
	vdp_cnt_bit_load g5412 (.Q(w5574), .D(w5573), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1), .R(1'b0), .CI(w5527), .L(w5526), .nL(w5571), .CO(w6499) );
	vdp_aon22 g5413 (.Z(w5458), .B2(w5528), .B1(DB[11]), .A1(w5569), .A2(w5546) );
	vdp_aon22 g5414 (.Z(w5529), .B2(w5530), .B1(w5558), .A1(w5557), .A2(w5549) );
	vdp_aon22 g5415 (.Z(w5461), .B2(w5528), .B1(DB[12]), .A1(w5566), .A2(w5546) );
	vdp_aon22 g5416 (.Z(w5531), .B2(w5530), .B1(w5554), .A1(w5555), .A2(w5549) );
	vdp_aon22 g5417 (.Z(w5462), .B2(w5528), .B1(DB[13]), .A1(w5565), .A2(w5546) );
	vdp_aon22 g5418 (.Z(w5532), .B2(w5530), .B1(w5547), .A1(w5548), .A2(w5549) );
	vdp_aon22 g5419 (.Z(w5464), .B2(w5528), .B1(DB[14]), .A1(w5562), .A2(w5546) );
	vdp_aon22 g5420 (.Z(w5533), .B2(w5530), .B1(w5538), .A1(w5539), .A2(w5549) );
	vdp_aon22 g5421 (.Z(w5445), .B2(w5528), .B1(DB[3]), .A1(w5561), .A2(w5546) );
	vdp_aon22 g5422 (.Z(w5534), .B2(w5530), .B1(w5557), .A1(w5558), .A2(w5549) );
	vdp_aon22 g5423 (.Z(w5449), .B2(w5528), .B1(DB[4]), .A1(w5556), .A2(w5546) );
	vdp_aon22 g5424 (.Z(w5535), .B2(w5530), .B1(w5555), .A1(w5554), .A2(w5549) );
	vdp_aon22 g5425 (.Z(w5450), .B2(w5528), .B1(DB[5]), .A1(w5550), .A2(w5546) );
	vdp_aon22 g5426 (.Z(w5536), .B2(w5530), .B1(w5548), .A1(w5547), .A2(w5549) );
	vdp_aon22 g5427 (.Z(w5453), .B2(w5528), .B1(DB[6]), .A1(w5545), .A2(w5546) );
	vdp_aon22 g5428 (.Z(w5537), .B2(w5530), .B1(w5539), .A1(w5538), .A2(w5549) );
	vdp_slatch g5429 (.Q(w6390), .D(w5582), .nC(w5525), .C(w5583) );
	vdp_dlatch_inv g5430 (.nQ(w5580), .D(w5579), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5431 (.nQ(nDCLK2), .D(w26), .nC(nHCLK1), .C(HCLK1) );
	vdp_xnor g5432 (.Z(w5508), .B(1'b0), .A(w5591) );
	vdp_xor g5433 (.Z(w5570), .B(w5579), .A(w5581) );
	vdp_aon22 g5434 (.Z(w6497), .B2(w5589), .B1(M5), .A1(w5596), .A2(w6498) );
	vdp_not g5435 (.nZ(w5597), .A(nDCLK2) );
	vdp_not g5436 (.nZ(w6498), .A(M5) );
	vdp_not g5437 (.nZ(w5525), .A(w5583) );
	vdp_not g5438 (.nZ(w6391), .A(w5586) );
	vdp_not g5439 (.nZ(w5507), .A(w5580) );
	vdp_not g5440 (.nZ(w5515), .A(w5593) );
	vdp_not g5441 (.nZ(w5527), .A(w5583) );
	vdp_comp_we g5442 (.nZ(w5546), .A(w4505), .Z(w5528) );
	vdp_comp_we g5443 (.nZ(w5549), .A(w5570), .Z(w5530) );
	vdp_comp_we g5444 (.nZ(w5571), .A(w5583), .Z(w5526) );
	vdp_and g5445 (.Z(w6394), .B(w6459), .A(w5597) );
	vdp_aoi21 g5446 (.Z(w5586), .B(w25), .A1(M5), .A2(w22) );
	vdp_sr_bit g5447 (.Q(w5581), .D(w5644), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_aon22 g5448 (.Z(w5652), .B2(w5646), .B1(w5645), .A1(w5642), .A2(w5590) );
	vdp_aon22 g5449 (.Z(w5651), .B2(w5646), .B1(w5649), .A1(w5647), .A2(w5590) );
	vdp_aon22 g5450 (.Z(w5648), .B2(w5646), .B1(w5647), .A1(w5649), .A2(w5590) );
	vdp_aon22 g5451 (.Z(w5653), .B2(w5646), .B1(w5642), .A1(w5645), .A2(w5590) );
	vdp_not g5452 (.nZ(w5608), .A(w5645) );
	vdp_not g5453 (.nZ(w5609), .A(w5649) );
	vdp_not g5454 (.nZ(w5614), .A(w5647) );
	vdp_not g5455 (.nZ(w5613), .A(w5642) );
	vdp_not g5456 (.nZ(w5541), .A(w5651) );
	vdp_not g5457 (.nZ(w5542), .A(w5652) );
	vdp_not g5458 (.nZ(w5543), .A(w5653) );
	vdp_not g5459 (.nZ(w5544), .A(w5648) );
	vdp_not g5460 (.nZ(w5588), .A(M5) );
	vdp_comp_we g5461 (.nZ(w5646), .A(w5581), .Z(w5590) );
	vdp_not g5462 (.nZ(w5583), .A(w5643) );
	vdp_not g5463 (.nZ(w5641), .A(w5640) );
	vdp_dlatch_inv g5464 (.nQ(w5640), .D(w5639), .nC(nHCLK1), .C(HCLK1) );
	vdp_aon2222 g5465 (.Z(w5540), .B2(w5542), .B1(w5602), .A1(w5601), .A2(w5541), .D2(w5544), .D1(w5620), .C1(w5618), .C2(w5543) );
	vdp_aon2222 g5466 (.Z(w5592), .B2(w5614), .B1(w5606), .A1(w5613), .A2(w5601), .D2(w5608), .D1(w5610), .C1(w5609), .C2(w5654) );
	vdp_aon2222 g5467 (.Z(w5560), .B2(w5542), .B1(w5607), .A1(w5606), .A2(w5541), .D2(w5544), .D1(w5611), .C1(w5619), .C2(w5543) );
	vdp_aon2222 g5468 (.Z(w5551), .B2(w5614), .B1(w5607), .A1(w5613), .A2(w5602), .D2(w5608), .D1(w5622), .C1(w5609), .C2(w5615) );
	vdp_aon2222 g5469 (.Z(w5568), .B2(w5542), .B1(w5615), .A1(w5654), .A2(w5541), .D2(w5544), .D1(w5617), .C1(w5616), .C2(w5543) );
	vdp_aon2222 g5470 (.Z(w5559), .B2(w5614), .B1(w5619), .A1(w5613), .A2(w5618), .D2(w5608), .D1(w5621), .C1(w5609), .C2(w5616) );
	vdp_aon2222 g5471 (.Z(w5578), .B2(w5542), .B1(w5622), .A1(w5610), .A2(w5541), .D2(w5544), .D1(w5623), .C1(w5621), .C2(w5543) );
	vdp_aon2222 g5472 (.Z(w5563), .B2(w5614), .B1(w5611), .A1(w5613), .A2(w5620), .D2(w5608), .D1(w5623), .C1(w5609), .C2(w5617) );
	vdp_aon2222 g5473 (.Z(w5552), .B2(w5542), .B1(w5625), .A1(w5624), .A2(w5541), .D2(w5544), .D1(w5637), .C1(w5626), .C2(w5543) );
	vdp_aon2222 g5474 (.Z(w5567), .B2(w5614), .B1(w5627), .A1(w5613), .A2(w5624), .D2(w5608), .D1(w5628), .C1(w5609), .C2(w5629) );
	vdp_aon2222 g5475 (.Z(w5564), .B2(w5542), .B1(w5631), .A1(w5627), .A2(w5541), .D2(w5544), .D1(w5630), .C1(w5632), .C2(w5543) );
	vdp_aon2222 g5476 (.Z(w5576), .B2(w5614), .B1(w5631), .A1(w5613), .A2(w5625), .D2(w5608), .D1(w5633), .C1(w5609), .C2(w5634) );
	vdp_aon2222 g5477 (.Z(w5575), .B2(w5542), .B1(w5634), .A1(w5629), .A2(w5541), .D2(w5544), .D1(w5635), .C1(w5636), .C2(w5543) );
	vdp_aon2222 g5478 (.Z(w5577), .B2(w5614), .B1(w5632), .A1(w5613), .A2(w5626), .D2(w5608), .D1(w5638), .C1(w5609), .C2(w5636) );
	vdp_aon2222 g5479 (.Z(w5585), .B2(w5542), .B1(w5633), .A1(w5628), .A2(w5541), .D2(w5544), .D1(w5650), .C1(w5638), .C2(w5543) );
	vdp_aon2222 g5480 (.Z(w5584), .B2(w5614), .B1(w5630), .A1(w5613), .A2(w5637), .D2(w5608), .D1(w5650), .C1(w5609), .C2(w5635) );
	vdp_aoi22 g5481 (.Z(w5538), .B2(w5600), .B1(w5540), .A1(w5553), .A2(w5592) );
	vdp_aoi22 g5482 (.Z(w5547), .B2(w5600), .B1(w5552), .A1(w5553), .A2(w5551) );
	vdp_aoi22 g5483 (.Z(w5554), .B2(w5600), .B1(w5560), .A1(w5553), .A2(w5559) );
	vdp_aoi22 g5484 (.Z(w5558), .B2(w5600), .B1(w5564), .A1(w5553), .A2(w5563) );
	vdp_aoi22 g5485 (.Z(w5539), .B2(w5600), .B1(w5568), .A1(w5553), .A2(w5567) );
	vdp_aoi22 g5486 (.Z(w5548), .B2(w5600), .B1(w5575), .A1(w5553), .A2(w5576) );
	vdp_aoi22 g5487 (.Z(w5555), .B2(w5600), .B1(w5578), .A1(w5553), .A2(w5577) );
	vdp_aoi22 g5488 (.Z(w5557), .B2(w5600), .B1(w5585), .A1(w5553), .A2(w5584) );
	vdp_nand g5489 (.Z(w5643), .B(w5641), .A(HCLK2) );
	vdp_nor g5490 (.Z(w5600), .B(w5588), .A(w5587) );
	vdp_nor g5491 (.Z(w5553), .B(M5), .A(w5587) );
	vdp_sr_bit g5492 (.Q(w5645), .D(w5649), .nC2(w5656), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5493 (.Q(w5649), .D(w5647), .nC2(w5656), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5494 (.Q(w5647), .D(w5642), .nC2(w5656), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5495 (.Q(w5642), .D(w5643), .nC2(w5656), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_dlatch_inv g5496 (.nQ(w5488), .D(w5645), .nC(nDCLK1), .C(DCLK1) );
	vdp_comp_str g5497 (.nZ(w5605), .A(w5657), .Z(w5659) );
	vdp_comp_str g5498 (.nZ(w5604), .A(w5657), .Z(w5662) );
	vdp_comp_str g5499 (.nZ(w5612), .A(w5657), .Z(w5663) );
	vdp_comp_str g5500 (.nZ(w5603), .A(w5657), .Z(w5658) );
	vdp_slatch g5501 (.D(w5672), .Q(w5601), .nC(w5603), .C(w5658) );
	vdp_slatch g5502 (.D(w6523), .Q(w5602), .nC(w5612), .C(w5663) );
	vdp_slatch g5503 (.D(w6522), .Q(w5618), .nC(w5604), .C(w5662) );
	vdp_slatch g5504 (.D(w6521), .Q(w5620), .nC(w5605), .C(w5659) );
	vdp_slatch g5505 (.D(w5671), .Q(w5606), .nC(w5603), .C(w5658) );
	vdp_slatch g5506 (.D(w6520), .Q(w5607), .nC(w5612), .C(w5663) );
	vdp_slatch g5507 (.D(w6519), .Q(w5619), .nC(w5604), .C(w5662) );
	vdp_slatch g5508 (.D(w6518), .Q(w5611), .nC(w5605), .C(w5659) );
	vdp_slatch g5509 (.D(w5670), .Q(w5654), .nC(w5603), .C(w5658) );
	vdp_slatch g5510 (.D(w6517), .Q(w5615), .nC(w5612), .C(w5663) );
	vdp_slatch g5511 (.D(w6516), .Q(w5616), .nC(w5604), .C(w5662) );
	vdp_slatch g5512 (.D(w6515), .Q(w5617), .nC(w5605), .C(w5659) );
	vdp_slatch g5513 (.D(w5669), .Q(w5610), .nC(w5603), .C(w5658) );
	vdp_slatch g5514 (.D(w6514), .Q(w5622), .nC(w5612), .C(w5663) );
	vdp_slatch g5515 (.D(w6513), .Q(w5621), .nC(w5604), .C(w5662) );
	vdp_slatch g5516 (.D(w6512), .Q(w5623), .nC(w5605), .C(w5659) );
	vdp_slatch g5517 (.D(w5668), .Q(w5624), .nC(w5603), .C(w5658) );
	vdp_slatch g5518 (.D(w6511), .Q(w5625), .nC(w5612), .C(w5663) );
	vdp_slatch g5519 (.D(w6510), .Q(w5626), .nC(w5604), .C(w5662) );
	vdp_slatch g5520 (.D(w6509), .Q(w5637), .nC(w5605), .C(w5659) );
	vdp_slatch g5521 (.D(w5667), .Q(w5627), .nC(w5603), .C(w5658) );
	vdp_slatch g5522 (.D(w6508), .Q(w5631), .nC(w5612), .C(w5663) );
	vdp_slatch g5523 (.D(w6507), .Q(w5632), .nC(w5604), .C(w5662) );
	vdp_slatch g5524 (.D(w6506), .Q(w5630), .nC(w5605), .C(w5659) );
	vdp_slatch g5525 (.D(w5666), .Q(w5629), .nC(w5603), .C(w5658) );
	vdp_slatch g5526 (.D(w6505), .Q(w5634), .nC(w5612), .C(w5663) );
	vdp_slatch g5527 (.D(w6504), .Q(w5636), .nC(w5604), .C(w5662) );
	vdp_slatch g5528 (.D(w6503), .Q(w5635), .nC(w5605), .C(w5659) );
	vdp_slatch g5529 (.D(w5665), .Q(w5628), .nC(w5603), .C(w5658) );
	vdp_slatch g5530 (.D(w6502), .Q(w5633), .nC(w5612), .C(w5663) );
	vdp_slatch g5531 (.D(w6501), .Q(w5638), .nC(w5604), .C(w5662) );
	vdp_slatch g5532 (.D(w6500), .nC(w5605), .C(w5659), .Q(w5650) );
	vdp_sr_bit g5533 (.Q(w5673), .D(w5674), .nC2(nDCLK1), .nC1(w5656), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g5534 (.Q(w6395), .D(w5673), .nC2(nDCLK1), .nC1(w5656), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g5535 (.Q(w5687), .D(w6395), .nC2(nDCLK1), .nC1(w5656), .C2(DCLK1), .C1(DCLK2) );
	vdp_comp_str g5536 (.nZ(w5677), .A(w5688), .Z(w5664) );
	vdp_comp_str g5537 (.nZ(w5680), .A(w5688), .Z(w5661) );
	vdp_comp_str g5538 (.nZ(w5682), .A(w5688), .Z(w5660) );
	vdp_dlatch_inv g5539 (.nQ(w5674), .D(w5683), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g5540 (.Z(w5657), .B(DCLK2), .A(w5687) );
	vdp_and g5541 (.Z(w5688), .B(DCLK2), .A(w5673) );
	vdp_and g5542 (.Z(w5689), .B(DCLK2), .A(w5674) );
	vdp_slatch g5543 (.Q(w6502), .D(w6526), .nC(w5677), .C(w5664) );
	vdp_slatch g5544 (.Q(w6501), .D(w6525), .nC(w5680), .C(w5661) );
	vdp_slatch g5545 (.Q(w6500), .D(w6524), .nC(w5682), .C(w5660) );
	vdp_slatch g5546 (.Q(w6505), .D(w6529), .nC(w5677), .C(w5664) );
	vdp_slatch g5547 (.Q(w6504), .D(w6528), .nC(w5680), .C(w5661) );
	vdp_slatch g5548 (.Q(w6503), .D(w6527), .nC(w5682), .C(w5660) );
	vdp_slatch g5549 (.Q(w6508), .D(w6532), .nC(w5677), .C(w5664) );
	vdp_slatch g5550 (.Q(w6507), .D(w6531), .nC(w5680), .C(w5661) );
	vdp_slatch g5551 (.Q(w6506), .D(w6530), .nC(w5682), .C(w5660) );
	vdp_slatch g5552 (.Q(w6511), .D(w6535), .nC(w5677), .C(w5664) );
	vdp_slatch g5553 (.Q(w6510), .D(w6534), .nC(w5680), .C(w5661) );
	vdp_slatch g5554 (.Q(w6509), .D(w6533), .nC(w5682), .C(w5660) );
	vdp_slatch g5555 (.Q(w6514), .D(w6538), .nC(w5677), .C(w5664) );
	vdp_slatch g5556 (.Q(w6513), .D(w6537), .nC(w5680), .C(w5661) );
	vdp_slatch g5557 (.Q(w6512), .D(w6536), .nC(w5682), .C(w5660) );
	vdp_slatch g5558 (.Q(w6517), .D(w6541), .nC(w5677), .C(w5664) );
	vdp_slatch g5559 (.Q(w6516), .D(w6540), .nC(w5680), .C(w5661) );
	vdp_slatch g5560 (.Q(w6515), .D(w6539), .nC(w5682), .C(w5660) );
	vdp_slatch g5561 (.Q(w6520), .D(w6544), .nC(w5677), .C(w5664) );
	vdp_slatch g5562 (.Q(w6519), .D(w6543), .nC(w5680), .C(w5661) );
	vdp_slatch g5563 (.Q(w6518), .D(w6542), .nC(w5682), .C(w5660) );
	vdp_slatch g5564 (.Q(w6523), .D(w6547), .nC(w5677), .C(w5664) );
	vdp_slatch g5565 (.Q(w6522), .D(w6546), .nC(w5680), .C(w5661) );
	vdp_slatch g5566 (.Q(w6521), .D(w6545), .nC(w5682), .C(w5660) );
	vdp_sr_bit g5567 (.Q(w5686), .D(w5685), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_dlatch_inv g5568 (.nQ(w5685), .D(w5684), .nC(nDCLK1), .C(DCLK1) );
	vdp_and g5569 (.Z(w5696), .B(w5685), .A(DCLK2) );
	vdp_nand g5570 (.Z(w5684), .B(w5589), .A(HCLK1) );
	vdp_nand g5571 (.Z(w5683), .B(w5598), .A(HCLK1) );
	vdp_and g5572 (.Z(w5695), .B(w5686), .A(DCLK2) );
	vdp_comp_str g5573 (.nZ(w5681), .A(w5696), .Z(w5694) );
	vdp_comp_str g5574 (.nZ(w5679), .A(w5695), .Z(w5693) );
	vdp_comp_str g5575 (.nZ(w5678), .A(w5689), .Z(w5692) );
	vdp_comp_str g5576 (.nZ(w5676), .A(w5688), .Z(w5691) );
	vdp_slatch g5577 (.D(S[7]), .Q(w5672), .nC(w5676), .C(w5691) );
	vdp_slatch g5578 (.D(S[7]), .Q(w6547), .nC(w5678), .C(w5692) );
	vdp_slatch g5579 (.D(S[7]), .Q(w6546), .nC(w5679), .C(w5693) );
	vdp_slatch g5580 (.D(S[7]), .Q(w6545), .nC(w5681), .C(w5694) );
	vdp_slatch g5581 (.D(S[5]), .Q(w5671), .nC(w5676), .C(w5691) );
	vdp_slatch g5582 (.D(S[5]), .Q(w6544), .nC(w5678), .C(w5692) );
	vdp_slatch g5583 (.D(S[5]), .Q(w6543), .nC(w5679), .C(w5693) );
	vdp_slatch g5584 (.D(S[5]), .Q(w6542), .nC(w5681), .C(w5694) );
	vdp_slatch g5585 (.D(S[3]), .Q(w5670), .nC(w5676), .C(w5691) );
	vdp_slatch g5586 (.D(S[3]), .Q(w6541), .nC(w5678), .C(w5692) );
	vdp_slatch g5587 (.D(S[3]), .Q(w6540), .nC(w5679), .C(w5693) );
	vdp_slatch g5588 (.D(S[3]), .Q(w6539), .nC(w5681), .C(w5694) );
	vdp_slatch g5589 (.D(S[1]), .Q(w5669), .nC(w5676), .C(w5691) );
	vdp_slatch g5590 (.D(S[1]), .Q(w6538), .nC(w5678), .C(w5692) );
	vdp_slatch g5591 (.D(S[1]), .Q(w6537), .nC(w5679), .C(w5693) );
	vdp_slatch g5592 (.D(S[1]), .Q(w6536), .nC(w5681), .C(w5694) );
	vdp_slatch g5593 (.D(S[6]), .Q(w5668), .nC(w5676), .C(w5691) );
	vdp_slatch g5594 (.D(S[6]), .Q(w6535), .nC(w5678), .C(w5692) );
	vdp_slatch g5595 (.D(S[6]), .Q(w6534), .nC(w5679), .C(w5693) );
	vdp_slatch g5596 (.D(S[6]), .Q(w6533), .nC(w5681), .C(w5694) );
	vdp_slatch g5597 (.D(S[4]), .Q(w5667), .nC(w5676), .C(w5691) );
	vdp_slatch g5598 (.D(S[4]), .Q(w6532), .nC(w5678), .C(w5692) );
	vdp_slatch g5599 (.D(S[4]), .Q(w6531), .nC(w5679), .C(w5693) );
	vdp_slatch g5600 (.D(S[4]), .Q(w6530), .nC(w5681), .C(w5694) );
	vdp_slatch g5601 (.D(S[2]), .Q(w5666), .nC(w5676), .C(w5691) );
	vdp_slatch g5602 (.D(S[2]), .Q(w6529), .nC(w5678), .C(w5692) );
	vdp_slatch g5603 (.D(S[2]), .Q(w6528), .nC(w5679), .C(w5693) );
	vdp_slatch g5604 (.D(S[2]), .Q(w6527), .nC(w5681), .C(w5694) );
	vdp_slatch g5605 (.D(S[0]), .Q(w5665), .nC(w5676), .C(w5691) );
	vdp_slatch g5606 (.D(S[0]), .Q(w6526), .nC(w5678), .C(w5692) );
	vdp_slatch g5607 (.D(S[0]), .Q(w6525), .nC(w5679), .C(w5693) );
	vdp_slatch g5608 (.D(S[0]), .nC(w5681), .C(w5694), .Q(w6524) );
	vdp_aon21_sr g5609 (.Q(w5752), .A1(w5711), .A2(w6723), .B(w6434), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5610 (.Q(w6434), .A1(w5319), .A2(w6723), .B(w6435), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5611 (.Q(w6435), .A1(w5317), .A2(w6723), .B(w6436), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5612 (.Q(w6436), .A1(w5712), .A2(w6723), .B(w6437), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5613 (.Q(w6437), .A1(w5741), .A2(w6723), .B(w6438), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5614 (.Q(w6438), .A1(w5703), .A2(w6723), .B(w6433), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5615 (.Q(w6433), .A1(w5704), .A2(w6723), .B(w6432), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5616 (.Q(w6432), .A1(w5705), .A2(w6723), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5617 (.Q(w6445), .A1(w5707), .A2(w6724), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5618 (.Q(w6444), .A1(w5708), .A2(w6724), .B(w6445), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5619 (.Q(w6443), .A1(w5722), .A2(w6724), .B(w6444), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5620 (.Q(w6442), .A1(w5709), .A2(w6724), .B(w6443), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5621 (.Q(w6441), .A1(w5710), .A2(w6724), .B(w6442), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5622 (.Q(w6440), .A1(w5318), .A2(w6724), .B(w6441), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5623 (.Q(w6439), .A1(w5320), .A2(w6724), .B(w6440), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5624 (.Q(w5756), .A1(w5339), .A2(w6724), .B(w6439), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5625 (.Q(w5761), .A1(w5718), .A2(w6725), .B(w6452), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5626 (.Q(w6452), .A1(w5714), .A2(w6725), .B(w6451), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5627 (.Q(w6451), .A1(w5713), .A2(w6725), .B(w6450), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5628 (.Q(w6450), .A1(w5720), .A2(w6725), .B(w6449), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5629 (.Q(w6449), .A1(w5721), .A2(w6725), .B(w6448), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5630 (.Q(w6448), .A1(w5723), .A2(w6725), .B(w6447), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5631 (.Q(w6447), .A1(w5735), .A2(w6725), .B(w6446), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon21_sr g5632 (.Q(w6446), .A1(w5736), .A2(w6725), .B(1'b0), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_or4 g5633 (.Z(w5744), .B(w5741), .A(w5301), .C(w5709), .D(w5721) );
	vdp_or4 g5634 (.Z(w5383), .B(w5712), .A(w5379), .C(w5710), .D(w5720) );
	vdp_aon22 g5635 (.Z(w5731), .B2(w4506), .B1(w5738), .A1(w5766), .A2(DB[0]) );
	vdp_aon22 g5636 (.Z(w5730), .B2(w4507), .B1(w5738), .A1(w5766), .A2(DB[1]) );
	vdp_aon22 g5637 (.Z(w5729), .B2(w4515), .B1(w5738), .A1(w5766), .A2(DB[2]) );
	vdp_aon22 g5638 (.Z(w5728), .B2(w4506), .B1(w5738), .A1(w5766), .A2(DB[8]) );
	vdp_aon22 g5639 (.Z(w5727), .B2(w4507), .B1(w5738), .A1(w5766), .A2(DB[9]) );
	vdp_aon22 g5640 (.Z(w5726), .B2(w4515), .B1(w5738), .A1(w5766), .A2(DB[10]) );
	vdp_or4 g5641 (.Z(w5753), .B(w5701), .A(w5702), .C(w5706), .D(w5740) );
	vdp_or4 g5642 (.Z(w5745), .B(w5715), .A(w5743), .C(w5716), .D(w5742) );
	vdp_or4 g5643 (.Z(w5760), .B(w5704), .A(w5303), .C(w5708), .D(w5735) );
	vdp_or4 g5644 (.Z(w5757), .B(w5722), .A(w5723), .C(w5703), .D(w5302) );
	vdp_or4 g5645 (.Z(w5767), .B(w5717), .A(w5719), .C(w5725), .D(w5724) );
	vdp_or4 g5646 (.Z(w5758), .B(w5733), .A(w5734), .C(w5737), .D(w5732) );
	vdp_or4 g5647 (.Z(w5769), .B(w5705), .A(w5304), .C(w5707), .D(w5736) );
	vdp_comp_we g5648 (.nZ(w5738), .A(w4505), .Z(w5766) );
	vdp_not g5649 (.nZ(w6723), .A(w5364) );
	vdp_not g5650 (.nZ(w6724), .A(w5364) );
	vdp_not g5651 (.nZ(w6725), .A(w5364) );
	vdp_slatch g5652 (.Q(w5742), .D(w5784), .nC(w5750), .C(w5783) );
	vdp_comp_str g5653 (.nZ(w5750), .A(w5395), .Z(w5783) );
	vdp_slatch g5654 (.Q(w5716), .D(w5786), .nC(w5750), .C(w5783) );
	vdp_slatch g5655 (.Q(w5715), .D(w5787), .nC(w5750), .C(w5783) );
	vdp_slatch g5656 (.Q(w5743), .D(w5788), .nC(w5750), .C(w5783) );
	vdp_slatch g5657 (.Q(w5702), .D(w5789), .nC(w5750), .C(w5783) );
	vdp_slatch g5658 (.Q(w5701), .D(w5791), .nC(w5750), .C(w5783) );
	vdp_slatch g5659 (.Q(w5706), .D(w5792), .nC(w5750), .C(w5783) );
	vdp_slatch g5660 (.Q(w5740), .D(w5793), .nC(w5750), .C(w5783) );
	vdp_slatch g5661 (.Q(w5732), .D(w5802), .nC(w5764), .C(w5801) );
	vdp_comp_str g5662 (.nZ(w5764), .A(w5395), .Z(w5801) );
	vdp_slatch g5663 (.Q(w5737), .D(w5804), .nC(w5764), .C(w5801) );
	vdp_slatch g5664 (.Q(w5733), .D(w5805), .nC(w5764), .C(w5801) );
	vdp_slatch g5665 (.Q(w5734), .D(w5806), .nC(w5764), .C(w5801) );
	vdp_slatch g5666 (.Q(w5719), .D(w5807), .nC(w5764), .C(w5801) );
	vdp_slatch g5667 (.Q(w5717), .D(w5809), .nC(w5764), .C(w5801) );
	vdp_slatch g5668 (.Q(w5725), .D(w5810), .nC(w5764), .C(w5801) );
	vdp_slatch g5669 (.Q(w5724), .D(w5811), .nC(w5764), .C(w5801) );
	vdp_comp_we g5670 (.nZ(w5747), .A(1'b0), .Z(w5381) );
	vdp_aon22 g5671 (.Z(w5813), .B2(w5747), .B1(w5768), .A1(w5767), .A2(w5381) );
	vdp_not g5672 (.nZ(w5364), .A(w4517) );
	vdp_not g5673 (.nZ(w5768), .A(w5769) );
	vdp_not g5674 (.nZ(w5759), .A(w5760) );
	vdp_not g5675 (.nZ(w5755), .A(w5757) );
	vdp_not g5676 (.nZ(w5746), .A(w5744) );
	vdp_and3 g5677 (.Z(w5773), .B(w5772), .A(w5745), .C(w5744) );
	vdp_aon22 g5678 (.Z(w5781), .B2(w5747), .B1(w5746), .A1(w5745), .A2(w5381) );
	vdp_notif0 g5679 (.A(w5748), .nZ(DB[4]), .nE(w5749) );
	vdp_aon2222 g5680 (.Z(w5748), .B2(w5741), .B1(w5779), .A1(w5780), .A2(w5704), .D2(w5711), .D1(w5777), .C1(w5778), .C2(w5317) );
	vdp_notif0 g5681 (.A(w5751), .nZ(DB[12]), .nE(w5749) );
	vdp_aon2222 g5682 (.Z(w5751), .B2(w5703), .B1(w5779), .A1(w5780), .A2(w5705), .D2(w5319), .D1(w5777), .C1(w5778), .C2(w5712) );
	vdp_notif0 g5683 (.A(w6429), .nZ(DB[13]), .nE(w5749) );
	vdp_aon2222 g5684 (.Z(w6429), .B2(w5722), .B1(w5779), .A1(w5780), .A2(w5707), .D2(w5320), .D1(w5777), .C1(w5778), .C2(w5710) );
	vdp_notif0 g5685 (.A(w5754), .nZ(DB[5]), .nE(w5749) );
	vdp_aon2222 g5686 (.Z(w5754), .B2(w5709), .B1(w5779), .A1(w5780), .A2(w5708), .D2(w5339), .D1(w5777), .C1(w5778), .C2(w5318) );
	vdp_notif0 g5687 (.A(w5763), .nZ(DB[14]), .nE(w5749) );
	vdp_aon2222 g5688 (.Z(w5763), .B2(w5723), .B1(w5779), .A1(w5780), .A2(w5736), .D2(w5714), .D1(w5777), .C1(w5778), .C2(w5720) );
	vdp_notif0 g5689 (.A(w5762), .nZ(DB[6]), .nE(w5749) );
	vdp_aon2222 g5690 (.Z(w5762), .B2(w5721), .B1(w5779), .A1(w5780), .A2(w5735), .D2(w5718), .D1(w5777), .C1(w5778), .C2(w5713) );
	vdp_aon22 g5691 (.Z(w5794), .B2(w5747), .B1(w5755), .A1(w5753), .A2(w5381) );
	vdp_aon22 g5692 (.Z(w5797), .B2(w5747), .B1(w5759), .A1(w5758), .A2(w5381) );
	vdp_and3 g5693 (.Z(w5775), .B(w5796), .A(w5753), .C(w5757) );
	vdp_and3 g5694 (.Z(w5776), .B(w5798), .A(w5758), .C(w5760) );
	vdp_and3 g5695 (.Z(w5774), .B(w5812), .A(w5767), .C(w5769) );
	vdp_not g5696 (.nZ(w5749), .A(w121) );
	vdp_slatch g5697 (.Q(w5807), .D(w5458), .nC(w5843), .C(w5808) );
	vdp_slatch g5698 (.Q(w5809), .D(w5461), .nC(w5843), .C(w5808) );
	vdp_slatch g5699 (.Q(w5810), .D(w5462), .nC(w5843), .C(w5808) );
	vdp_slatch g5700 (.Q(w5811), .D(w5464), .nC(w5843), .C(w5808) );
	vdp_comp_str g5701 (.nZ(w5843), .A(w5844), .Z(w5808) );
	vdp_slatch g5702 (.Q(w5802), .D(w5445), .nC(w5838), .C(w5803) );
	vdp_slatch g5703 (.Q(w5804), .D(w5449), .nC(w5838), .C(w5803) );
	vdp_slatch g5704 (.Q(w5805), .D(w5450), .nC(w5838), .C(w5803) );
	vdp_slatch g5705 (.Q(w5806), .D(w5453), .nC(w5838), .C(w5803) );
	vdp_comp_str g5706 (.nZ(w5838), .A(w5842), .Z(w5803) );
	vdp_slatch g5707 (.Q(w5789), .D(w5458), .nC(w5825), .C(w5790) );
	vdp_slatch g5708 (.Q(w5791), .D(w5461), .nC(w5825), .C(w5790) );
	vdp_slatch g5709 (.Q(w5792), .D(w5462), .nC(w5825), .C(w5790) );
	vdp_slatch g5710 (.Q(w5793), .D(w5464), .nC(w5825), .C(w5790) );
	vdp_comp_str g5711 (.nZ(w5825), .A(w6720), .Z(w5790) );
	vdp_slatch g5712 (.Q(w5784), .D(w5445), .nC(w5824), .C(w5785) );
	vdp_slatch g5713 (.Q(w5786), .D(w5449), .nC(w5824), .C(w5785) );
	vdp_slatch g5714 (.Q(w5787), .D(w5450), .nC(w5824), .C(w5785) );
	vdp_slatch g5715 (.Q(w5788), .D(w5453), .nC(w5824), .C(w5785) );
	vdp_comp_str g5716 (.nZ(w5824), .A(w5822), .Z(w5785) );
	vdp_dlatch_inv g5717 (.nQ(w6428), .D(w5817), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5718 (.Z(w5819), .B(w5436), .A(w6428) );
	vdp_sr_bit g5719 (.Q(w126), .D(w6426), .nC2(nDCLK1), .nC1(nDCLK2), .C2(DCLK1), .C1(DCLK2) );
	vdp_sr_bit g5720 (.Q(w5816), .D(w5752), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5721 (.nQ(w5821), .D(w5782), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5722 (.nQ(w6421), .D(w5795), .nC(nDCLK2), .C(DCLK2) );
	vdp_dlatch_inv g5723 (.nQ(w6423), .D(w5831), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5724 (.Z(w6422), .B(w6423), .A(w5436) );
	vdp_sr_bit g5725 (.Q(w6431), .D(w5756), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5726 (.nQ(w5799), .D(w6718), .nC(nDCLK1), .C(DCLK1) );
	vdp_xor g5727 (.Z(w6424), .B(w5799), .A(w5436) );
	vdp_sr_bit g5728 (.Q(w5835), .D(w5761), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5729 (.nQ(w5832), .D(w6427), .nC(nDCLK2), .C(DCLK2) );
	vdp_not g5730 (.nZ(w5848), .A(w5436) );
	vdp_not g5731 (.nZ(w5800), .A(w83) );
	vdp_not g5732 (.nZ(w5836), .A(w82) );
	vdp_dlatch_inv g5733 (.nQ(w5846), .D(w6425), .nC(nDCLK2), .C(DCLK2) );
	vdp_and g5734 (.Z(w5812), .B(w5848), .A(w5437) );
	vdp_aoi21 g5735 (.Z(w6425), .B(w5833), .A1(w5813), .A2(w5812) );
	vdp_and g5736 (.Z(w5698), .B(w5846), .A(DCLK1) );
	vdp_and g5737 (.Z(w5699), .B(w5832), .A(DCLK1) );
	vdp_and g5738 (.Z(w5798), .B(w6424), .A(w5437) );
	vdp_aoi21 g5739 (.Z(w6427), .B(w5833), .A1(w5797), .A2(w5798) );
	vdp_and g5740 (.Z(w5796), .B(w6422), .A(w5437) );
	vdp_aoi21 g5741 (.Z(w5795), .B(w5820), .A1(w5794), .A2(w5796) );
	vdp_and g5742 (.Z(w5772), .B(w5437), .A(w5819) );
	vdp_aoi21 g5743 (.Z(w5782), .B(w5820), .A1(w5781), .A2(w5772) );
	vdp_and g5744 (.Z(w5739), .B(DCLK1), .A(w5821) );
	vdp_and g5745 (.Z(w5700), .B(w6421), .A(DCLK1) );
	vdp_and g5746 (.Z(w5777), .B(w5800), .A(w5836) );
	vdp_and g5747 (.Z(w5779), .B(w83), .A(w5836) );
	vdp_and g5748 (.Z(w5778), .B(w5800), .A(w82) );
	vdp_and g5749 (.Z(w5780), .B(w83), .A(w82) );
	vdp_or8 g5750 (.Z(w6426), .B(w5773), .A(w5430), .C(w5774), .D(w5814), .F(w5776), .E(w5771), .G(w5414), .H(w5775) );
	vdp_sr_bit g5751 (.Q(w5493), .D(w5854), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5752 (.Q(w5818), .D(w5493), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5753 (.Q(w5492), .D(w5830), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5754 (.Q(w5849), .D(w5492), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5755 (.Q(w5512), .D(w6411), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5756 (.Q(w5837), .D(w5512), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_comp_we g5757 (.nZ(w5852), .A(M5), .Z(w5851) );
	vdp_not g5758 (.nZ(w5844), .A(w5845) );
	vdp_or g5759 (.Z(w5516), .B(w5847), .A(w5456) );
	vdp_and3 g5760 (.Z(w5847), .B(w5508), .A(w5515), .C(w5507) );
	vdp_and3 g5761 (.Z(w5840), .B(w5508), .A(w5515), .C(w5519) );
	vdp_and3 g5762 (.Z(w6718), .B(w5513), .A(w5501), .C(w5514) );
	vdp_and3 g5763 (.Z(w5827), .B(w5520), .A(w5515), .C(w5507) );
	vdp_and3 g5764 (.Z(w5829), .B(w5520), .A(w5515), .C(w5519) );
	vdp_aoi21 g5765 (.Z(w5817), .B(w5446), .A1(w5435), .A2(w5518) );
	vdp_aon22 g5766 (.Z(w5854), .B2(w5752), .B1(w5852), .A1(w5851), .A2(w5816) );
	vdp_aon22 g5767 (.Z(w5830), .B2(w5756), .B1(w5852), .A1(w5851), .A2(w6431) );
	vdp_aon22 g5768 (.Z(w6411), .B2(w5761), .B1(w5852), .A1(w5851), .A2(w5835) );
	vdp_bufif0 g5769 (.A(w5849), .Z(COL[2]), .nE(w5853) );
	vdp_oai21 g5770 (.Z(w5828), .B(DCLK2), .A1(w5841), .A2(w5829) );
	vdp_and g5771 (.Z(w5831), .B(w5513), .A(w5501) );
	vdp_or g5772 (.Z(w5841), .B(w5827), .A(w5456) );
	vdp_bufif0 g5773 (.A(w5837), .Z(COL[3]), .nE(w5853) );
	vdp_oai21 g5774 (.Z(w5839), .B(DCLK2), .A1(w5841), .A2(w5840) );
	vdp_oai21 g5775 (.Z(w5845), .B(DCLK2), .A1(w5840), .A2(w5516) );
	vdp_not g5776 (.nZ(w5519), .A(w5507) );
	vdp_not g5777 (.nZ(w5842), .A(w5839) );
	vdp_not g5778 (.nZ(w5517), .A(w82) );
	vdp_not g5779 (.nZ(w5520), .A(w5508) );
	vdp_not g5780 (.nZ(w6720), .A(w5828) );
	vdp_not g5781 (.nZ(w5518), .A(w5514) );
	vdp_not g5782 (.nZ(w5822), .A(w5823) );
	vdp_bufif0 g5783 (.A(w5818), .Z(COL[1]), .nE(w5853) );
	vdp_oai21 g5784 (.Z(w5823), .B(DCLK2), .A1(w5499), .A2(w5829) );
	vdp_not g5785 (.nZ(w5853), .A(SPR_PRIO) );
	vdp_nand3 g5786 (.Z(w5826), .B(w120), .A(w83), .C(w5517) );
	vdp_nand g5787 (.Z(w5820), .B(w5511), .A(w5826) );
	vdp_nand3 g5788 (.Z(w5834), .B(w120), .A(w83), .C(w82) );
	vdp_nand g5789 (.Z(w5833), .B(w5511), .A(w5834) );
	vdp_sr_bit g5790 (.Q(w5881), .D(w5922), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5791 (.Q(w5882), .D(w5920), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5792 (.Q(w5879), .D(w5927), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5793 (.Q(w5880), .D(w5919), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5794 (.Z(w4512), .B2(w5881), .B1(w5916), .A1(w5915), .A2(w81), .C1(w5870), .C2(w5882) );
	vdp_aon222 g5795 (.Z(w4511), .B2(w5879), .B1(w5916), .A1(w5915), .A2(w80), .C1(w5870), .C2(w5880) );
	vdp_sr_bit g5796 (.Q(w5877), .D(w5926), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5797 (.Q(w5878), .D(w5918), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5798 (.Z(w4510), .B2(w5877), .B1(w5916), .A1(w5915), .A2(w79), .C1(w5870), .C2(w5878) );
	vdp_sr_bit g5799 (.Q(w5875), .D(w5925), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5800 (.Q(w5876), .D(w5917), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5801 (.Z(w4509), .B2(w5875), .B1(w5916), .A1(w5915), .A2(w78), .C1(w5870), .C2(w5876) );
	vdp_sr_bit g5802 (.Q(w5871), .D(w5924), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5803 (.Q(w5874), .D(w5928), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5804 (.Z(w4508), .B2(w5871), .B1(w5916), .A1(w5915), .A2(w77), .C1(w5870), .C2(w5874) );
	vdp_sr_bit g5805 (.Q(w5872), .D(w5923), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5806 (.Q(w5873), .D(w5914), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_aon222 g5807 (.Z(w4513), .B2(w5872), .B1(w5916), .A1(w5915), .A2(w76), .C1(w5870), .C2(w5873) );
	vdp_sr_bit g5808 (.Q(w5501), .D(w6697), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_slatch g5809 (.Q(w6697), .D(w5595), .nC(w5906), .C(w5867) );
	vdp_sr_bit g5810 (.Q(w5513), .D(w6695), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_slatch g5811 (.Q(w6695), .D(w5573), .nC(w5906), .C(w5867) );
	vdp_sr_bit g5812 (.Q(w5514), .D(w6696), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_slatch g5813 (.Q(w6696), .D(w5582), .nC(w5906), .C(w5867) );
	vdp_sr_bit g5814 (.Q(w5883), .D(w26), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5815 (.Q(w5866), .D(w5883), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5816 (.Q(w5865), .D(w5911), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5817 (.Q(w5899), .D(w5909), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5818 (.Q(w5898), .D(w5908), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5819 (.Q(w5862), .D(w4517), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5820 (.Q(w5861), .D(w5894), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5821 (.Q(w5889), .D(w6455), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5822 (.Q(w6455), .D(w5930), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_xor g5823 (.Z(w5891), .B(w5889), .A(w5890) );
	vdp_dlatch_inv g5824 (.nQ(w5860), .D(w5894), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5825 (.nQ(w5892), .D(w5891), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5826 (.nQ(w5863), .D(w5864), .nC(nDCLK1), .C(DCLK1) );
	vdp_dlatch_inv g5827 (.nQ(w5897), .D(w5896), .nC(nHCLK1), .C(HCLK1) );
	vdp_comp_str g5828 (.nZ(w5906), .A(w5903), .Z(w5867) );
	vdp_oai21 g5829 (.Z(w6454), .B(w5893), .A1(w5930), .A2(w5889) );
	vdp_and g5830 (.Z(w4506), .B(w5887), .A(w5859) );
	vdp_not g5831 (.nZ(w5436), .A(w5892) );
	vdp_not g5832 (.nZ(w5894), .A(w6454) );
	vdp_and g5833 (.Z(w4507), .B(w5886), .A(w5859) );
	vdp_and g5834 (.Z(w4515), .B(w5885), .A(w5859) );
	vdp_or g5835 (.Z(w5895), .B(w5861), .A(w5894) );
	vdp_not g5836 (.nZ(w5913), .A(w4505) );
	vdp_not g5837 (.nZ(w4517), .A(w5896) );
	vdp_not g5838 (.nZ(w5929), .A(M5) );
	vdp_not g5839 (.nZ(w5916), .A(w6688) );
	vdp_not g5840 (.nZ(w5868), .A(w5867) );
	vdp_not g5841 (.nZ(w5915), .A(w5913) );
	vdp_not g5842 (.nZ(w5870), .A(w5869) );
	vdp_or4 g5843 (.Z(w4514), .B(w4517), .A(w4505), .C(w5862), .D(w5895) );
	vdp_or4 g5844 (.Z(w5896), .B(w5899), .A(w5859), .C(w5865), .D(w5898) );
	vdp_nand g5845 (.Z(w5864), .B(w5897), .A(HCLK2) );
	vdp_nand g5846 (.Z(w5511), .B(w5913), .A(w5863) );
	vdp_nor g5847 (.Z(w5437), .B(w5860), .A(w4505) );
	vdp_nand g5848 (.Z(w5869), .B(w5913), .A(w5868) );
	vdp_nand g5849 (.Z(w6688), .B(w5913), .A(w5859) );
	vdp_aoi22 g5850 (.Z(w5859), .B2(w5929), .B1(w26), .A1(M5), .A2(w5866) );
	vdp_cnt_bit_load g5851 (.Q(w5959), .D(w5907), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w7), .CI(w6021), .L(w5905), .nL(w5952) );
	vdp_cnt_bit_load g5852 (.Q(w5904), .D(w5956), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w7), .CI(w5900), .L(w5905), .nL(w5952), .CO(w6021) );
	vdp_sr_bit g5853 (.Q(w5893), .D(w6418), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5854 (.SUM(w5911), .CO(w6676), .CI(1'b1), .A(HPOS[0]), .B(M5) );
	vdp_fa g5855 (.SUM(w5909), .CO(w6677), .CI(w6676), .A(HPOS[1]), .B(1'b0) );
	vdp_fa g5856 (.SUM(w5908), .CO(w6678), .CI(w6677), .A(HPOS[2]), .B(1'b1) );
	vdp_fa g5857 (.SUM(w5914), .CO(w6679), .CI(w6678), .A(w5964), .B(M5) );
	vdp_fa g5858 (.SUM(w5928), .CO(w6680), .CI(w6679), .A(HPOS[4]), .B(w5968) );
	vdp_fa g5859 (.SUM(w5917), .CO(w6681), .CI(w6680), .A(HPOS[5]), .B(1'b1) );
	vdp_fa g5860 (.SUM(w5918), .CO(w6682), .CI(w6681), .A(HPOS[6]), .B(1'b1) );
	vdp_fa g5861 (.SUM(w5919), .CO(w6683), .CI(w6682), .A(HPOS[7]), .B(1'b1) );
	vdp_fa g5862 (.SUM(w5920), .CI(w6683), .A(HPOS[8]), .B(1'b1) );
	vdp_not g5863 (.nZ(w5968), .A(M5) );
	vdp_aoi33 g5864 (.Z(w6418), .B2(w6694), .B1(w5922), .A1(H40), .A2(w5922), .A3(w5921), .B3(w6694) );
	vdp_not g5865 (.nZ(w6694), .A(H40) );
	vdp_or g5866 (.Z(w5921), .B(w5926), .A(w5927) );
	vdp_and g5867 (.Z(w5902), .B(w5900), .A(w5901) );
	vdp_sr_bit g5868 (.Q(w5900), .D(w6453), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5869 (.Q(w6453), .D(w5639), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5870 (.nQ(w5949), .D(w5488), .nC(nDCLK2), .C(DCLK2) );
	vdp_slatch g5871 (.Q(w5948), .D(w5935), .nC(w5888), .C(w5939) );
	vdp_slatch g5872 (.Q(w5887), .D(w5948), .nC(w5884), .C(w5941) );
	vdp_slatch g5873 (.Q(w5942), .D(w5933), .nC(w5888), .C(w5939) );
	vdp_slatch g5874 (.Q(w5885), .D(w5942), .nC(w5884), .C(w5941) );
	vdp_slatch g5875 (.Q(w5943), .D(w5934), .nC(w5888), .C(w5939) );
	vdp_slatch g5876 (.Q(w5886), .D(w5943), .nC(w5884), .C(w5941) );
	vdp_slatch g5877 (.Q(w6456), .D(w5644), .nC(w5888), .C(w5939) );
	vdp_sr_bit g5878 (.Q(w5890), .D(w6456), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_and g5879 (.Z(w5932), .B(DCLK2), .A(w5488) );
	vdp_comp_str g5880 (.nZ(w5884), .A(w5932), .Z(w5941) );
	vdp_comp_str g5881 (.nZ(w5888), .A(w5903), .Z(w5939) );
	vdp_not g5882 (.nZ(w5930), .A(w5949) );
	vdp_comp_we g5883 (.nZ(w5952), .A(w5902), .Z(w5905) );
	vdp_and3 g5884 (.Z(w5903), .B(HCLK1), .A(w5901), .C(w5900) );
	vdp_nand g5885 (.Z(w5956), .B(w5937), .A(M5) );
	vdp_nand g5886 (.Z(w5907), .B(w5936), .A(M5) );
	vdp_nor g5887 (.Z(w5901), .B(w5959), .A(w5904) );
	vdp_fa g5888 (.SUM(w5922), .CI(w5978), .A(w5977), .B(w5990) );
	vdp_aon22 g5889 (.Z(w5977), .B2(w5982), .B1(w5976), .A1(w6014), .A2(w5945) );
	vdp_sr_bit g5890 (.Q(w5976), .D(w5922), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5891 (.Q(w6014), .D(w6015), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5892 (.SUM(w6015), .CI(w5974), .A(w5975), .B(w6010) );
	vdp_aon22 g5893 (.Z(w5975), .B2(w5987), .B1(w6013), .A1(1'b0), .A2(w5938) );
	vdp_fa g5894 (.SUM(w5927), .CO(w5978), .CI(w5973), .A(w5972), .B(w5990) );
	vdp_aon22 g5895 (.Z(w5972), .B2(w5982), .B1(w5971), .A1(w6011), .A2(w5945) );
	vdp_sr_bit g5896 (.Q(w5971), .D(w5927), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5897 (.Q(w6011), .D(w6017), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5898 (.SUM(w6017), .CO(w5974), .CI(w5970), .A(w5969), .B(w6010) );
	vdp_aon22 g5899 (.Z(w5969), .B2(w5987), .B1(w6008), .A1(w6009), .A2(w5938) );
	vdp_fa g5900 (.SUM(w5926), .CO(w5973), .CI(w5967), .A(w5966), .B(w5990) );
	vdp_aon22 g5901 (.Z(w5966), .B2(w5982), .B1(w5965), .A1(w6007), .A2(w5945) );
	vdp_fa g5902 (.SUM(w6018), .CO(w5970), .CI(w5963), .A(w5962), .B(w5993) );
	vdp_aon22 g5903 (.Z(w5962), .B2(w5987), .B1(w6005), .A1(w6006), .A2(w5938) );
	vdp_sr_bit g5904 (.Q(w5965), .D(w5926), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5905 (.Q(w6007), .D(w6018), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5906 (.SUM(w5979), .CO(w5967), .CI(w5980), .A(w5961), .B(w5990) );
	vdp_aon22 g5907 (.Z(w5961), .B2(w5982), .B1(w5960), .A1(w6004), .A2(w5945) );
	vdp_sr_bit g5908 (.Q(w5960), .D(w5979), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5909 (.Q(w6004), .D(w6003), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5910 (.SUM(w6003), .CO(w5963), .CI(w5957), .A(w5958), .B(w5993) );
	vdp_aon22 g5911 (.Z(w5958), .B2(w5987), .B1(w6691), .A1(w6002), .A2(w5938) );
	vdp_fa g5912 (.SUM(w5924), .CO(w5980), .CI(w5954), .A(w5955), .B(w5990) );
	vdp_aon22 g5913 (.Z(w5955), .B2(w5982), .B1(w5953), .A1(w6001), .A2(w5945) );
	vdp_sr_bit g5914 (.Q(w5953), .D(w5924), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5915 (.Q(w6001), .D(w6684), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5916 (.SUM(w6684), .CO(w5957), .CI(w5951), .A(w5950), .B(w6000) );
	vdp_aon22 g5917 (.Z(w5950), .B2(w5987), .B1(w6019), .A1(w5999), .A2(w5938) );
	vdp_fa g5918 (.SUM(w5923), .CO(w5954), .CI(w5947), .A(w5946), .B(w5990) );
	vdp_aon22 g5919 (.Z(w5946), .B2(w5982), .B1(w5944), .A1(w5998), .A2(w5945) );
	vdp_sr_bit g5920 (.Q(w5944), .D(w5923), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5921 (.Q(w5998), .D(w5997), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_fa g5922 (.SUM(w5997), .CO(w5951), .CI(w5995), .A(w5940), .B(w5992) );
	vdp_aon22 g5923 (.Z(w5940), .B2(w5987), .B1(w5994), .A1(w5996), .A2(w5938) );
	vdp_aon22 g5924 (.Z(w5595), .B2(w5987), .B1(w5991), .A1(w6016), .A2(w5938) );
	vdp_aon22 g5925 (.Z(w5573), .B2(w5987), .B1(w5986), .A1(w5989), .A2(w5938) );
	vdp_aon22 g5926 (.Z(w5582), .B2(w5987), .B1(w5985), .A1(w5988), .A2(w5938) );
	vdp_and g5927 (.Z(w5947), .B(w5984), .A(w6690) );
	vdp_comp_we g5928 (.nZ(w5938), .A(M5), .Z(w5987) );
	vdp_comp_we g5929 (.nZ(w5982), .A(w6689), .Z(w5945) );
	vdp_sr_bit g5930 (.Q(w6689), .D(w5903), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5931 (.Q(w5983), .D(w5949), .nC2(nDCLK2), .nC1(nDCLK1), .C2(DCLK2), .C1(DCLK1) );
	vdp_sr_bit g5932 (.Q(w6031), .D(w6034), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5933 (.Q(w6034), .D(w6035), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5934 (.Q(w6035), .D(w6039), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5935 (.Q(w6039), .D(w6040), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5936 (.Q(w6040), .D(w6041), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5937 (.nQ(w6041), .D(w6044), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5938 (.nZ(w5991), .A(w6031) );
	vdp_sr_bit g5939 (.Q(w6045), .D(w6046), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5940 (.Q(w6046), .D(w6050), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5941 (.Q(w6050), .D(w6051), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5942 (.Q(w6051), .D(w6053), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5943 (.Q(w6053), .D(w6056), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5944 (.nQ(w6056), .D(w6055), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5945 (.nZ(w5994), .A(w6045) );
	vdp_sr_bit g5946 (.Q(w6057), .D(w6457), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5947 (.Q(w6457), .D(w6060), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5948 (.Q(w6060), .D(w6062), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5949 (.Q(w6062), .D(w6063), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5950 (.Q(w6063), .D(w6064), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5951 (.nQ(w6064), .D(w6068), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5952 (.nZ(w6019), .A(w6057) );
	vdp_sr_bit g5953 (.Q(w6069), .D(w6072), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5954 (.Q(w6072), .D(w6076), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5955 (.Q(w6076), .D(w6075), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5956 (.Q(w6075), .D(w6077), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5957 (.Q(w6077), .D(w6080), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5958 (.nQ(w6080), .D(w6081), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5959 (.nZ(w6691), .A(w6069) );
	vdp_sr_bit g5960 (.Q(w6084), .D(w6087), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5961 (.Q(w6087), .D(w6088), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5962 (.Q(w6088), .D(w6089), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5963 (.Q(w6089), .D(w6113), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5964 (.Q(w6113), .D(w6114), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5965 (.nQ(w6114), .D(w6094), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5966 (.nZ(w6005), .A(w6084) );
	vdp_sr_bit g5967 (.Q(w6115), .D(w6109), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5968 (.Q(w6109), .D(w6108), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5969 (.Q(w6108), .D(w6106), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5970 (.Q(w6106), .D(w6105), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5971 (.Q(w6105), .D(w6103), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5972 (.nQ(w6103), .D(w6093), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5973 (.nZ(w6008), .A(w6115) );
	vdp_sr_bit g5974 (.Q(w6692), .D(w6099), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5975 (.Q(w6099), .D(w6100), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5976 (.Q(w6100), .D(w6096), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5977 (.Q(w6096), .D(w6095), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5978 (.Q(w6095), .D(w6091), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5979 (.nQ(w6091), .D(w6092), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5980 (.nZ(w6013), .A(w6692) );
	vdp_and g5981 (.Z(w5990), .B(w5984), .A(w5890) );
	vdp_and g5982 (.Z(w6027), .B(w5644), .A(w5937) );
	vdp_and g5983 (.Z(w6028), .B(w5995), .A(w5936) );
	vdp_or g5984 (.Z(w5992), .B(w6027), .A(w5993) );
	vdp_and g5985 (.B(w6030), .A(M5) );
	vdp_or g5986 (.Z(w6000), .B(w6028), .A(w5993) );
	vdp_and g5987 (.Z(w5993), .B(w23), .A(w6701) );
	vdp_or g5988 (.Z(w6010), .B(w5993), .A(M5) );
	vdp_not g5989 (.nZ(w6701), .A(M5) );
	vdp_not g5990 (.nZ(w6690), .A(w5890) );
	vdp_nor g5991 (.Z(w5984), .B(w6689), .A(w5983) );
	vdp_sr_bit g5992 (.Q(w6043), .D(w6047), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5993 (.Q(w6047), .D(w6048), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5994 (.Q(w6048), .D(w6049), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5995 (.Q(w6049), .D(w6052), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g5996 (.Q(w6052), .D(w6693), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g5997 (.nQ(w6693), .D(w6122), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g5998 (.nZ(w5934), .A(w6043) );
	vdp_sr_bit g5999 (.Q(w6032), .D(w6033), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6000 (.Q(w6033), .D(w6036), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6001 (.Q(w6036), .D(w6037), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6002 (.Q(w6037), .D(w6038), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6003 (.Q(w6038), .D(w6042), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6004 (.nQ(w6042), .D(w6121), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6005 (.nZ(w5935), .A(w6032) );
	vdp_sr_bit g6006 (.Q(w6022), .D(w6023), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6007 (.Q(w6023), .D(w6024), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6008 (.Q(w6024), .D(w6026), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6009 (.Q(w6026), .D(w6025), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6010 (.Q(w6025), .D(w6029), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6011 (.nQ(w6029), .D(w6120), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6012 (.nZ(w6030), .A(w6022) );
	vdp_sr_bit g6013 (.Q(w6054), .D(w6058), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6014 (.Q(w6058), .D(w6059), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6015 (.Q(w6059), .D(w6061), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6016 (.Q(w6061), .D(w6065), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6017 (.Q(w6065), .D(w6066), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6018 (.nQ(w6066), .D(w6127), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6019 (.nZ(w5933), .A(w6054) );
	vdp_sr_bit g6020 (.Q(w6067), .D(w6070), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6021 (.Q(w6070), .D(w6071), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6022 (.Q(w6071), .D(w6073), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6023 (.Q(w6073), .D(w6074), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6024 (.Q(w6074), .D(w6078), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6025 (.nQ(w6078), .D(w6123), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6026 (.nZ(w5937), .A(w6067) );
	vdp_sr_bit g6027 (.Q(w6079), .D(w6082), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6028 (.Q(w6082), .D(w6083), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6029 (.Q(w6083), .D(w6085), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6030 (.Q(w6085), .D(w6086), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6031 (.Q(w6086), .D(w6090), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6032 (.nQ(w6090), .D(w6124), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6033 (.nZ(w5936), .A(w6079) );
	vdp_sr_bit g6034 (.Q(w6111), .D(w6112), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6035 (.Q(w6112), .D(w6116), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6036 (.Q(w6116), .D(w6117), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6037 (.Q(w6117), .D(w6110), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6038 (.Q(w6110), .D(w6107), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6039 (.nQ(w6107), .D(w6125), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6040 (.nZ(w5985), .A(w6111) );
	vdp_sr_bit g6041 (.Q(w6102), .D(w6104), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6042 (.Q(w6104), .D(w6101), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6043 (.Q(w6101), .D(w6098), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6044 (.Q(w6098), .D(w6097), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6045 (.Q(w6097), .D(w6118), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6046 (.nQ(w6118), .D(w6126), .nC(nHCLK2), .C(HCLK2) );
	vdp_not g6047 (.nZ(w5986), .A(w6102) );
	vdp_slatch g6048 (.D(w6152), .nC(w6190), .C(w6130), .nQ(w5988) );
	vdp_slatch g6049 (.D(S[1]), .nC(w6191), .C(w6134), .Q(w6151) );
	vdp_slatch g6050 (.D(S[1]), .nC(w6192), .C(w6133), .Q(w6150) );
	vdp_aoi22 g6051 (.Z(w6149), .B2(w6196), .B1(w6151), .A1(w6150), .A2(w6131) );
	vdp_slatch g6052 (.D(S[0]), .nC(w6191), .C(w6134), .Q(w6154) );
	vdp_slatch g6053 (.D(S[0]), .nC(w6192), .C(w6133), .Q(w6153) );
	vdp_aoi22 g6054 (.Z(w6152), .B2(w6196), .B1(w6154), .A1(w6153), .A2(w6131) );
	vdp_slatch g6055 (.D(w6149), .nC(w6190), .C(w6130), .nQ(w5989) );
	vdp_slatch g6056 (.D(S[2]), .nC(w6191), .C(w6134), .Q(w6148) );
	vdp_slatch g6057 (.D(S[2]), .nC(w6192), .C(w6133), .Q(w6147) );
	vdp_aoi22 g6058 (.Z(w6233), .B2(w6196), .B1(w6148), .A1(w6147), .A2(w6131) );
	vdp_slatch g6059 (.D(w6233), .nC(w6190), .C(w6130), .nQ(w6016) );
	vdp_slatch g6060 (.D(S[3]), .nC(w6191), .C(w6134), .Q(w6146) );
	vdp_slatch g6061 (.D(S[3]), .nC(w6192), .C(w6133), .Q(w6145) );
	vdp_aoi22 g6062 (.Z(w6144), .B2(w6196), .B1(w6146), .A1(w6145), .A2(w6131) );
	vdp_slatch g6063 (.D(w6144), .nC(w6190), .C(w6130), .nQ(w5996) );
	vdp_slatch g6064 (.D(S[4]), .nC(w6191), .C(w6134), .Q(w6143) );
	vdp_slatch g6065 (.D(S[4]), .nC(w6192), .C(w6133), .Q(w6142) );
	vdp_aoi22 g6066 (.Z(w6141), .B2(w6196), .B1(w6143), .A1(w6142), .A2(w6131) );
	vdp_slatch g6067 (.D(w6141), .nC(w6190), .C(w6130), .nQ(w5999) );
	vdp_slatch g6068 (.D(S[5]), .nC(w6191), .C(w6134), .Q(w6140) );
	vdp_slatch g6069 (.D(S[5]), .nC(w6192), .C(w6133), .Q(w6139) );
	vdp_aoi22 g6070 (.Z(w6138), .B2(w6196), .B1(w6140), .A1(w6139), .A2(w6131) );
	vdp_slatch g6071 (.D(w6138), .nC(w6190), .C(w6130), .nQ(w6002) );
	vdp_slatch g6072 (.D(S[6]), .nC(w6191), .C(w6134), .Q(w6137) );
	vdp_slatch g6073 (.D(S[6]), .nC(w6192), .C(w6133), .Q(w6135) );
	vdp_aoi22 g6074 (.Z(w6136), .B2(w6196), .B1(w6137), .A1(w6135), .A2(w6131) );
	vdp_slatch g6075 (.D(w6136), .nC(w6190), .C(w6130), .nQ(w6006) );
	vdp_slatch g6076 (.D(S[7]), .nC(w6191), .C(w6134), .Q(w6132) );
	vdp_slatch g6077 (.D(S[7]), .nC(w6192), .C(w6133), .Q(w6128) );
	vdp_aoi22 g6078 (.Z(w6129), .B2(w6196), .B1(w6132), .A1(w6128), .A2(w6131) );
	vdp_slatch g6079 (.D(w6129), .nC(w6190), .C(w6130), .nQ(w6009) );
	vdp_comp_str g6080 (.nZ(w6190), .A(w5639), .Z(w6130) );
	vdp_comp_str g6081 (.nZ(w6191), .A(w4969), .Z(w6134) );
	vdp_comp_str g6082 (.nZ(w6192), .A(w4973), .Z(w6133) );
	vdp_comp_we g6083 (.nZ(w6196), .A(w6189), .Z(w6131) );
	vdp_sr_bit g6084 (.Q(w6187), .D(w6183), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6085 (.Z(w6183), .B(w6188), .A(w6155) );
	vdp_fa g6086 (.SUM(w6188), .CI(w6157), .A(w6187), .B(1'b0) );
	vdp_sr_bit g6087 (.Q(w6222), .D(w6178), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6088 (.Z(w6178), .B(w6184), .A(w6155) );
	vdp_fa g6089 (.SUM(w6184), .CO(w6157), .CI(w6158), .A(w6222), .B(1'b0) );
	vdp_sr_bit g6090 (.Q(w6179), .D(w6202), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6091 (.Z(w6202), .B(w6180), .A(w6155) );
	vdp_fa g6092 (.SUM(w6180), .CO(w6158), .CI(w6160), .A(w6179), .B(w6159) );
	vdp_sr_bit g6093 (.Q(w6175), .D(w6174), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_and g6094 (.Z(w6174), .B(w6176), .A(w6155) );
	vdp_fa g6095 (.SUM(w6176), .CO(w6160), .CI(w6162), .A(w6175), .B(w6161) );
	vdp_sr_bit g6096 (.Q(w6165), .D(w6698), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6097 (.Q(w6698), .D(w22), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6098 (.nQ(w6163), .D(w6165), .nC(nHCLK1), .C(HCLK1) );
	vdp_dlatch_inv g6099 (.nQ(w6155), .D(w6164), .nC(nHCLK1), .C(HCLK1) );
	vdp_and g6100 (.Z(w6159), .B(w6162), .A(w6171) );
	vdp_and g6101 (.Z(w6161), .B(w6162), .A(w6170) );
	vdp_and g6102 (.Z(w4595), .B(w6698), .A(w6247) );
	vdp_or g6103 (.Z(w6164), .B(w6168), .A(w6234) );
	vdp_not g6104 (.nZ(w6167), .A(M5) );
	vdp_not g6105 (.nZ(w6162), .A(w6163) );
	vdp_fa g6106 (.SUM(w6207), .CO(w6210), .CI(w6208), .A(w6261), .B(w6181) );
	vdp_aoi22 g6107 (.Z(w6273), .B2(w6193), .B1(w6209), .A1(w6207), .A2(w6257) );
	vdp_notif0 g6108 (.A(w6273), .nZ(VRAMA[9]), .nE(w6250) );
	vdp_fa g6109 (.SUM(w6198), .CO(w6208), .CI(w6204), .A(w6260), .B(w6185) );
	vdp_aoi22 g6110 (.Z(w6206), .B2(w6193), .B1(w6207), .A1(w6198), .A2(w6257) );
	vdp_notif0 g6111 (.A(w6206), .nZ(VRAMA[8]), .nE(w6250) );
	vdp_fa g6112 (.SUM(w6194), .CO(w6204), .CI(w6197), .A(w6259), .B(w6177) );
	vdp_aoi22 g6113 (.Z(w6205), .B2(w6193), .B1(w6198), .A1(w6194), .A2(w6257) );
	vdp_notif0 g6114 (.A(w6205), .nZ(VRAMA[7]), .nE(w6250) );
	vdp_fa g6115 (.SUM(w6200), .CO(w6197), .CI(1'b0), .A(w6258), .B(w6173) );
	vdp_aoi22 g6116 (.Z(w6195), .B2(w6193), .B1(w6194), .A1(w6200), .A2(w6257) );
	vdp_notif0 g6117 (.A(w6195), .nZ(VRAMA[6]), .nE(w6250) );
	vdp_not g6118 (.nZ(w6250), .A(w6264) );
	vdp_ha g6119 (.SUM(w6209), .B(w6262), .A(w6210), .CO(w6211) );
	vdp_aoi22 g6120 (.Z(w6213), .B2(w6193), .B1(w6212), .A1(w6209), .A2(w6257) );
	vdp_notif0 g6121 (.A(w6213), .nZ(VRAMA[10]), .nE(w6267) );
	vdp_ha g6122 (.SUM(w6212), .B(w6263), .A(w6211), .CO(w6214) );
	vdp_aoi22 g6123 (.Z(w6215), .B2(w6193), .B1(w6223), .A1(w6212), .A2(w6257) );
	vdp_notif0 g6124 (.A(w6215), .nZ(VRAMA[11]), .nE(w6267) );
	vdp_ha g6125 (.SUM(w6223), .B(w6266), .A(w6214), .CO(w6216) );
	vdp_aoi22 g6126 (.Z(w6218), .B2(w6193), .B1(w6217), .A1(w6223), .A2(w6257) );
	vdp_notif0 g6127 (.A(w6218), .nZ(VRAMA[12]), .nE(w6267) );
	vdp_ha g6128 (.SUM(w6217), .B(w6265), .A(w6216), .CO(w6220) );
	vdp_aoi22 g6129 (.Z(w6221), .B2(w6193), .B1(w6219), .A1(w6217), .A2(w6257) );
	vdp_notif0 g6130 (.A(w6221), .nZ(VRAMA[13]), .nE(w6267) );
	vdp_ha g6131 (.SUM(w6219), .B(w6269), .A(w6220), .CO(w6226) );
	vdp_aoi22 g6132 (.Z(w6224), .B2(w6193), .B1(w6225), .A1(w6219), .A2(w6257) );
	vdp_notif0 g6133 (.A(w6224), .nZ(VRAMA[14]), .nE(w6267) );
	vdp_ha g6134 (.SUM(w6225), .B(w6268), .A(w6226), .CO(w6227) );
	vdp_aoi22 g6135 (.Z(w6230), .B2(w6193), .B1(w6231), .A1(w6225), .A2(w6257) );
	vdp_notif0 g6136 (.A(w6230), .nZ(VRAMA[15]), .nE(w6267) );
	vdp_ha g6137 (.SUM(w6231), .B(w6271), .A(w6227) );
	vdp_aoi22 g6138 (.Z(w6229), .B2(w6193), .B1(w5245), .A1(w6231), .A2(w6257) );
	vdp_notif0 g6139 (.A(w6229), .nZ(VRAMA[16]), .nE(w6267) );
	vdp_not g6140 (.nZ(w6267), .A(w6264) );
	vdp_sr_bit g6141 (.Q(w6264), .D(w6417), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_dlatch_inv g6142 (.nQ(w4516), .D(w6228), .nC(nHCLK2), .C(HCLK2) );
	vdp_and g6143 (.Z(w6417), .B(M5), .A(w22) );
	vdp_or9 g6144 (.Z(w6228), .B(w6126), .A(w6125), .C(w6044), .D(w6055), .F(w6081), .E(w6068), .G(w6094), .H(w6093), .I(w6092) );
	vdp_sr_bit g6145 (.Q(w4589), .D(w6562), .nC2(nHCLK1), .nC1(nHCLK2), .C2(HCLK1), .C1(HCLK2) );
	vdp_sr_bit g6146 (.D(w6699), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_fa g6147 (.SUM(w6173), .CO(w6685), .CI(1'b0), .A(w6245), .B(w6174) );
	vdp_fa g6148 (.SUM(w6177), .CO(w6686), .CI(w6685), .A(w6246), .B(w6202) );
	vdp_fa g6149 (.SUM(w6185), .CO(w6687), .CI(w6686), .A(1'b0), .B(w6178) );
	vdp_fa g6150 (.SUM(w6181), .CI(w6687), .A(1'b0), .B(w6183) );
	vdp_notif0 g6151 (.A(1'b1), .nZ(VRAMA[0]), .nE(w6250) );
	vdp_notif0 g6152 (.A(1'b1), .nZ(VRAMA[1]), .nE(w6250) );
	vdp_not g6153 (.nZ(w6182), .A(w6251) );
	vdp_notif0 g6154 (.A(w6182), .nZ(VRAMA[2]), .nE(w6250) );
	vdp_not g6155 (.nZ(w6186), .A(w6253) );
	vdp_notif0 g6156 (.A(w6186), .nZ(VRAMA[3]), .nE(w6250) );
	vdp_not g6157 (.nZ(w6199), .A(w6252) );
	vdp_notif0 g6158 (.A(w6199), .nZ(VRAMA[4]), .nE(w6250) );
	vdp_notif0 g6159 (.A(w6201), .nZ(VRAMA[5]), .nE(w6250) );
	vdp_aoi22 g6160 (.Z(w6201), .B2(w6193), .B1(w6200), .A1(w6243), .A2(w6257) );
	vdp_comp_we g6161 (.nZ(w6193), .A(w1), .Z(w6257) );
	vdp_aon22 g6162 (.Z(w6245), .B2(w6169), .B1(w6243), .A1(w6241), .A2(w6244) );
	vdp_aon22 g6163 (.Z(w6246), .B2(w6169), .B1(w6241), .A1(w6240), .A2(w6244) );
	vdp_comp_we g6164 (.nZ(w6169), .A(w1), .Z(w6244) );
	vdp_or g6165 (.Z(w6699), .B(w6234), .A(w4595) );
	vdp_nor g6166 (.Z(w6562), .B(w6168), .A(w6167) );
	vdp_comp_str g6167 (.nZ(w6297), .A(w6254), .Z(w6270) );
	vdp_slatch g6168 (.D(w6300), .nC(w6297), .C(w6270), .Q(w6125) );
	vdp_aon22 g6169 (.Z(w6301), .B2(w6274), .B1(w6153), .A1(DB[0]), .A2(w6255) );
	vdp_slatch g6170 (.D(w6302), .nC(w6297), .C(w6270), .Q(w6126) );
	vdp_aon22 g6171 (.Z(w6303), .B2(w6274), .B1(w6150), .A1(DB[1]), .A2(w6255) );
	vdp_slatch g6172 (.D(w6304), .nC(w6297), .C(w6270), .Q(w6044) );
	vdp_aon22 g6173 (.Z(w6305), .B2(w6274), .B1(w6147), .A1(DB[2]), .A2(w6255) );
	vdp_slatch g6174 (.D(w6306), .nC(w6297), .C(w6270), .Q(w6055) );
	vdp_aon22 g6175 (.Z(w6307), .B2(w6274), .B1(w6145), .A1(DB[3]), .A2(w6255) );
	vdp_slatch g6176 (.D(w6308), .nC(w6297), .C(w6270), .Q(w6068) );
	vdp_aon22 g6177 (.Z(w6309), .B2(w6274), .B1(w6142), .A1(DB[4]), .A2(w6255) );
	vdp_slatch g6178 (.D(w6310), .nC(w6297), .C(w6270), .Q(w6081) );
	vdp_aon22 g6179 (.Z(w6311), .B2(w6274), .B1(w6139), .A1(DB[5]), .A2(w6255) );
	vdp_slatch g6180 (.D(w6312), .nC(w6297), .C(w6270), .Q(w6094) );
	vdp_aon22 g6181 (.Z(w6313), .B2(w6274), .B1(w6135), .A1(DB[6]), .A2(w6255) );
	vdp_slatch g6182 (.D(w6315), .nC(w6297), .C(w6270), .Q(w6093) );
	vdp_aon22 g6183 (.Z(w6316), .B2(w6274), .B1(w6128), .A1(DB[7]), .A2(w6255) );
	vdp_slatch g6184 (.D(w6314), .nC(w6297), .C(w6270), .Q(w6092) );
	vdp_aon22 g6185 (.Z(w6317), .B2(w6274), .B1(w5084), .A1(DB[8]), .A2(w6255) );
	vdp_slatch g6186 (.D(w6288), .nC(w6285), .C(w6256), .Q(w6260) );
	vdp_aon22 g6187 (.Z(w6324), .B2(w6274), .B1(w6148), .A1(DB[2]), .A2(w6255) );
	vdp_slatch g6188 (.D(w6287), .nC(w6285), .C(w6256), .Q(w6261) );
	vdp_aon22 g6189 (.Z(w6319), .B2(w6274), .B1(w6146), .A1(DB[3]), .A2(w6255) );
	vdp_slatch g6190 (.D(w6294), .nC(w6285), .C(w6256), .Q(w6262) );
	vdp_aon22 g6191 (.Z(w6320), .B2(w6274), .B1(w6143), .A1(DB[4]), .A2(w6255) );
	vdp_slatch g6192 (.D(w6293), .nC(w6285), .C(w6256), .Q(w6263) );
	vdp_aon22 g6193 (.Z(w6323), .B2(w6274), .B1(w6140), .A1(DB[5]), .A2(w6255) );
	vdp_slatch g6194 (.D(w6291), .nC(w6285), .C(w6256), .Q(w6266) );
	vdp_aon22 g6195 (.Z(w6325), .B2(w6274), .B1(w6137), .A1(DB[6]), .A2(w6255) );
	vdp_slatch g6196 (.D(w6292), .nC(w6285), .C(w6256), .Q(w6265) );
	vdp_aon22 g6197 (.Z(w6326), .B2(w6274), .B1(w6132), .A1(DB[7]), .A2(w6255) );
	vdp_slatch g6198 (.D(w6290), .nC(w6285), .C(w6256), .Q(w6269) );
	vdp_aon22 g6199 (.Z(w6327), .B2(w6274), .B1(w5024), .A1(DB[8]), .A2(w6255) );
	vdp_slatch g6200 (.D(w6283), .nC(w6285), .C(w6256), .Q(w6268) );
	vdp_aon22 g6201 (.Z(w6282), .B2(w6274), .B1(w5085), .A1(DB[9]), .A2(w6255) );
	vdp_slatch g6202 (.D(w6298), .nC(w6285), .C(w6256), .Q(w6271) );
	vdp_aon22 g6203 (.Z(w6299), .B2(w6274), .B1(w5093), .A1(DB[10]), .A2(w6255) );
	vdp_slatch g6204 (.D(w6286), .nC(w6285), .C(w6256), .Q(w6258) );
	vdp_aon22 g6205 (.Z(w6321), .B2(w6274), .B1(w6154), .A1(DB[0]), .A2(w6255) );
	vdp_slatch g6206 (.D(w6329), .nC(w6285), .C(w6256), .Q(w6259) );
	vdp_aon22 g6207 (.Z(w6322), .B2(w6274), .B1(w6151), .A1(DB[1]), .A2(w6255) );
	vdp_comp_str g6208 (.nZ(w6285), .A(w6254), .Z(w6256) );
	vdp_not g6209 (.nZ(w6254), .A(w6412) );
	vdp_oai21 g6210 (.Z(w6412), .B(HCLK1), .A1(w6168), .A2(w122) );
	vdp_sr_bit g6211 (.Q(w6413), .D(w6415), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6212 (.Q(w5639), .D(w6414), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6213 (.Q(w6189), .D(w6416), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6214 (.Q(w6318), .D(w5598), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_cnt_bit_load g6215 (.Q(w6237), .D(w6242), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w6234), .CI(w22), .L(w6239), .nL(w6277), .CO(w6278) );
	vdp_cnt_bit_load g6216 (.Q(w6276), .D(w6238), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w6234), .CI(w6278), .L(w6239), .nL(w6277) );
	vdp_comp_we g6217 (.nZ(w6277), .A(w6168), .Z(w6239) );
	vdp_not g6218 (.nZ(w6242), .A(w6279) );
	vdp_not g6219 (.nZ(w6238), .A(w6275) );
	vdp_not g6220 (.nZ(w6235), .A(w125) );
	vdp_nand g6221 (.Z(w6330), .B(w125), .A(w4589) );
	vdp_nand g6222 (.Z(w6236), .B(w6235), .A(w4589) );
	vdp_not g6223 (.nZ(w6274), .A(w6236) );
	vdp_nor g6224 (.Z(w6247), .B(w6276), .A(w6237) );
	vdp_and g6225 (.Z(w6168), .B(w6247), .A(w22) );
	vdp_rs_FF g6226 (.Q(w6415), .R(w6248), .S(w6234) );
	vdp_and3 g6227 (.Z(w6414), .B(w5598), .A(w4596), .C(w6413) );
	vdp_cnt_bit g6228 (.Q(w6416), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1), .R(w7), .CI(w6318) );
	vdp_not g6229 (.nZ(w6255), .A(w6330) );
	vdp_not g6230 (.nZ(w6281), .A(w4551) );
	vdp_not g6231 (.nZ(w6284), .A(w4552) );
	vdp_comp_str g6232 (.nZ(w6280), .A(w6254), .Z(w6332) );
	vdp_not g6233 (.nZ(w6340), .A(w122) );
	vdp_aon22 g6234 (.Z(w6342), .B2(w6274), .B1(w5145), .A1(DB[0]), .A2(w6255) );
	vdp_slatch g6235 (.D(w6331), .nC(w6280), .C(w6332), .Q(w6120) );
	vdp_bufif0 g6236 (.A(w6339), .Z(DB[0]), .nE(w6340) );
	vdp_aon222 g6237 (.Z(w6339), .B2(w4553), .B1(w6125), .A1(w6120), .A2(w6281), .C1(w6258), .C2(w6284) );
	vdp_aon22 g6238 (.Z(w6345), .B2(w6274), .B1(w5226), .A1(DB[1]), .A2(w6255) );
	vdp_slatch g6239 (.D(w6341), .nC(w6280), .C(w6332), .Q(w6121) );
	vdp_bufif0 g6240 (.A(w6343), .Z(DB[1]), .nE(w6340) );
	vdp_aon222 g6241 (.Z(w6343), .B2(w4553), .B1(w6126), .A1(w6121), .A2(w6281), .C1(w6259), .C2(w6284) );
	vdp_aon22 g6242 (.Z(w6347), .B2(w6274), .B1(w5246), .A1(DB[2]), .A2(w6255) );
	vdp_slatch g6243 (.D(w6344), .nC(w6280), .C(w6332), .Q(w6122) );
	vdp_bufif0 g6244 (.A(w6346), .Z(DB[2]), .nE(w6340) );
	vdp_aon222 g6245 (.Z(w6346), .B2(w4553), .B1(w6044), .A1(w6122), .A2(w6281), .C1(w6260), .C2(w6284) );
	vdp_aon22 g6246 (.Z(w6356), .B2(w6274), .B1(w5211), .A1(DB[3]), .A2(w6255) );
	vdp_slatch g6247 (.D(w6348), .nC(w6280), .C(w6332), .Q(w6127) );
	vdp_bufif0 g6248 (.A(w6355), .Z(DB[3]), .nE(w6340) );
	vdp_aon222 g6249 (.Z(w6355), .B2(w4553), .B1(w6055), .A1(w6127), .A2(w6281), .C1(w6261), .C2(w6284) );
	vdp_aon22 g6250 (.Z(w6353), .B2(w6274), .B1(w4533), .A1(DB[4]), .A2(w6255) );
	vdp_slatch g6251 (.D(w6279), .nC(w6280), .C(w6332), .Q(w6123) );
	vdp_bufif0 g6252 (.A(w6354), .Z(DB[4]), .nE(w6340) );
	vdp_aon222 g6253 (.Z(w6354), .B2(w4553), .B1(w6068), .A1(w6123), .A2(w6281), .C1(w6262), .C2(w6284) );
	vdp_aon22 g6254 (.Z(w6351), .B2(w6274), .B1(w4579), .A1(DB[5]), .A2(w6255) );
	vdp_slatch g6255 (.D(w6275), .nC(w6280), .C(w6332), .Q(w6124) );
	vdp_bufif0 g6256 (.A(w6352), .Z(DB[5]), .nE(w6340) );
	vdp_aon222 g6257 (.Z(w6352), .B2(w4553), .B1(w6081), .A1(w6124), .A2(w6281), .C1(w6263), .C2(w6284) );
	vdp_aon22 g6258 (.Z(w6349), .B2(w6274), .B1(w4534), .A1(DB[6]), .A2(w6255) );
	vdp_slatch g6259 (.D(w6350), .nC(w6280), .C(w6332), .Q(w6170) );
	vdp_bufif0 g6260 (.A(w6372), .Z(DB[6]), .nE(w6340) );
	vdp_aon222 g6261 (.Z(w6372), .B2(w4553), .B1(w6094), .A1(w6170), .A2(w6281), .C1(w6266), .C2(w6284) );
	vdp_aon22 g6262 (.Z(w6368), .B2(w6274), .B1(w4529), .A1(DB[7]), .A2(w6255) );
	vdp_slatch g6263 (.D(w6369), .nC(w6289), .C(w6370), .Q(w6171) );
	vdp_bufif0 g6264 (.A(w6371), .Z(DB[7]), .nE(w6340) );
	vdp_aon222 g6265 (.Z(w6371), .B2(w4553), .B1(w6093), .A1(w6171), .A2(w6281), .C1(w6265), .C2(w6284) );
	vdp_aon22 g6266 (.Z(w6366), .B2(w6274), .B1(w6333), .A1(DB[8]), .A2(w6255) );
	vdp_slatch g6267 (.D(w6367), .nC(w6289), .C(w6370), .Q(w6251) );
	vdp_bufif0 g6268 (.A(w6700), .Z(DB[8]), .nE(w6340) );
	vdp_aon222 g6269 (.Z(w6700), .B2(w4553), .B1(w6092), .A1(w6251), .A2(w6281), .C1(w6269), .C2(w6284) );
	vdp_aon22 g6270 (.Z(w6364), .B2(w6274), .B1(w6338), .A1(DB[9]), .A2(w6255) );
	vdp_slatch g6271 (.D(w6365), .nC(w6289), .C(w6370), .Q(w6253) );
	vdp_bufif0 g6272 (.A(w6373), .Z(DB[9]), .nE(w6340) );
	vdp_aon222 g6273 (.Z(w6373), .B2(w4553), .B1(1'b0), .A1(w6253), .A2(w6281), .C1(w6268), .C2(w6284) );
	vdp_aon22 g6274 (.Z(w6362), .B2(w6274), .B1(w6337), .A1(DB[10]), .A2(w6255) );
	vdp_slatch g6275 (.D(w6363), .nC(w6289), .C(w6370), .Q(w6252) );
	vdp_bufif0 g6276 (.A(w6374), .Z(DB[10]), .nE(w6340) );
	vdp_aon222 g6277 (.Z(w6374), .B2(w4553), .B1(1'b0), .A1(w6252), .A2(w6281), .C1(w6271), .C2(w6284) );
	vdp_aon22 g6278 (.Z(w6360), .B2(w6274), .B1(w6336), .A1(DB[11]), .A2(w6255) );
	vdp_slatch g6279 (.D(w6361), .nC(w6289), .C(w6370), .Q(w6243) );
	vdp_bufif0 g6280 (.A(w6243), .Z(DB[11]), .nE(w6340) );
	vdp_aon22 g6281 (.Z(w6359), .B2(w6274), .B1(w6335), .A1(DB[12]), .A2(w6255) );
	vdp_slatch g6282 (.D(w6375), .nC(w6289), .C(w6370), .Q(w6241) );
	vdp_bufif0 g6283 (.A(w6241), .Z(DB[12]), .nE(w6340) );
	vdp_aon22 g6284 (.Z(w6357), .B2(w6274), .B1(w6334), .A1(DB[13]), .A2(w6255) );
	vdp_slatch g6285 (.D(w6358), .nC(w6289), .C(w6370), .Q(w6240) );
	vdp_bufif0 g6286 (.A(w6240), .Z(DB[13]), .nE(w6340) );
	vdp_comp_str g6287 (.nZ(w6289), .A(w6254), .Z(w6370) );
	vdp_sr_bit g6288 (.Q(w4698), .D(w131), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6289 (.Q(w4699), .D(VRAMA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6290 (.Q(w6383), .D(w6377), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6291 (.Q(w4691), .D(VRAMA[3]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6292 (.Q(w4693), .D(VRAMA[4]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6293 (.Q(w4694), .D(VRAMA[5]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6294 (.Q(w4695), .D(VRAMA[6]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6295 (.Q(w4696), .D(VRAMA[7]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6296 (.Q(w4697), .D(VRAMA[8]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6297 (.Q(w4638), .D(w6381), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6298 (.Q(w4637), .D(w6382), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_and g6299 (.Z(w6381), .B(w134), .A(w5210) );
	vdp_and g6300 (.Z(w6382), .B(w133), .A(w5210) );
	vdp_sr_bit g6301 (.Q(w6396), .D(RD_DATA[0]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6302 (.Q(w6397), .D(RD_DATA[1]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6303 (.Q(w6399), .D(w324), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_sr_bit g6304 (.Q(w6398), .D(RD_DATA[2]), .nC2(nHCLK2), .nC1(nHCLK1), .C2(HCLK2), .C1(HCLK1) );
	vdp_V_PLA g6305 (.o[0](w1886), .o[1](w1887), .o[2](w1888), .o[3](w1889), .o[4](w1890), .o[5](w1891), .o[6](w1892), .o[7](w1893), .o[8](w1894), .o[9](w1895), .o[10](w1896), .o[11](w1897), .o[12](w1898), .o[13](w1899), .o[14](w1900), .o[15](w6818), .o[16](w6819), .o[17](w6820), .o[18](w1901), .o[19](w1902), .o[20](w1903), .o[21](w1904), .o[22](w6821), .o[23](w1905), .o[24](w1980), .o[25](w1906), .o[26](w1907), .o[27](w1981), .o[28](w1995), .o[29](w1994), .o[30](w2014), .o[31](w1923), .o[32](w1885), .o[33](w1884), .o[34](w1924), .o[35](w1908), .o[36](w1925), .o[37](w1926), .o[38](w1883), .o[39](w1882), .o[40](w1929), .o[41](w1927), .o[42](w1928), .o[43](w1880), .o[44](w1879), .o[45](w1878), .o[46](w1877), .o[47](w6707), .Vcnt[0](w1702), .Vcnt[1](w1845), .Vcnt[2](w1937), .Vcnt[3](w1830), .Vcnt[4](w1936), .Vcnt[5](w1785), .Vcnt[6](w1748), .Vcnt[7](w1819), .Vcnt[8](w1846), .ODD_EVEN(ODD/EVEN), .LS0(LS0), .PAL(PAL), .nPAL(w1838), .2(w1837), .3(w1826), .M5(M5) );
	vdp_not g6306 (.A(w592), .nZ(w6705) );
	vdp_not g6307 (.A(w966), .nZ(w6706) );
	vdp_not g6308 (.nZ(w2451), .A(w6705) );
	vdp_not g6309 (.nZ(w2452), .A(w6706) );
	vdp_cram g6310 (.q[8](w2750), .D[8](w2751), .q[7](w2852), .D[7](w2752), .q[6](w2749), .D[6](w2753), .q[5](w2755), .D[5](w2754), .q[4](w2748), .D[4](w2756), .q[3](w2757), .D[3](w2981), .q[2](w2747), .D[2](w2758), .q[1](w2746), .D[1](w2759), .q[0](w2744), .D[0](w2760), .A[0](w2780), .A[1](w2784), .CLK(HCLK1), .A[2](w2790), .A[3](w2799), .A[4](w2820), .A[5](w2819), .B(w2826), .A(w2825) );
	vdp_linebuf_ram g6311 (.q[0](w5335), .D[0](w5731), .q[1](w5324), .D[1](w5730), .q[2](w5312), .D[2](w5729), .q[3](w5301), .D[3](w5742), .q[4](w5741), .D[4](w5716), .q[5](w5709), .D[5](w5715), .q[6](w5721), .D[6](w5743), .q[7](w5334), .D[7](w5728), .q[8](w5325), .D[8](w5727), .q[9](w5311), .D[9](w5726), .q[10](w5302), .D[10](w5702), .q[11](w5703), .D[11](w5701), .q[12](w5722), .D[12](w5706), .q[13](w5723), .D[13](w5740), .q[14](w5333), .D[14](w5731), .q[15](w5326), .D[15](w5730), .q[16](w5310), .D[16](w5729), .q[17](w5303), .D[17](w5732), .q[18](w5704), .D[18](w5737), .q[19](w5708), .D[19](w5733), .q[20](w5735), .D[20](w5734), .q[21](w5332), .D[21](w5728), .q[22](w5327), .D[22](w5727), .q[23](w5309), .D[23](w5726), .q[24](w5304), .D[24](w5719), .q[25](w5705), .D[25](w5717), .q[26](w5707), .D[26](w5725), .q[27](w5736), .D[27](w5724), .CLK(w4514), .A[5](w4508), .A[4](w4509), .A[3](w4510), .A[2](w4511), .A[1](w4512), .A[0](w4513), .A(w5739), .B(w5700), .C(w5699), .D(w5698) );
	vdp_linebuf_ram g6312 (.q[0](w5370), .D[0](w5731), .q[1](w5341), .D[1](w5730), .q[2](w5316), .D[2](w5729), .q[3](w5299), .D[3](w5365), .q[4](w5340), .D[4](w5331), .q[5](w5339), .D[5](w5330), .q[6](w5718), .D[6](w5387), .q[7](w5338), .D[7](w5728), .q[8](w5321), .D[8](w5727), .q[9](w5315), .D[9](w5726), .q[10](w5378), .D[10](w5363), .q[11](w5319), .D[11](w5329), .q[12](w5320), .D[12](w5328), .q[13](w5714), .D[13](w5359), .q[14](w5337), .D[14](w5731), .q[15](w5322), .D[15](w5730), .q[16](w5314), .D[16](w5729), .q[17](w5384), .D[17](w5345), .q[18](w5317), .D[18](w5308), .q[19](w5318), .D[19](w5343), .q[20](w5713), .D[20](w5344), .q[21](w5336), .D[21](w5728), .q[22](w5323), .D[22](w5727), .q[23](w5313), .D[23](w5726), .q[24](w5379), .D[24](w6379), .q[25](w5712), .D[25](w5307), .q[26](w5710), .D[26](w5306), .q[27](w5720), .D[27](w5305), .A[0](w4513), .CLK(w4514), .A[5](w4508), .A[3](w4510), .A[4](w4509), .A[2](w4511), .A[1](w4512), .A(w5429), .B(w5413), .C(w5425), .D(w5415) );
	vdp_att_cashe_ram2 g6313 (.q[0](w4715), .D[0](FIFOo[0]), .q[1](w4714), .D[1](FIFOo[1]), .q[2](w4713), .D[2](FIFOo[2]), .q[3](w4712), .D[3](FIFOo[3]), .q[4](w4688), .D[4](FIFOo[4]), .q[5](w4687), .D[5](w172), .q[6](w4682), .D[6](FIFOo[6]), .q[7](w4856), .D[7](w6396), .q[8](w4894), .D[8](w6397), .q[9](w4879), .D[9](w6398), .q[10](w4876), .D[10](w6399), .CLK(HCLK1), .A[6](w6404), .A[5](w6405), .A[1](w6410), .A[0](w6409), .A[4](w6406), .A[3](w6407), .A[2](w6408), .A(w6401), .B(w4701) );
	vdp_att_cashe_ram1 g6314 (.q[0](w4747), .D[0](FIFOo[0]), .q[1](w4750), .D[1](FIFOo[1]), .q[2](w4743), .D[2](FIFOo[2]), .q[3](w4744), .D[3](FIFOo[3]), .q[4](w4726), .D[4](FIFOo[4]), .q[5](w4718), .D[5](w172), .q[6](w4719), .D[6](FIFOo[6]), .q[7](w4717), .D[7](FIFOo[7]), .q[8](w4716), .D[8](w6396), .q[9](w4711), .D[9](w6397), .CLK(HCLK1), .A[0](w6409), .A[1](w6410), .A[2](w6408), .A[3](w6407), .A[4](w6406), .A[5](w6405), .A[6](w6404), .A(w6403), .B(w6402) );
	vdp_att_temp_ram g6315 (.A[4](w4613), .A[0](w4617), .A[1](w4616), .A[2](w4615), .A[3](w4614), .q[0](w6286), .D[0](w6321), .q[1](w6329), .D[1](w6322), .q[2](w6288), .D[2](w6324), .q[3](w6287), .D[3](w6319), .q[4](w6294), .D[4](w6320), .q[5](w6293), .D[5](w6323), .q[6](w6291), .D[6](w6325), .q[7](w6292), .D[7](w6326), .q[8](w6290), .D[8](w6327), .q[9](w6283), .D[9](w6282), .q[10](w6298), .D[10](w6299), .q[11](w6300), .D[11](w6301), .q[12](w6302), .D[12](w6303), .q[13](w6304), .D[13](w6305), .q[14](w6306), .D[14](w6307), .q[15](w6308), .D[15](w6309), .q[16](w6310), .D[16](w6311), .q[17](w6312), .D[17](w6313), .q[18](w6315), .D[18](w6316), .q[19](w6314), .D[19](w6317), .q[20](w6331), .D[20](w6342), .q[21](w6341), .D[21](w6345), .q[22](w6344), .D[22](w6347), .q[23](w6348), .D[23](w6356), .q[24](w6279), .D[24](w6353), .q[25](w6275), .D[25](w6351), .q[26](w6350), .D[26](w6349), .q[26](w6369), .D[26](w6368), .q[27](w6367), .D[27](w6366), .q[28](w6365), .D[28](w6364), .q[29](w6363), .D[29](w6362), .q[30](w6361), .D[30](w6360), .q[31](w6375), .D[31](w6359), .q[32](w6358), .D[32](w6357), .CLK(HCLK1), .A(w4580), .B(w4581), .C(w4585) );
	vdp_vsram g6316 (.CLK(HCLK1), .D[10](w4001), .q[10](w3959), .D[9](w4005), .q[9](w3952), .D[8](w4003), .q[8](w3978), .D[7](w4002), .q[7](w3944), .D[6](w3990), .q[6](w3940), .D[5](w3988), .q[5](w3932), .D[4](w3995), .q[4](w3928), .D[3](w3997), .q[3](w3925), .D[2](w4000), .q[2](w3983), .D[1](w3958), .q[1](w3920), .D[0](w3976), .q[0](w3915), .A[1](w3732), .A[2](w3704), .A[3](w3703), .A[4](w3702), .A[5](w3701), .A[0](w3733), .A(w3700), .B(w3699) );
	vdp_not g6317 (.nZ(w1820), .A(w6707) );
	vdp_not g6318 (.nZ(PAL), .A(w6708) );
	vdp_H_PLA g6319 (.HPLA[0](w1939), .HPLA[1](w1920), .HPLA[2](w1912), .HPLA[3](w1749), .HPLA[4](w1910), .HPLA[5](w1913), .HPLA[7](w1750), .HPLA[8](w1751), .HPLA[9](w1870), .HPLA[6](w1752), .HPLA[10](w1873), .HPLA[11](w1916), .HPLA[16](w1874), .HPLA[15](w1918), .HPLA[14](w1917), .HPLA[13](w1921), .HPLA[12](w1922), .i0(w59), .HPLA[17](w1772), .HPLA[18](w1771), .HPLA[19](w1872), .HPLA[20](w1871), .HPLA[21](w1914), .HPLA[22](w1909), .Hcnt[0](w1940), .Hcnt[1](w1686), .Hcnt[2](w1691), .Hcnt[3](w1690), .Hcnt[4](w1735), .Hcnt[5](w1769), .Hcnt[6](w1915), .Hcnt[7](w1746), .Hcnt[8](w1774), .H40(H40), .M5(M5), .B(w1773), .C(w1670), .A(w1740), .HPLA[23](w1689), .HPLA[24](w1687), .HPLA[25](w1688), .HPLA[26](w1685), .HPLA[27](w1875), .HPLA[28](w1868), .HPLA[29](w1671), .HPLA[30](w1724), .HPLA[31](w1672), .HPLA[32](w1911), .HPLA[33](w1766), .3(w1919), .HPLA[35](w1802), .HPLA[36](w1764), .HPLA[34](w1941) );
	vdp_slatch g5073 (.D(S[4]), .nC(w5029), .C(w5030), .Q(w5225) );
endmodule // VDP

// Module Definitions [It is possible to wrap here on your primitives]

module vdp_slatch (  nQ, D, C, nC);

	output wire nQ;
	input wire D;
	input wire C;
	input wire nC;

endmodule // vdp_slatch

module vdp_sr_bit (  D, C2, C1, Q, nC2, nC1);

	input wire D;
	input wire C2;
	input wire C1;
	output wire Q;
	input wire nC2;
	input wire nC1;

endmodule // vdp_sr_bit

module vdp_notif0 (  A, nZ, nE);

	input wire A;
	output wire nZ;
	input wire nE;

endmodule // vdp_notif0

module vdp_aon22 (  Z, A1, A2, B1, B2);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire B1;
	input wire B2;

endmodule // vdp_aon22

module vdp_not (  A, nZ);

	input wire A;
	output wire nZ;

endmodule // vdp_not

module vdp_comp_str (  A, Z, nZ);

	input wire A;
	output wire Z;
	output wire nZ;

endmodule // vdp_comp_str

module vdp_comp_we (  A, Z, nZ);

	input wire A;
	output wire Z;
	output wire nZ;

endmodule // vdp_comp_we

module vdp_and (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_and

module vdp_nand (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_nand

module vdp_and3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_and3

module vdp_fa (  SUM, A, B, CO, CI);

	output wire SUM;
	input wire A;
	input wire B;
	output wire CO;
	input wire CI;

endmodule // vdp_fa

module vdp_comp_dff (  D, C2, C1, Q, nC2, nC1);

	input wire D;
	input wire C2;
	input wire C1;
	output wire Q;
	input wire nC2;
	input wire nC1;

endmodule // vdp_comp_dff

module vdp_or (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_or

module vdp_xor (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_xor

module vdp_aoi21 (  Z, B, A1, A2);

	output wire Z;
	input wire B;
	input wire A1;
	input wire A2;

endmodule // vdp_aoi21

module vdp_nor (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // vdp_nor

module vdp_and5 (  Z, A, B, C, D, E);

	output wire Z;
	input wire A;
	input wire B;
	input wire C;
	input wire D;
	input wire E;

endmodule // vdp_and5

module vdp_aon2222 (  C2, B2, A2, C1, B1, A1, Z, D2, D1);

	input wire C2;
	input wire B2;
	input wire A2;
	input wire C1;
	input wire B1;
	input wire A1;
	output wire Z;
	input wire D2;
	input wire D1;

endmodule // vdp_aon2222

module vdp_cnt_bit (  R, Q, C1, C2, nC1, nC2, CI);

	input wire R;
	output wire Q;
	input wire C1;
	input wire C2;
	input wire nC1;
	input wire nC2;
	input wire CI;

endmodule // vdp_cnt_bit

module vdp_oai21 (  A1, Z, A2, B);

	input wire A1;
	output wire Z;
	input wire A2;
	input wire B;

endmodule // vdp_oai21

module vdp_comb1 (  Z, A1, B, A2, C);

	output wire Z;
	input wire A1;
	input wire B;
	input wire A2;
	input wire C;

endmodule // vdp_comb1

module vdp_rs_ff (  Q, R, S);

	output wire Q;
	input wire R;
	input wire S;

endmodule // vdp_rs_ff

module vdp_and4 (  A, Z, B, C, D);

	input wire A;
	output wire Z;
	input wire B;
	input wire C;
	input wire D;

endmodule // vdp_and4

module vdp_or3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_or3

module vdp_bufif0 (  A, Z, nE);

	input wire A;
	output wire Z;
	input wire nE;

endmodule // vdp_bufif0

module vdp_aoi221 (  Z, A2, B1, B2, A1, C);

	output wire Z;
	input wire A2;
	input wire B1;
	input wire B2;
	input wire A1;
	input wire C;

endmodule // vdp_aoi221

module vdp_aon33 (  Z, A2, B1, B2, A1, A3, B3);

	output wire Z;
	input wire A2;
	input wire B1;
	input wire B2;
	input wire A1;
	input wire A3;
	input wire B3;

endmodule // vdp_aon33

module vdp_dlatch_inv (  D, C, Q, nC);

	input wire D;
	input wire C;
	output wire Q;
	input wire nC;

endmodule // vdp_dlatch_inv

module vdp_cnt_bit_load (  D, nL, L, R, Q, C1, C2, nC1, nC2, CI, CO);

	input wire D;
	input wire nL;
	input wire L;
	input wire R;
	output wire Q;
	input wire C1;
	input wire C2;
	input wire nC1;
	input wire nC2;
	input wire CI;
	output wire CO;

endmodule // vdp_cnt_bit_load

module vdp_nand3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_nand3

module vdp_nor3 (  Z, B, A, C);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;

endmodule // vdp_nor3

module vdp_dff (  Q, R, C, D);

	output wire Q;
	input wire R;
	input wire C;
	input wire D;

endmodule // vdp_dff

module vdp_ha (  SUM, A, B, CO);

	output wire SUM;
	input wire A;
	input wire B;
	output wire CO;

endmodule // vdp_ha

module vdp_slatch_r (  Q, D, R, C, nC);

	output wire Q;
	input wire D;
	input wire R;
	input wire C;
	input wire nC;

endmodule // vdp_slatch_r

module vdp_rs_FF (  nQ, R, S, Q);

	output wire nQ;
	input wire R;
	input wire S;
	output wire Q;

endmodule // vdp_rs_FF

module vdp_or5 (  C, A, B, Z, D, E);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;
	input wire E;

endmodule // vdp_or5

module vdp_2a3oi (  A1, B, Z, A2, C);

	input wire A1;
	input wire B;
	output wire Z;
	input wire A2;
	input wire C;

endmodule // vdp_2a3oi

module vdp_nor5 (  C, A, B, Z, D, E);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;
	input wire E;

endmodule // vdp_nor5

module vdp_or4 (  C, A, B, Z, D);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;

endmodule // vdp_or4

module vdp_aoi22 (  Z, A1, A2, B1, B2);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire B1;
	input wire B2;

endmodule // vdp_aoi22

module vdp_aon222 (  C2, B2, A2, C1, B1, A1, Z);

	input wire C2;
	input wire B2;
	input wire A2;
	input wire C1;
	input wire B1;
	input wire A1;
	output wire Z;

endmodule // vdp_aon222

module vdp_dslatch (  D, C, Q, nC);

	input wire D;
	input wire C;
	output wire Q;
	input wire nC;

endmodule // vdp_dslatch

module vdp_comp_DFF (  D, C2, C1, Q, nC2, nC1);

	input wire D;
	input wire C2;
	input wire C1;
	output wire Q;
	input wire nC2;
	input wire nC1;

endmodule // vdp_comp_DFF

module vdp_nor4 (  C, A, B, Z, D);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;

endmodule // vdp_nor4

module vdp_and6 (  C, A, B, Z, D, E, F);

	input wire C;
	input wire A;
	input wire B;
	output wire Z;
	input wire D;
	input wire E;
	input wire F;

endmodule // vdp_and6

module vdp_g1622 (  Z, A);

	output wire Z;
	input wire A;

endmodule // vdp_g1622

module vdp_g1623 (  Z, A);

	output wire Z;
	input wire A;

endmodule // vdp_g1623

module vdp_g1624 (  A, Z);

	input wire A;
	output wire Z;

endmodule // vdp_g1624

module vdp_g1625 (  A, Z);

	input wire A;
	output wire Z;

endmodule // vdp_g1625

module vdp_g1626 (  Z, A);

	output wire Z;
	input wire A;

endmodule // vdp_g1626

module vdp_g1627 (  Z, A);

	output wire Z;
	input wire A;

endmodule // vdp_g1627

module vdp_g1628 (  Z, A);

	output wire Z;
	input wire A;

endmodule // vdp_g1628

module vdp_g1629 (  Z, A);

	output wire Z;
	input wire A;

endmodule // vdp_g1629

module vdp_2?3?I (  Z, A1, A2, C, B);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire C;
	input wire B;

endmodule // vdp_2?3?I

module vdp_RS (  Q, S, R);

	output wire Q;
	input wire S;
	input wire R;

endmodule // vdp_RS

module vdp_TFF (  C2, C1, nC2, nC1, CI, R, A, Q);

	input wire C2;
	input wire C1;
	input wire nC2;
	input wire nC1;
	input wire CI;
	input wire R;
	input wire A;
	output wire Q;

endmodule // vdp_TFF

module vdp_comp_ (  Q, D, nC1, C1, nC2, C2);

	output wire Q;
	input wire D;
	input wire nC1;
	input wire C1;
	input wire nC2;
	input wire C2;

endmodule // vdp_comp_

module vdp_SDELAY8 (  Q, D, nC1, C1, nC2, C2, nC3, C3, nC4, C4, nC5, C5, nC6, C6, nC7, C7, nC8, C8, nC9, C9, nC10, C10, nC11, C11, nC12, C12, nC13, C13, nC14, C14, nC15, C15, nC16, C16);

	output wire Q;
	input wire D;
	input wire nC1;
	input wire C1;
	input wire nC2;
	input wire C2;
	input wire nC3;
	input wire C3;
	input wire nC4;
	input wire C4;
	input wire nC5;
	input wire C5;
	input wire nC6;
	input wire C6;
	input wire nC7;
	input wire C7;
	input wire nC8;
	input wire C8;
	input wire nC9;
	input wire C9;
	input wire nC10;
	input wire C10;
	input wire nC11;
	input wire C11;
	input wire nC12;
	input wire C12;
	input wire nC13;
	input wire C13;
	input wire nC14;
	input wire C14;
	input wire nC15;
	input wire C15;
	input wire nC16;
	input wire C16;

endmodule // vdp_SDELAY8

module vdp_SDELAY7 (  Q, D, C1, nC1, C2, nC2, nC3, C4, nC4, C5, nC5, C6, nC6, C7, nC7, C8, nC8, C9, nC9, C10, nC10, C11, nC11, C12, nC12, C13, nC13, C14, nC14, C3);

	output wire Q;
	input wire D;
	input wire C1;
	input wire nC1;
	input wire C2;
	input wire nC2;
	input wire nC3;
	input wire C4;
	input wire nC4;
	input wire C5;
	input wire nC5;
	input wire C6;
	input wire nC6;
	input wire C7;
	input wire nC7;
	input wire C8;
	input wire nC8;
	input wire C9;
	input wire nC9;
	input wire C10;
	input wire nC10;
	input wire C11;
	input wire nC11;
	input wire C12;
	input wire nC12;
	input wire C13;
	input wire nC13;
	input wire C14;
	input wire nC14;
	input wire C3;

endmodule // vdp_SDELAY7

module vdp_or8 (  Z, A, B, C, D, E, F, G, H);

	output wire Z;
	input wire A;
	input wire B;
	input wire C;
	input wire D;
	input wire E;
	input wire F;
	input wire G;
	input wire H;

endmodule // vdp_or8

module vdp_or7 (  Z, A, B, C, D, E, F, G);

	output wire Z;
	input wire A;
	input wire B;
	input wire C;
	input wire D;
	input wire E;
	input wire F;
	input wire G;

endmodule // vdp_or7

module vdp_dlatch (  Q, C, D, nC);

	output wire Q;
	input wire C;
	input wire D;
	input wire nC;

endmodule // vdp_dlatch

module vdp_clkgen (  PH, CLK1, nCLK1, CLK2, nCLK2);

	input wire PH;
	output wire CLK1;
	output wire nCLK1;
	output wire CLK2;
	output wire nCLK2;

endmodule // vdp_clkgen

module vdp_cgi2a (  Z, A, C, B);

	output wire Z;
	input wire A;
	input wire C;
	input wire B;

endmodule // vdp_cgi2a

module vdp_nand4 (  Z, A, B, D, C);

	output wire Z;
	input wire A;
	input wire B;
	input wire D;
	input wire C;

endmodule // vdp_nand4

module vdp_lfsr_bit (  Q, A, C2, C1, nC2, nC1, C, B);

	output wire Q;
	input wire A;
	input wire C2;
	input wire C1;
	input wire nC2;
	input wire nC1;
	input wire C;
	input wire B;

endmodule // vdp_lfsr_bit

module vdp_aoi222 (  Z, A1, B1, B2, A2, C1, C2);

	output wire Z;
	input wire A1;
	input wire B1;
	input wire B2;
	input wire A2;
	input wire C1;
	input wire C2;

endmodule // vdp_aoi222

module vdp_aon333 (  Z, A1, A2, A3, B1, B2, B3, C1, C2, C3);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire A3;
	input wire B1;
	input wire B2;
	input wire B3;
	input wire C1;
	input wire C2;
	input wire C3;

endmodule // vdp_aon333

module vdp_aoi33 (  Z, A1, A2, A3, B1, B2, B3);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire A3;
	input wire B1;
	input wire B2;
	input wire B3;

endmodule // vdp_aoi33

module vdp_comp_strong (  nZ, Z, A);

	output wire nZ;
	output wire Z;
	input wire A;

endmodule // vdp_comp_strong

module vdp_neg_dff (  Q, C, D, R);

	output wire Q;
	input wire C;
	input wire D;
	input wire R;

endmodule // vdp_neg_dff

module vdp_buf (  Z, A);

	output wire Z;
	input wire A;

endmodule // vdp_buf

module vdp_g2925 (  Z, A, B, C, D);

	output wire Z;
	input wire A;
	input wire B;
	input wire C;
	input wire D;

endmodule // vdp_g2925

module vdp_g2938 (  A, Z);

	input wire A;
	output wire Z;

endmodule // vdp_g2938

module vdp_aon2*8 (  Z, A1, B1, C1, D2, A2, B2, C2, D1, E2, F1, E1, F2, G1, H2, G2, H1);

	output wire Z;
	input wire A1;
	input wire B1;
	input wire C1;
	input wire D2;
	input wire A2;
	input wire B2;
	input wire C2;
	input wire D1;
	input wire E2;
	input wire F1;
	input wire E1;
	input wire F2;
	input wire G1;
	input wire H2;
	input wire G2;
	input wire H1;

endmodule // vdp_aon2*8

module vdp_xnor (  Z, A, B);

	output wire Z;
	input wire A;
	input wire B;

endmodule // vdp_xnor

module vdp_oai211 (  Z, A1, A2, B, C);

	output wire Z;
	input wire A1;
	input wire A2;
	input wire B;
	input wire C;

endmodule // vdp_oai211

module vdp_aoi31 (  Z, B3, B2, B1, A);

	output wire Z;
	input wire B3;
	input wire B2;
	input wire B1;
	input wire A;

endmodule // vdp_aoi31

module vdp_AOI222 (  Z, B1, A1, B2, A2, C1, C2);

	output wire Z;
	input wire B1;
	input wire A1;
	input wire B2;
	input wire A2;
	input wire C1;
	input wire C2;

endmodule // vdp_AOI222

module vdp_SR_bit (  Q, D, C1, C2, nC1, nC2);

	output wire Q;
	input wire D;
	input wire C1;
	input wire C2;
	input wire nC1;
	input wire nC2;

endmodule // vdp_SR_bit

module vdp_cnt_bit_rev (  nC2, nC1, C2, C1, Q, CI, B, A);

	input wire nC2;
	input wire nC1;
	input wire C2;
	input wire C1;
	output wire Q;
	input wire CI;
	input wire B;
	input wire A;

endmodule // vdp_cnt_bit_rev

module vdp_2x_sr_bit (  Q, D, nC2, nC1, C2, C1, nC4, nC3, C4, C3);

	output wire Q;
	input wire D;
	input wire nC2;
	input wire nC1;
	input wire C2;
	input wire C1;
	input wire nC4;
	input wire nC3;
	input wire C4;
	input wire C3;

endmodule // vdp_2x_sr_bit

module vdp_and9 (  Z, B, A, C, D, F, E, G, H, I);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;
	input wire I;

endmodule // vdp_and9

module vdp_nor12 (  Z, B, A, C, D, F, E, G, H, J, I, K, L);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;
	input wire J;
	input wire I;
	input wire K;
	input wire L;

endmodule // vdp_nor12

module vdp_noif0 (  A, nZ, nE);

	input wire A;
	output wire nZ;
	input wire nE;

endmodule // vdp_noif0

module vdp_nor8 (  Z, B, A, C, D, F, E, G, H);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;

endmodule // vdp_nor8

module vdp_aon21_sr (  Q, A1, A2, B, nC2, nC1, C2, C1);

	output wire Q;
	input wire A1;
	input wire A2;
	input wire B;
	input wire nC2;
	input wire nC1;
	input wire C2;
	input wire C1;

endmodule // vdp_aon21_sr

module vdp_or9 (  Z, B, A, C, D, F, E, G, H, I);

	output wire Z;
	input wire B;
	input wire A;
	input wire C;
	input wire D;
	input wire F;
	input wire E;
	input wire G;
	input wire H;
	input wire I;

endmodule // vdp_or9

module vdp_V_PLA (  o[0], o[1], o[2], o[3], o[4], o[5], o[6], o[7], o[8], o[9], o[10], o[11], o[12], o[13], o[14], o[15], o[16], o[17], o[18], o[19], o[20], o[21], o[22], o[23], o[24], o[25], o[26], o[27], o[28], o[29], o[30], o[31], o[32], o[33], o[34], o[35], o[36], o[37], o[38], o[39], o[40], o[41], o[42], o[43], o[44], o[45], o[46], o[47], Vcnt[0], Vcnt[1], Vcnt[2], Vcnt[3], Vcnt[4], Vcnt[5], Vcnt[6], Vcnt[7], Vcnt[8], ODD_EVEN, LS0, PAL, nPAL, 2, 3, M5);

	output wire o[0];
	output wire o[1];
	output wire o[2];
	output wire o[3];
	output wire o[4];
	output wire o[5];
	output wire o[6];
	output wire o[7];
	output wire o[8];
	output wire o[9];
	output wire o[10];
	output wire o[11];
	output wire o[12];
	output wire o[13];
	output wire o[14];
	output wire o[15];
	output wire o[16];
	output wire o[17];
	output wire o[18];
	output wire o[19];
	output wire o[20];
	output wire o[21];
	output wire o[22];
	output wire o[23];
	output wire o[24];
	output wire o[25];
	output wire o[26];
	output wire o[27];
	output wire o[28];
	output wire o[29];
	output wire o[30];
	output wire o[31];
	output wire o[32];
	output wire o[33];
	output wire o[34];
	output wire o[35];
	output wire o[36];
	output wire o[37];
	output wire o[38];
	output wire o[39];
	output wire o[40];
	output wire o[41];
	output wire o[42];
	output wire o[43];
	output wire o[44];
	output wire o[45];
	output wire o[46];
	output wire o[47];
	input wire Vcnt[0];
	input wire Vcnt[1];
	input wire Vcnt[2];
	input wire Vcnt[3];
	input wire Vcnt[4];
	input wire Vcnt[5];
	input wire Vcnt[6];
	input wire Vcnt[7];
	input wire Vcnt[8];
	input wire ODD_EVEN;
	input wire LS0;
	input wire PAL;
	input wire nPAL;
	input wire 2;
	input wire 3;
	input wire M5;

endmodule // vdp_V_PLA

module vdp_cram (  q[8], D[8], q[7], D[7], q[6], D[6], q[5], D[5], q[4], D[4], q[3], D[3], q[2], D[2], q[1], D[1], q[0], D[0], A[0], A[1], CLK, A[2], A[3], A[4], A[5], B, A);

	output wire q[8];
	input wire D[8];
	output wire q[7];
	input wire D[7];
	output wire q[6];
	input wire D[6];
	output wire q[5];
	input wire D[5];
	output wire q[4];
	input wire D[4];
	output wire q[3];
	input wire D[3];
	output wire q[2];
	input wire D[2];
	output wire q[1];
	input wire D[1];
	output wire q[0];
	input wire D[0];
	input wire A[0];
	input wire A[1];
	input wire CLK;
	input wire A[2];
	input wire A[3];
	input wire A[4];
	input wire A[5];
	input wire B;
	input wire A;

endmodule // vdp_cram

module vdp_linebuf_ram (  q[0], D[0], q[1], D[1], q[2], D[2], q[3], D[3], q[4], D[4], q[5], D[5], q[6], D[6], q[7], D[7], q[8], D[8], q[9], D[9], q[10], D[10], q[11], D[11], q[12], D[12], q[13], D[13], q[14], D[14], q[15], D[15], q[16], D[16], q[17], D[17], q[18], D[18], q[19], D[19], q[20], D[20], q[21], D[21], q[22], D[22], q[23], D[23], q[24], D[24], q[25], D[25], q[26], D[26], q[27], D[27], CLK, A[5], A[4], A[3], A[2], A[1], A[0], A, B, C, D);

	output wire q[0];
	input wire D[0];
	output wire q[1];
	input wire D[1];
	output wire q[2];
	input wire D[2];
	output wire q[3];
	input wire D[3];
	output wire q[4];
	input wire D[4];
	output wire q[5];
	input wire D[5];
	output wire q[6];
	input wire D[6];
	output wire q[7];
	input wire D[7];
	output wire q[8];
	input wire D[8];
	output wire q[9];
	input wire D[9];
	output wire q[10];
	input wire D[10];
	output wire q[11];
	input wire D[11];
	output wire q[12];
	input wire D[12];
	output wire q[13];
	input wire D[13];
	output wire q[14];
	input wire D[14];
	output wire q[15];
	input wire D[15];
	output wire q[16];
	input wire D[16];
	output wire q[17];
	input wire D[17];
	output wire q[18];
	input wire D[18];
	output wire q[19];
	input wire D[19];
	output wire q[20];
	input wire D[20];
	output wire q[21];
	input wire D[21];
	output wire q[22];
	input wire D[22];
	output wire q[23];
	input wire D[23];
	output wire q[24];
	input wire D[24];
	output wire q[25];
	input wire D[25];
	output wire q[26];
	input wire D[26];
	output wire q[27];
	input wire D[27];
	input wire CLK;
	input wire A[5];
	input wire A[4];
	input wire A[3];
	input wire A[2];
	input wire A[1];
	input wire A[0];
	input wire A;
	input wire B;
	input wire C;
	input wire D;

endmodule // vdp_linebuf_ram

module vdp_att_cashe_ram2 (  q[0], D[0], q[1], D[1], q[2], D[2], q[3], D[3], q[4], D[4], q[5], D[5], q[6], D[6], q[7], D[7], q[8], D[8], q[9], D[9], q[10], D[10], CLK, A[6], A[5], A[1], A[0], A[4], A[3], A[2], A, B);

	output wire q[0];
	input wire D[0];
	output wire q[1];
	input wire D[1];
	output wire q[2];
	input wire D[2];
	output wire q[3];
	input wire D[3];
	output wire q[4];
	input wire D[4];
	output wire q[5];
	input wire D[5];
	output wire q[6];
	input wire D[6];
	output wire q[7];
	input wire D[7];
	output wire q[8];
	input wire D[8];
	output wire q[9];
	input wire D[9];
	output wire q[10];
	input wire D[10];
	input wire CLK;
	input wire A[6];
	input wire A[5];
	input wire A[1];
	input wire A[0];
	input wire A[4];
	input wire A[3];
	input wire A[2];
	input wire A;
	input wire B;

endmodule // vdp_att_cashe_ram2

module vdp_att_cashe_ram1 (  q[0], D[0], q[1], D[1], q[2], D[2], q[3], D[3], q[4], D[4], q[5], D[5], q[6], D[6], q[7], D[7], q[8], D[8], q[9], D[9], CLK, A[0], A[1], A[2], A[3], A[4], A[5], A[6], A, B);

	output wire q[0];
	input wire D[0];
	output wire q[1];
	input wire D[1];
	output wire q[2];
	input wire D[2];
	output wire q[3];
	input wire D[3];
	output wire q[4];
	input wire D[4];
	output wire q[5];
	input wire D[5];
	output wire q[6];
	input wire D[6];
	output wire q[7];
	input wire D[7];
	output wire q[8];
	input wire D[8];
	output wire q[9];
	input wire D[9];
	input wire CLK;
	input wire A[0];
	input wire A[1];
	input wire A[2];
	input wire A[3];
	input wire A[4];
	input wire A[5];
	input wire A[6];
	input wire A;
	input wire B;

endmodule // vdp_att_cashe_ram1

module vdp_att_temp_ram (  A[4], A[0], A[1], A[2], A[3], q[0], D[0], q[1], D[1], q[2], D[2], q[3], D[3], q[4], D[4], q[5], D[5], q[6], D[6], q[7], D[7], q[8], D[8], q[9], D[9], q[10], D[10], q[11], D[11], q[12], D[12], q[13], D[13], q[14], D[14], q[15], D[15], q[16], D[16], q[17], D[17], q[18], D[18], q[19], D[19], q[20], D[20], q[21], D[21], q[22], D[22], q[23], D[23], q[24], D[24], q[25], D[25], q[26], D[26], q[26], D[26], q[27], D[27], q[28], D[28], q[29], D[29], q[30], D[30], q[31], D[31], q[32], D[32], CLK, A, B, C);

	input wire A[4];
	input wire A[0];
	input wire A[1];
	input wire A[2];
	input wire A[3];
	output wire q[0];
	input wire D[0];
	output wire q[1];
	input wire D[1];
	output wire q[2];
	input wire D[2];
	output wire q[3];
	input wire D[3];
	output wire q[4];
	input wire D[4];
	output wire q[5];
	input wire D[5];
	output wire q[6];
	input wire D[6];
	output wire q[7];
	input wire D[7];
	output wire q[8];
	input wire D[8];
	output wire q[9];
	input wire D[9];
	output wire q[10];
	input wire D[10];
	output wire q[11];
	input wire D[11];
	output wire q[12];
	input wire D[12];
	output wire q[13];
	input wire D[13];
	output wire q[14];
	input wire D[14];
	output wire q[15];
	input wire D[15];
	output wire q[16];
	input wire D[16];
	output wire q[17];
	input wire D[17];
	output wire q[18];
	input wire D[18];
	output wire q[19];
	input wire D[19];
	output wire q[20];
	input wire D[20];
	output wire q[21];
	input wire D[21];
	output wire q[22];
	input wire D[22];
	output wire q[23];
	input wire D[23];
	output wire q[24];
	input wire D[24];
	output wire q[25];
	input wire D[25];
	output wire q[26];
	input wire D[26];
	output wire q[26];
	input wire D[26];
	output wire q[27];
	input wire D[27];
	output wire q[28];
	input wire D[28];
	output wire q[29];
	input wire D[29];
	output wire q[30];
	input wire D[30];
	output wire q[31];
	input wire D[31];
	output wire q[32];
	input wire D[32];
	input wire CLK;
	input wire A;
	input wire B;
	input wire C;

endmodule // vdp_att_temp_ram

module vdp_vsram (  CLK, D[10], q[10], D[9], q[9], D[8], q[8], D[7], q[7], D[6], q[6], D[5], q[5], D[4], q[4], D[3], q[3], D[2], q[2], D[1], q[1], D[0], q[0], A[1], A[2], A[3], A[4], A[5], A[0], A, B);

	input wire CLK;
	input wire D[10];
	output wire q[10];
	input wire D[9];
	output wire q[9];
	input wire D[8];
	output wire q[8];
	input wire D[7];
	output wire q[7];
	input wire D[6];
	output wire q[6];
	input wire D[5];
	output wire q[5];
	input wire D[4];
	output wire q[4];
	input wire D[3];
	output wire q[3];
	input wire D[2];
	output wire q[2];
	input wire D[1];
	output wire q[1];
	input wire D[0];
	output wire q[0];
	input wire A[1];
	input wire A[2];
	input wire A[3];
	input wire A[4];
	input wire A[5];
	input wire A[0];
	input wire A;
	input wire B;

endmodule // vdp_vsram

module vdp_H_PLA (  HPLA[0], HPLA[1], HPLA[2], HPLA[3], HPLA[4], HPLA[5], HPLA[7], HPLA[8], HPLA[9], HPLA[6], HPLA[10], HPLA[11], HPLA[16], HPLA[15], HPLA[14], HPLA[13], HPLA[12], i0, HPLA[17], HPLA[18], HPLA[19], HPLA[20], HPLA[21], HPLA[22], Hcnt[0], Hcnt[1], Hcnt[2], Hcnt[3], Hcnt[4], Hcnt[5], Hcnt[6], Hcnt[7], Hcnt[8], H40, M5, B, C, A, HPLA[23], HPLA[24], HPLA[25], HPLA[26], HPLA[27], HPLA[28], HPLA[29], HPLA[30], HPLA[31], HPLA[32], HPLA[33], 3, HPLA[35], HPLA[36], HPLA[34]);

	output wire HPLA[0];
	output wire HPLA[1];
	output wire HPLA[2];
	output wire HPLA[3];
	output wire HPLA[4];
	output wire HPLA[5];
	output wire HPLA[7];
	output wire HPLA[8];
	output wire HPLA[9];
	output wire HPLA[6];
	output wire HPLA[10];
	output wire HPLA[11];
	output wire HPLA[16];
	output wire HPLA[15];
	output wire HPLA[14];
	output wire HPLA[13];
	output wire HPLA[12];
	input wire i0;
	output wire HPLA[17];
	output wire HPLA[18];
	output wire HPLA[19];
	output wire HPLA[20];
	output wire HPLA[21];
	output wire HPLA[22];
	input wire Hcnt[0];
	input wire Hcnt[1];
	input wire Hcnt[2];
	input wire Hcnt[3];
	input wire Hcnt[4];
	input wire Hcnt[5];
	input wire Hcnt[6];
	input wire Hcnt[7];
	input wire Hcnt[8];
	input wire H40;
	input wire M5;
	input wire B;
	input wire C;
	input wire A;
	output wire HPLA[23];
	output wire HPLA[24];
	output wire HPLA[25];
	output wire HPLA[26];
	output wire HPLA[27];
	output wire HPLA[28];
	output wire HPLA[29];
	output wire HPLA[30];
	output wire HPLA[31];
	output wire HPLA[32];
	output wire HPLA[33];
	input wire 3;
	output wire HPLA[35];
	output wire HPLA[36];
	output wire HPLA[34];

endmodule // vdp_H_PLA



// ERROR: conflicting wire VRAMA[8]
// WARNING: wire not driving anything w128
// ERROR: conflicting wire AD_DATA[7]
// ERROR: conflicting wire AD_DATA[6]
// ERROR: conflicting wire AD_DATA[4]
// ERROR: conflicting wire RD_DATA[2]
// ERROR: conflicting wire RD_DATA[1]
// ERROR: conflicting wire RD_DATA[0]
// ERROR: conflicting wire AD_DATA[5]
// ERROR: conflicting wire nDCLK2
// ERROR: conflicting wire DB[0]
// ERROR: conflicting wire DB[1]
// ERROR: conflicting wire DB[2]
// ERROR: conflicting wire DB[3]
// ERROR: conflicting wire DB[4]
// ERROR: conflicting wire DB[5]
// ERROR: conflicting wire DB[6]
// ERROR: conflicting wire DB[7]
// ERROR: conflicting wire DB[8]
// ERROR: conflicting wire DB[9]
// ERROR: conflicting wire AD_DATA[3]
// ERROR: conflicting wire AD_DATA[2]
// ERROR: conflicting wire AD_DATA[1]
// ERROR: conflicting wire AD_DATA[0]
// ERROR: conflicting wire DB[14]
// ERROR: conflicting wire DB[13]
// ERROR: conflicting wire DB[12]
// ERROR: conflicting wire DB[11]
// ERROR: conflicting wire DB[10]
// ERROR: floating wire w172
// ERROR: floating wire w190
// ERROR: conflicting wire RD_DATA[4]
// ERROR: floating wire w221
// ERROR: conflicting wire RD_DATA[6]
// ERROR: floating wire w237
// ERROR: conflicting wire w239
// ERROR: conflicting wire w247
// ERROR: conflicting wire w256
// ERROR: conflicting wire w264
// ERROR: conflicting wire w281
// ERROR: conflicting wire w290
// ERROR: conflicting wire w291
// ERROR: conflicting wire w300
// ERROR: conflicting wire w308
// ERROR: conflicting wire w324
// ERROR: floating wire w337
// ERROR: conflicting wire RD_DATA[5]
// ERROR: floating wire w353
// ERROR: conflicting wire DB[15]
// ERROR: conflicting wire w358
// ERROR: floating wire w461
// ERROR: conflicting wire VRAMA[0]
// ERROR: floating wire w576
// ERROR: conflicting wire VRAMA[7]
// ERROR: conflicting wire VRAMA[9]
// ERROR: conflicting wire VRAMA[10]
// ERROR: conflicting wire VRAMA[6]
// ERROR: conflicting wire VRAMA[5]
// ERROR: conflicting wire VRAMA[11]
// ERROR: conflicting wire VRAMA[12]
// ERROR: conflicting wire VRAMA[4]
// ERROR: conflicting wire VRAMA[13]
// ERROR: conflicting wire VRAMA[3]
// ERROR: conflicting wire VRAMA[14]
// ERROR: conflicting wire VRAMA[2]
// ERROR: conflicting wire CA[14]
// ERROR: conflicting wire VRAMA[15]
// ERROR: conflicting wire VRAMA[1]
// ERROR: conflicting wire VRAMA[16]
// ERROR: floating wire w798
// ERROR: floating wire w800
// ERROR: floating wire w813
// ERROR: floating wire w814
// ERROR: floating wire w831
// ERROR: floating wire w927
// ERROR: floating wire w929
// ERROR: floating wire w1075
// ERROR: floating wire w1081
// ERROR: conflicting wire COL[0]
// ERROR: conflicting wire COL[1]
// ERROR: conflicting wire COL[2]
// ERROR: conflicting wire COL[3]
// ERROR: conflicting wire COL[4]
// ERROR: conflicting wire COL[5]
// ERROR: conflicting wire COL[6]
// ERROR: floating wire w1098
// ERROR: floating wire w1099
// ERROR: floating wire w1187
// ERROR: floating wire w1208
// ERROR: floating wire w1226
// ERROR: floating wire w1300
// ERROR: floating wire w1307
// ERROR: floating wire w1315
// ERROR: floating wire w1332
// ERROR: floating wire w1363
// ERROR: floating wire w1387
// ERROR: floating wire w1607
// ERROR: floating wire w1684
// ERROR: floating wire w1742
// ERROR: floating wire w1743
// ERROR: floating wire w1787
// ERROR: floating wire w1829
// ERROR: floating wire w1839
// ERROR: floating wire w1984
// ERROR: floating wire w2074
// ERROR: floating wire w2260
// ERROR: floating wire w2295
// ERROR: floating wire w2483
// ERROR: floating wire w2629
// ERROR: floating wire w2635
// ERROR: floating wire w2796
// ERROR: floating wire w3115
// ERROR: floating wire w3121
// ERROR: floating wire w3456
// ERROR: floating wire w3526
// ERROR: floating wire w3606
// ERROR: floating wire w3663
// ERROR: floating wire w3673
// ERROR: floating wire w3674
// ERROR: floating wire w3706
// ERROR: floating wire w3749
// ERROR: floating wire w3754
// ERROR: floating wire w3809
// ERROR: floating wire w3811
// ERROR: floating wire w3887
// ERROR: floating wire w3913
// ERROR: floating wire w3968
// ERROR: floating wire w4087
// ERROR: floating wire w4420
// ERROR: floating wire w4432
// ERROR: floating wire w4505
// ERROR: floating wire w4590
// ERROR: floating wire w4659
// ERROR: floating wire w4664
// ERROR: floating wire w4702
// ERROR: floating wire w4705
// ERROR: floating wire w4760
// ERROR: floating wire w4765
// ERROR: floating wire w4794
// ERROR: floating wire w4838
// ERROR: floating wire w4896
// ERROR: floating wire w4911
// ERROR: floating wire w4918
// ERROR: floating wire w4957
// ERROR: floating wire w5150
// ERROR: floating wire w5207
// ERROR: floating wire w5347
// ERROR: floating wire w5362
// ERROR: floating wire w5366
// ERROR: floating wire w5374
// ERROR: floating wire w5404
// ERROR: floating wire w5468
// ERROR: floating wire w5494
// ERROR: floating wire w5524
// ERROR: floating wire w5572
// ERROR: floating wire w5644
// ERROR: floating wire w5656
// ERROR: floating wire w5711
// ERROR: floating wire w5765
// ERROR: floating wire w5910
// ERROR: floating wire w5912
// ERROR: floating wire w5925
// ERROR: floating wire w5964
// ERROR: floating wire w5995
// ERROR: floating wire w6012
// ERROR: floating wire w6156
// ERROR: floating wire w6172
// ERROR: floating wire w6203
// ERROR: floating wire w6249
// ERROR: floating wire w6295
// ERROR: floating wire w6296
// ERROR: floating wire w6604
// ERROR: floating wire w6719
// ERROR: floating wire w6721
// ERROR: floating wire w6722
// WARNING: Cell vdp_fa:g385 port CO not connected.
// WARNING: Cell vdp_and:g527 port Z not connected.
// WARNING: Cell vdp_cnt_bit_load:g871 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g873 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g1405 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g1406 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1407 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1408 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1409 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1410 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1411 port Q not connected.
// WARNING: Cell vdp_cnt_bit_load:g1412 port Q not connected.
// WARNING: Cell vdp_or:g1576 port Z not connected.
// WARNING: Cell vdp_cnt_bit_load:g1959 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g1960 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2145 port CO not connected.
// WARNING: Cell vdp_ha:g2278 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2280 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2282 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2284 port CO not connected.
// WARNING: Cell vdp_cnt_bit:g2286 port CO not connected.
// WARNING: Cell vdp_rs_ff:g2380 port nQ not connected.
// WARNING: Cell vdp_rs_ff:g2381 port nQ not connected.
// WARNING: Cell vdp_comp_we:g2612 port nZ not connected.
// WARNING: Cell vdp_fa:g3842 port CO not connected.
// WARNING: Cell vdp_fa:g4058 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g4437 port CO not connected.
// WARNING: Cell vdp_fa:g4453 port CO not connected.
// WARNING: Cell vdp_fa:g4463 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g5851 port CO not connected.
// WARNING: Cell vdp_fa:g5862 port CO not connected.
// WARNING: Cell vdp_fa:g5888 port CO not connected.
// WARNING: Cell vdp_fa:g5892 port CO not connected.
// WARNING: Cell vdp_fa:g6086 port CO not connected.
// WARNING: Cell vdp_ha:g6137 port CO not connected.
// WARNING: Cell vdp_sr_bit:g6146 port Q not connected.
// WARNING: Cell vdp_fa:g6150 port CO not connected.
// WARNING: Cell vdp_cnt_bit_load:g6216 port CO not connected.
