module IO (  VD15_i, VD15_d, VD15_o, VA1_i, VA1_d, VA1_o, VA2_i, VA2_d, VA2_o, VA3_i, VA3_d, VA3_o, VA4_i, VA4_d, VA4_o, VA5_i, VA5_d, VA5_o, VA6_i, VA6_d, VA6_o, VA7_i, VA7_d, VA7_o, n_FRES, n_DISK, PC0_i, PC0_d, PC0_o, PC1_i, PC1_d, PC1_o, PC2_i, PC2_d, PC2_o, PC3_i, PC3_d, PC3_o, PC4_i, PC4_d, PC4_o, PC5_i, PC5_d, PC5_o, PC6_i, PC6_d, PC6_o, TEST, n_HL, n_LWR, n_CAS0, VCLK, n_JAP, NTSC, n_M3, n_IO, n_SRES, n_ZTOV, n_VTOZ, ZD7_i, ZD7_d, ZD7_o, ZD6_i, ZD6_d, ZD6_o, ZD5_i, ZD5_d, ZD5_o, ZD4_i, ZD4_d, ZD4_o, ZD3_i, ZD3_d, ZD3_o, ZD2_i, ZD2_d, ZD2_o, ZD1_i, ZD1_d, ZD1_o, ZD0_i, ZD0_d, ZD0_o, ZA0, ZA1_i, ZA1_d, ZA1_o, ZA2_i, ZA2_d, ZA2_o, ZA3_i, ZA3_d, ZA3_o, ZA4_i, ZA4_d, ZA4_o, ZA5_i, ZA5_d, ZA5_o, ZA6_i, ZA6_d, ZA6_o, ZA7_i, ZA7_d, ZA7_o, PA0_i, PA0_d, PA0_o, PA1_i, PA1_d, PA1_o, PA2_i, PA2_d, PA2_o, PA3_i, PA3_d, PA3_o, PA4_i, PA4_d, PA4_o, PA5_i, PA5_d, PA5_o, PA6_i, PA6_d, PA6_o, PB0_i, PB0_d, PB0_o, PB1_i, PB1_d, PB1_o, PB2_i, PB2_d, PB2_o, PB3_i, PB3_d, PB3_o, PB4_i, PB4_d, PB4_o, PB5_i, PB5_d, PB5_o, PB6_i, PB6_d, PB6_o, VD0_i, VD0_d, VD0_o, VD1_i, VD1_d, VD1_o, VD2_i, VD2_d, VD2_o, VD3_i, VD3_d, VD3_o, VD4_i, VD4_d, VD4_o, VD5_i, VD5_d, VD5_o, VD6_i, VD6_d, VD6_o, VD7_i, VD7_d, VD7_o, VD8_i, VD8_d, VD8_o, VD9_i, VD9_d, VD9_o, VD10_i, VD10_d, VD10_o, VD11_i, VD11_d, VD11_o, VD12_i, VD12_d, VD12_o, VD13_i, VD13_d, VD13_o, VD14_i, VD14_d, VD14_o);

	input wire VD15_i;
	output wire VD15_d;
	output wire VD15_o;
	input wire VA1_i;
	output wire VA1_d;
	output wire VA1_o;
	input wire VA2_i;
	output wire VA2_d;
	output wire VA2_o;
	input wire VA3_i;
	output wire VA3_d;
	output wire VA3_o;
	input wire VA4_i;
	output wire VA4_d;
	output wire VA4_o;
	input wire VA5_i;
	output wire VA5_d;
	output wire VA5_o;
	input wire VA6_i;
	output wire VA6_d;
	output wire VA6_o;
	input wire VA7_i;
	output wire VA7_d;
	output wire VA7_o;
	output wire n_FRES;
	input wire n_DISK;
	input wire PC0_i;
	output wire PC0_d;
	output wire PC0_o;
	input wire PC1_i;
	output wire PC1_d;
	output wire PC1_o;
	input wire PC2_i;
	output wire PC2_d;
	output wire PC2_o;
	input wire PC3_i;
	output wire PC3_d;
	output wire PC3_o;
	input wire PC4_i;
	output wire PC4_d;
	output wire PC4_o;
	input wire PC5_i;
	output wire PC5_d;
	output wire PC5_o;
	input wire PC6_i;
	output wire PC6_d;
	output wire PC6_o;
	input wire TEST;
	output wire n_HL;
	input wire n_LWR;
	input wire n_CAS0;
	input wire VCLK;
	input wire n_JAP;
	input wire NTSC;
	input wire n_M3;
	input wire n_IO;
	input wire n_SRES;
	input wire n_ZTOV;
	input wire n_VTOZ;
	input wire ZD7_i;
	output wire ZD7_d;
	output wire ZD7_o;
	input wire ZD6_i;
	output wire ZD6_d;
	output wire ZD6_o;
	input wire ZD5_i;
	output wire ZD5_d;
	output wire ZD5_o;
	input wire ZD4_i;
	output wire ZD4_d;
	output wire ZD4_o;
	input wire ZD3_i;
	output wire ZD3_d;
	output wire ZD3_o;
	input wire ZD2_i;
	output wire ZD2_d;
	output wire ZD2_o;
	input wire ZD1_i;
	output wire ZD1_d;
	output wire ZD1_o;
	input wire ZD0_i;
	output wire ZD0_d;
	output wire ZD0_o;
	input wire ZA0;
	input wire ZA1_i;
	output wire ZA1_d;
	output wire ZA1_o;
	input wire ZA2_i;
	output wire ZA2_d;
	output wire ZA2_o;
	input wire ZA3_i;
	output wire ZA3_d;
	output wire ZA3_o;
	input wire ZA4_i;
	output wire ZA4_d;
	output wire ZA4_o;
	input wire ZA5_i;
	output wire ZA5_d;
	output wire ZA5_o;
	input wire ZA6_i;
	output wire ZA6_d;
	output wire ZA6_o;
	input wire ZA7_i;
	output wire ZA7_d;
	output wire ZA7_o;
	input wire PA0_i;
	output wire PA0_d;
	output wire PA0_o;
	input wire PA1_i;
	output wire PA1_d;
	output wire PA1_o;
	input wire PA2_i;
	output wire PA2_d;
	output wire PA2_o;
	input wire PA3_i;
	output wire PA3_d;
	output wire PA3_o;
	input wire PA4_i;
	output wire PA4_d;
	output wire PA4_o;
	input wire PA5_i;
	output wire PA5_d;
	output wire PA5_o;
	input wire PA6_i;
	output wire PA6_d;
	output wire PA6_o;
	input wire PB0_i;
	output wire PB0_d;
	output wire PB0_o;
	input wire PB1_i;
	output wire PB1_d;
	output wire PB1_o;
	input wire PB2_i;
	output wire PB2_d;
	output wire PB2_o;
	input wire PB3_i;
	output wire PB3_d;
	output wire PB3_o;
	input wire PB4_i;
	output wire PB4_d;
	output wire PB4_o;
	input wire PB5_i;
	output wire PB5_d;
	output wire PB5_o;
	input wire PB6_i;
	output wire PB6_d;
	output wire PB6_o;
	input wire VD0_i;
	output wire VD0_d;
	output wire VD0_o;
	input wire VD1_i;
	output wire VD1_d;
	output wire VD1_o;
	input wire VD2_i;
	output wire VD2_d;
	output wire VD2_o;
	input wire VD3_i;
	output wire VD3_d;
	output wire VD3_o;
	input wire VD4_i;
	output wire VD4_d;
	output wire VD4_o;
	input wire VD5_i;
	output wire VD5_d;
	output wire VD5_o;
	input wire VD6_i;
	output wire VD6_d;
	output wire VD6_o;
	input wire VD7_i;
	output wire VD7_d;
	output wire VD7_o;
	input wire VD8_i;
	output wire VD8_d;
	output wire VD8_o;
	input wire VD9_i;
	output wire VD9_d;
	output wire VD9_o;
	input wire VD10_i;
	output wire VD10_d;
	output wire VD10_o;
	input wire VD11_i;
	output wire VD11_d;
	output wire VD11_o;
	input wire VD12_i;
	output wire VD12_d;
	output wire VD12_o;
	input wire VD13_i;
	output wire VD13_d;
	output wire VD13_o;
	input wire VD14_i;
	output wire VD14_d;
	output wire VD14_o;

	// Wires

	wire w1;
	wire w2;
	wire w3;
	wire w4;
	wire w5;
	wire w6;
	wire w7;
	wire w8;
	wire w9;
	wire w10;
	wire w11;
	wire w12;
	wire w13;
	wire w14;
	wire w15;
	wire w16;
	wire w17;
	wire w18;
	wire w19;
	wire w20;
	wire w21;
	wire w22;
	wire w23;
	wire w24;
	wire w25;
	wire w26;
	wire w27;
	wire w28;
	wire w29;
	wire w30;
	wire w31;
	wire w32;
	wire w33;
	wire w34;
	wire w35;
	wire w36;
	wire w37;
	wire w38;
	wire w39;
	wire w40;
	wire w41;
	wire w42;
	wire w43;
	wire w44;
	wire w45;
	wire w46;
	wire w47;
	wire w48;
	wire w49;
	wire w50;
	wire w51;
	wire w52;
	wire w53;
	wire w54;
	wire w55;
	wire w56;
	wire w57;
	wire w58;
	wire w59;
	wire w60;
	wire w61;
	wire w62;
	wire w63;
	wire w64;
	wire w65;
	wire w66;
	wire w67;
	wire w68;
	wire w69;
	wire w70;
	wire w71;
	wire w72;
	wire w73;
	wire w74;
	wire w75;
	wire w76;
	wire w77;
	wire w78;
	wire w79;
	wire w80;
	wire w81;
	wire w82;
	wire w83;
	wire w84;
	wire w85;
	wire w86;
	wire w87;
	wire w88;
	wire w89;
	wire w90;
	wire w91;
	wire w92;
	wire w93;
	wire w94;
	wire w95;
	wire w96;
	wire w97;
	wire w98;
	wire w99;
	wire w100;
	wire w101;
	wire w102;
	wire w103;
	wire w104;
	wire w105;
	wire w106;
	wire w107;
	wire w108;
	wire w109;
	wire w110;
	wire w111;
	wire w112;
	wire w113;
	wire w114;
	wire w115;
	wire w116;
	wire w117;
	wire w118;
	wire w119;
	wire w120;
	wire w121;
	wire w122;
	wire w123;
	wire w124;
	wire w125;
	wire w126;
	wire w127;
	wire w128;
	wire w129;
	wire w130;
	wire w131;
	wire w132;
	wire w133;
	wire w134;
	wire w135;
	wire w136;
	wire w137;
	wire w138;
	wire w139;
	wire w140;
	wire w141;
	wire w142;
	wire w143;
	wire w144;
	wire w145;
	wire w146;
	wire w147;
	wire w148;
	wire w149;
	wire w150;
	wire w151;
	wire w152;
	wire w153;
	wire w154;
	wire w155;
	wire w156;
	wire w157;
	wire w158;
	wire w159;
	wire w160;
	wire w161;
	wire w162;
	wire w163;
	wire w164;
	wire w165;
	wire w166;
	wire w167;
	wire w168;
	wire w169;
	wire w170;
	wire w171;
	wire w172;
	wire w173;
	wire w174;
	wire w175;
	wire w176;
	wire w177;
	wire w178;
	wire w179;
	wire w180;
	wire w181;
	wire w182;
	wire w183;
	wire w184;
	wire w185;
	wire w186;
	wire w187;
	wire w188;
	wire w189;
	wire w190;
	wire w191;
	wire w192;
	wire w193;
	wire w194;
	wire w195;
	wire w196;
	wire w197;
	wire w198;
	wire w199;
	wire w200;
	wire w201;
	wire w202;
	wire w203;
	wire w204;
	wire w205;
	wire w206;
	wire w207;
	wire w208;
	wire w209;
	wire w210;
	wire w211;
	wire w212;
	wire w213;
	wire w214;
	wire w215;
	wire w216;
	wire w217;
	wire w218;
	wire w219;
	wire w220;
	wire w221;
	wire w222;
	wire w223;
	wire w224;
	wire w225;
	wire w226;
	wire w227;
	wire w228;
	wire w229;
	wire w230;
	wire w231;
	wire w232;
	wire w233;
	wire w234;
	wire w235;
	wire w236;
	wire w237;
	wire w238;
	wire w239;
	wire w240;
	wire w241;
	wire w242;
	wire w243;
	wire w244;
	wire w245;
	wire w246;
	wire w247;
	wire w248;
	wire w249;
	wire w250;
	wire w251;
	wire w252;
	wire w253;
	wire w254;
	wire w255;
	wire w256;
	wire w257;
	wire w258;
	wire w259;
	wire w260;
	wire w261;
	wire w262;
	wire w263;
	wire w264;
	wire w265;
	wire w266;
	wire w267;
	wire w268;
	wire w269;
	wire w270;
	wire w271;
	wire w272;
	wire w273;
	wire w274;
	wire w275;
	wire w276;
	wire w277;
	wire w278;
	wire w279;
	wire w280;
	wire w281;
	wire w282;
	wire w283;
	wire w284;
	wire w285;
	wire w286;
	wire w287;
	wire w288;
	wire w289;
	wire w290;
	wire w291;
	wire w292;
	wire w293;
	wire w294;
	wire w295;
	wire w296;
	wire w297;
	wire w298;
	wire w299;
	wire w300;
	wire w301;
	wire w302;
	wire w303;
	wire w304;
	wire w305;
	wire w306;
	wire w307;
	wire w308;
	wire w309;
	wire w310;
	wire w311;
	wire w312;
	wire w313;
	wire w314;
	wire w315;
	wire w316;
	wire w317;
	wire w318;
	wire w319;
	wire w320;
	wire w321;
	wire w322;
	wire w323;
	wire w324;
	wire w325;
	wire w326;
	wire w327;
	wire w328;
	wire w329;
	wire w330;
	wire w331;
	wire w332;
	wire w333;
	wire w334;
	wire w335;
	wire w336;
	wire w337;
	wire w338;
	wire w339;
	wire w340;
	wire w341;
	wire w342;
	wire w343;
	wire w344;
	wire w345;
	wire w346;
	wire w347;
	wire w348;
	wire w349;
	wire w350;
	wire w351;
	wire w352;
	wire w353;
	wire w354;
	wire w355;
	wire w356;
	wire w357;
	wire w358;
	wire w359;
	wire w360;
	wire w361;
	wire w362;
	wire w363;
	wire w364;
	wire w365;
	wire w366;
	wire w367;
	wire w368;
	wire w369;
	wire w370;
	wire w371;
	wire w372;
	wire w373;
	wire w374;
	wire w375;
	wire w376;
	wire w377;
	wire w378;
	wire w379;
	wire w380;
	wire w381;
	wire w382;
	wire w383;
	wire w384;
	wire w385;
	wire w386;
	wire w387;
	wire w388;
	wire w389;
	wire w390;
	wire w391;
	wire w392;
	wire w393;
	wire w394;
	wire w395;
	wire w396;
	wire w397;
	wire w398;
	wire w399;
	wire w400;
	wire w401;
	wire w402;
	wire w403;
	wire w404;
	wire w405;
	wire w406;
	wire w407;
	wire w408;
	wire w409;
	wire w410;
	wire w411;
	wire w412;
	wire w413;
	wire w414;
	wire w415;
	wire w416;
	wire w417;
	wire w418;
	wire w419;
	wire w420;
	wire w421;
	wire w422;
	wire w423;
	wire w424;
	wire w425;
	wire w426;
	wire w427;
	wire w428;
	wire w429;
	wire w430;
	wire w431;
	wire w432;
	wire w433;
	wire w434;
	wire w435;
	wire w436;
	wire w437;
	wire w438;
	wire w439;
	wire w440;
	wire w441;
	wire w442;
	wire w443;
	wire w444;
	wire w445;
	wire w446;
	wire w447;
	wire w448;
	wire w449;
	wire w450;
	wire w451;
	wire w452;
	wire w453;
	wire w454;
	wire w455;
	wire w456;
	wire w457;
	wire w458;
	wire w459;
	wire w460;
	wire w461;
	wire w462;
	wire w463;
	wire w464;
	wire w465;
	wire w466;
	wire w467;
	wire w468;
	wire w469;
	wire w470;
	wire w471;
	wire w472;
	wire w473;
	wire w474;
	wire w475;
	wire w476;
	wire w477;
	wire w478;
	wire w479;
	wire w480;
	wire w481;
	wire w482;
	wire w483;
	wire w484;
	wire w485;
	wire w486;
	wire w487;
	wire w488;
	wire w489;
	wire w490;
	wire w491;
	wire w492;
	wire w493;
	wire w494;
	wire w495;
	wire w496;
	wire w497;
	wire w498;
	wire w499;
	wire w500;
	wire w501;
	wire w502;
	wire w503;
	wire w504;
	wire w505;
	wire w506;
	wire w507;
	wire w508;
	wire w509;
	wire w510;
	wire w511;
	wire w512;
	wire w513;
	wire w514;
	wire w515;
	wire w516;
	wire w517;
	wire w518;
	wire w519;
	wire w520;
	wire w521;
	wire w522;
	wire w523;
	wire w524;
	wire w525;
	wire w526;
	wire w527;
	wire w528;
	wire w529;
	wire w530;
	wire w531;
	wire w532;
	wire w533;
	wire w534;
	wire w535;
	wire w536;
	wire w537;
	wire w538;
	wire w539;
	wire w540;
	wire w541;
	wire w542;
	wire w543;
	wire w544;
	wire w545;
	wire w546;
	wire w547;
	wire w548;
	wire w549;
	wire w550;
	wire w551;
	wire w552;
	wire w553;
	wire w554;
	wire w555;
	wire w556;
	wire w557;
	wire w558;
	wire w559;
	wire w560;
	wire w561;
	wire w562;
	wire w563;
	wire w564;
	wire w565;
	wire w566;
	wire w567;
	wire w568;
	wire w569;
	wire w570;
	wire w571;
	wire w572;
	wire w573;
	wire w574;
	wire w575;
	wire w576;
	wire w577;
	wire w578;
	wire w579;
	wire w580;
	wire w581;
	wire w582;
	wire w583;
	wire w584;
	wire w585;
	wire w586;
	wire w587;
	wire w588;
	wire w589;
	wire w590;
	wire w591;
	wire w592;
	wire w593;
	wire w594;
	wire w595;
	wire w596;
	wire w597;
	wire w598;
	wire w599;
	wire w600;
	wire w601;
	wire w602;
	wire w603;
	wire w604;
	wire w605;
	wire w606;
	wire w607;
	wire w608;
	wire w609;
	wire w610;
	wire w611;
	wire w612;
	wire w613;
	wire w614;
	wire w615;
	wire w616;
	wire w617;
	wire w618;
	wire w619;
	wire w620;
	wire w621;
	wire w622;
	wire w623;
	wire w624;
	wire w625;
	wire w626;
	wire w627;
	wire w628;
	wire w629;
	wire w630;
	wire w631;
	wire w632;
	wire w633;
	wire w634;
	wire w635;
	wire w636;
	wire w637;
	wire w638;
	wire w639;
	wire w640;
	wire w641;
	wire w642;
	wire w643;
	wire w644;
	wire w645;
	wire w646;
	wire w647;
	wire w648;
	wire w649;
	wire w650;
	wire w651;
	wire w652;
	wire w653;
	wire w654;
	wire w655;
	wire w656;
	wire w657;
	wire w658;
	wire w659;
	wire w660;
	wire w661;
	wire w662;
	wire w663;
	wire w664;
	wire w665;
	wire w666;
	wire w667;
	wire w668;
	wire w669;
	wire w670;
	wire w671;
	wire w672;
	wire w673;
	wire w674;
	wire w675;
	wire w676;
	wire w677;
	wire w678;
	wire w679;
	wire w680;
	wire w681;
	wire w682;
	wire w683;
	wire w684;
	wire w685;
	wire w686;
	wire w687;
	wire w688;
	wire w689;
	wire w690;
	wire w691;
	wire w692;
	wire w693;
	wire w694;
	wire w695;
	wire w696;
	wire w697;
	wire w698;
	wire w699;
	wire w700;
	wire w701;
	wire w702;
	wire w703;
	wire w704;
	wire w705;
	wire w706;
	wire w707;
	wire w708;
	wire w709;
	wire w710;
	wire w711;
	wire w712;
	wire w713;
	wire w714;
	wire w715;
	wire w716;
	wire w717;
	wire w718;
	wire w719;
	wire w720;
	wire w721;
	wire w722;
	wire w723;
	wire w724;
	wire w725;
	wire w726;
	wire w727;
	wire w728;
	wire w729;
	wire w730;
	wire w731;
	wire w732;
	wire w733;
	wire w734;
	wire w735;
	wire w736;
	wire w737;
	wire w738;
	wire w739;
	wire w740;
	wire w741;
	wire w742;
	wire w743;
	wire w744;
	wire w745;
	wire w746;
	wire w747;
	wire w748;
	wire w749;
	wire w750;
	wire w751;
	wire w752;
	wire w753;
	wire w754;
	wire w755;
	wire w756;
	wire w757;
	wire w758;
	wire w759;
	wire w760;
	wire w761;
	wire w762;
	wire w763;
	wire w764;
	wire w765;
	wire w766;
	wire w767;
	wire w768;
	wire w769;
	wire w770;
	wire w771;
	wire w772;
	wire w773;
	wire w774;
	wire w775;
	wire w776;
	wire w777;
	wire w778;
	wire w779;
	wire w780;
	wire w781;
	wire w782;
	wire w783;
	wire w784;
	wire w785;
	wire w786;
	wire w787;
	wire w788;
	wire w789;
	wire w790;
	wire w791;
	wire w792;
	wire w793;
	wire w794;
	wire w795;
	wire w796;
	wire w797;
	wire w798;
	wire w799;
	wire w800;
	wire w801;
	wire w802;
	wire w803;
	wire w804;
	wire w805;
	wire w806;
	wire w807;
	wire w808;
	wire w809;
	wire w810;
	wire w811;
	wire w812;
	wire w813;
	wire w814;
	wire w815;
	wire w816;
	wire w817;
	wire w818;
	wire w819;
	wire w820;
	wire w821;
	wire w822;
	wire w823;
	wire w824;
	wire w825;
	wire w826;
	wire w827;
	wire w828;
	wire w829;
	wire w830;
	wire w831;
	wire w832;
	wire w833;
	wire w834;
	wire w835;
	wire w836;
	wire w837;
	wire w838;
	wire w839;
	wire w840;
	wire w841;
	wire w842;
	wire w843;
	wire w844;
	wire w845;
	wire w846;
	wire w847;
	wire w848;
	wire w849;
	wire w850;
	wire w851;
	wire w852;
	wire w853;
	wire w854;
	wire w855;
	wire w856;
	wire w857;
	wire w858;
	wire w859;
	wire w860;
	wire w861;
	wire w862;
	wire w863;
	wire w864;
	wire w865;
	wire w866;
	wire w867;
	wire w868;
	wire w869;
	wire w870;
	wire w871;
	wire w872;
	wire w873;
	wire w874;
	wire w875;
	wire w876;
	wire w877;
	wire w878;
	wire w879;
	wire w880;
	wire w881;
	wire w882;
	wire w883;
	wire w884;
	wire w885;
	wire w886;
	wire w887;
	wire w888;
	wire w889;
	wire w890;
	wire w891;
	wire w892;
	wire w893;
	wire w894;
	wire w895;
	wire w896;
	wire w897;
	wire w898;
	wire w899;
	wire w900;
	wire w901;
	wire w902;
	wire w903;
	wire w904;
	wire w905;
	wire w906;
	wire w907;
	wire w908;
	wire w909;
	wire w910;
	wire w911;
	wire w912;
	wire w913;
	wire w914;
	wire w915;
	wire w916;
	wire w917;
	wire w918;
	wire w919;
	wire w920;
	wire w921;
	wire w922;
	wire w923;
	wire w924;
	wire w925;
	wire w926;
	wire w927;
	wire w928;
	wire w929;
	wire w930;
	wire w931;
	wire w932;
	wire w933;
	wire w934;

	assign w217 = VD15_i;
	assign VD15_d = w208;
	assign VD15_o = w205;
	assign w57 = VA1_i;
	assign VA1_d = w291;
	assign VA1_o = w224;
	assign w54 = VA2_i;
	assign VA2_d = w291;
	assign VA2_o = w223;
	assign w66 = VA3_i;
	assign VA3_d = w291;
	assign VA3_o = w55;
	assign w102 = VA4_i;
	assign VA4_d = w291;
	assign VA4_o = w222;
	assign w103 = VA5_i;
	assign VA5_d = w291;
	assign VA5_o = w88;
	assign w104 = VA6_i;
	assign VA6_d = w291;
	assign VA6_o = w246;
	assign w106 = VA7_i;
	assign VA7_d = w291;
	assign VA7_o = w259;
	assign n_FRES = w300;
	assign w306 = n_DISK;
	assign w307 = PC0_i;
	assign PC0_d = w308;
	assign PC0_o = w330;
	assign w157 = PC1_i;
	assign PC1_d = w310;
	assign PC1_o = w309;
	assign w257 = PC2_i;
	assign PC2_d = w331;
	assign PC2_o = w311;
	assign w314 = PC3_i;
	assign PC3_d = w313;
	assign PC3_o = w312;
	assign w317 = PC4_i;
	assign PC4_d = w316;
	assign PC4_o = w315;
	assign w318 = PC5_i;
	assign PC5_d = w319;
	assign PC5_o = w320;
	assign w321 = PC6_i;
	assign PC6_d = w322;
	assign PC6_o = w323;
	assign w324 = TEST;
	assign n_HL = w245;
	assign w325 = n_LWR;
	assign w268 = n_CAS0;
	assign w115 = VCLK;
	assign w153 = n_JAP;
	assign w293 = NTSC;
	assign w8 = n_M3;
	assign w266 = n_IO;
	assign w292 = n_SRES;
	assign w291 = n_ZTOV;
	assign w98 = n_VTOZ;
	assign w289 = ZD7_i;
	assign ZD7_d = w232;
	assign ZD7_o = w290;
	assign w288 = ZD6_i;
	assign ZD6_d = w232;
	assign ZD6_o = w287;
	assign w286 = ZD5_i;
	assign ZD5_d = w232;
	assign ZD5_o = w285;
	assign w283 = ZD4_i;
	assign ZD4_d = w232;
	assign ZD4_o = w284;
	assign w229 = ZD3_i;
	assign ZD3_d = w232;
	assign ZD3_o = w278;
	assign w280 = ZD2_i;
	assign ZD2_d = w232;
	assign ZD2_o = w279;
	assign w228 = ZD1_i;
	assign ZD1_d = w232;
	assign ZD1_o = w281;
	assign w226 = ZD0_i;
	assign ZD0_d = w232;
	assign ZD0_o = w282;
	assign w188 = ZA0;
	assign w35 = ZA1_i;
	assign ZA1_d = w98;
	assign ZA1_o = w57;
	assign w99 = ZA2_i;
	assign ZA2_d = w98;
	assign ZA2_o = w54;
	assign w100 = ZA3_i;
	assign ZA3_d = w98;
	assign ZA3_o = w66;
	assign w101 = ZA4_i;
	assign ZA4_d = w98;
	assign ZA4_o = w102;
	assign w90 = ZA5_i;
	assign ZA5_d = w98;
	assign ZA5_o = w103;
	assign w91 = ZA6_i;
	assign ZA6_d = w98;
	assign ZA6_o = w104;
	assign w105 = ZA7_i;
	assign ZA7_d = w98;
	assign ZA7_o = w106;
	assign w107 = PA0_i;
	assign PA0_d = w84;
	assign PA0_o = w85;
	assign w160 = PA1_i;
	assign PA1_d = w79;
	assign PA1_o = w932;
	assign w258 = PA2_i;
	assign PA2_d = w80;
	assign PA2_o = w81;
	assign w76 = PA3_i;
	assign PA3_d = w83;
	assign PA3_o = w82;
	assign w73 = PA4_i;
	assign PA4_d = w155;
	assign PA4_o = w74;
	assign w71 = PA5_i;
	assign PA5_d = w72;
	assign PA5_o = w75;
	assign w70 = PA6_i;
	assign PA6_d = w69;
	assign PA6_o = w68;
	assign w65 = PB0_i;
	assign PB0_d = w64;
	assign PB0_o = w67;
	assign w63 = PB1_i;
	assign PB1_d = w62;
	assign PB1_o = w58;
	assign w61 = PB2_i;
	assign PB2_d = w60;
	assign PB2_o = w59;
	assign w28 = PB3_i;
	assign PB3_d = w26;
	assign PB3_o = w27;
	assign w242 = PB4_i;
	assign PB4_d = w13;
	assign PB4_o = w15;
	assign w23 = PB5_i;
	assign PB5_d = w25;
	assign PB5_o = w24;
	assign w189 = PB6_i;
	assign PB6_d = w96;
	assign PB6_o = w190;
	assign w191 = VD0_i;
	assign VD0_d = w192;
	assign VD0_o = w193;
	assign w195 = VD1_i;
	assign VD1_d = w192;
	assign VD1_o = w194;
	assign w197 = VD2_i;
	assign VD2_d = w192;
	assign VD2_o = w196;
	assign w198 = VD3_i;
	assign VD3_d = w192;
	assign VD3_o = w213;
	assign w199 = VD4_i;
	assign VD4_d = w192;
	assign VD4_o = w200;
	assign w202 = VD5_i;
	assign VD5_d = w192;
	assign VD5_o = w201;
	assign w204 = VD6_i;
	assign VD6_d = w192;
	assign VD6_o = w203;
	assign w206 = VD7_i;
	assign VD7_d = w192;
	assign VD7_o = w205;
	assign w209 = VD8_i;
	assign VD8_d = w208;
	assign VD8_o = w207;
	assign w210 = VD9_i;
	assign VD9_d = w208;
	assign VD9_o = w194;
	assign w211 = VD10_i;
	assign VD10_d = w208;
	assign VD10_o = w196;
	assign w212 = VD11_i;
	assign VD11_d = w208;
	assign VD11_o = w213;
	assign w214 = VD12_i;
	assign VD12_d = w208;
	assign VD12_o = w200;
	assign w215 = VD13_i;
	assign VD13_d = w208;
	assign VD13_o = w201;
	assign w216 = VD14_i;
	assign VD14_d = w208;
	assign VD14_o = w203;

	// Instances

	io_AND g_1 (.Z(w1), .B(w2), .A(w8) );
	io_OR g_2 (.A(w1), .Z(w129), .B(w10) );
	io_NOR g_3 (.Z(w10), .B(w8), .A(w5) );
	io_NOT g_4 (.A(w9), .nZ(w5) );
	io_OR g_5 (.B(w5), .Z(w12), .A(w6) );
	io_AND g_6 (.Z(w173), .B(w6), .A(w11) );
	io_OR4 g_7 (.Z(w11), .D(w8), .C(w4), .B(w3), .A(w7) );
	io_OR g_8 (.B(w2), .Z(w4), .A(w20) );
	io_OR3 g_9 (.Z(w6), .C(w8), .B(w14), .A(w16) );
	io_NAND g_10 (.A(w161), .B(w930), .Z(w3) );
	io_NOT g_11 (.A(w161), .nZ(w22) );
	io_NOT g_12 (.A(w930), .nZ(w21) );
	io_NAND8 g_13 (.Z(w14), .D(w22), .C(w21), .B(w20), .A(1'b1), .E(w2), .F(w18), .G(w17), .H(w32) );
	io_AND3 g_14 (.Z(w31), .C(w32), .B(w17), .A(w18) );
	io_NOR g_15 (.Z(w7), .B(w31), .A(w30) );
	io_NOR3 g_16 (.Z(w30), .C(w17), .B(w32), .A(w18) );
	io_DFFRPOS g_17 (.Q(w29), .nRES(1'b1), .D(w186), .C(w33) );
	io_DFFRPOS g_18 (.Q(w27), .nRES(1'b1), .D(w156), .C(w33) );
	io_NOT g_19 (.A(w221), .nZ(w26) );
	io_DFFRPOS g_20 (.Q(w59), .nRES(1'b1), .D(w108), .C(w33) );
	io_DFFRPOS g_21 (.Q(w58), .nRES(1'b1), .D(w336), .C(w33) );
	io_NOT g_22 (.A(w120), .nZ(w62) );
	io_MUX4BIT g_23 (.S(w8), .Z0(w32), .A0(w100), .B0(w102), .A1(w99), .B1(w66), .Z1(w17), .Z2(w2), .B2(w54), .A2(w35), .A3(w188), .B3(w57), .Z3(w9) );
	io_NOT g_24 (.A(w166), .nZ(w60) );
	io_NOT g_25 (.A(w134), .nZ(w64) );
	io_DFFRPOS g_26 (.Q(w67), .nRES(1'b1), .D(w143), .C(w33) );
	io_DFFSPOS g_27 (.C(w12), .D(w130), .nSET(w122), .Q(w131) );
	io_MUX4BIT g_28 (.C(w8), .Z0(w190), .A0(w163), .B0(w133), .A1(w131), .B1(w124), .Z1(w24), .Z2(w68), .B2(w126), .A2(w162), .A3(w132), .B3(w123), .Z3(w75) );
	io_DFFSPOS g_29 (.C(w12), .D(w138), .nSET(w122), .Q(w163) );
	io_DFFSPOS g_30 (.C(w12), .D(w165), .nSET(w122), .Q(w162) );
	io_OR g_31 (.B(w153), .Z(w145), .A(w72) );
	io_AND g_32 (.Z(w147), .B(w145), .A(w71) );
	io_OR g_33 (.B(w153), .Z(w929), .A(w25) );
	io_MUX4BIT g_34 (.S(w8), .Z0(w154), .A0(w151), .B0(w28), .A1(w242), .B1(w61), .Z1(w150), .Z2(w149), .B2(w63), .A2(w28), .A3(w61), .B3(w65), .Z3(w152) );
	io_AND g_35 (.Z(w151), .A(w23), .B(w929) );
	io_DFFRPOS g_36 (.Q(w82), .nRES(1'b1), .D(w156), .C(w142) );
	io_NOT g_37 (.A(w77), .nZ(w83) );
	io_DFFRPOS g_38 (.Q(w81), .nRES(1'b1), .D(w108), .C(w142) );
	io_DFFRPOS g_39 (.Q(w85), .nRES(1'b1), .D(w143), .C(w142) );
	io_DFFRPOS g_40 (.Q(w932), .nRES(1'b1), .D(w336), .C(w142) );
	io_NOT g_41 (.A(w249), .nZ(w84) );
	io_DFFRPOS g_42 (.nRES(w112), .D(1'b0), .C(w86) );
	io_MUX4BIT g_43 (.S(w8), .A0(1'b0), .B0(1'b0), .A1(w91), .B1(w105), .Z1(w259), .Z2(w246), .B2(w91), .A2(w90), .A3(w101), .B3(w90), .Z3(w88) );
	io_DFFRPOS g_44 (.nRES(w112), .D(1'b0), .C(w86) );
	io_MUX4BIT g_45 (.S(w8), .Z0(w161), .A0(w105), .B0(1'b0), .A1(w91), .B1(w106), .Z1(w930), .Z2(w20), .B2(w104), .A2(w90), .A3(w101), .B3(w103), .Z3(w18) );
	io_NOR4 g_46 (.Z(w174), .D(w161), .C(w930), .B(w20), .A(w18) );
	io_DFFRPOS g_47 (.Q(w50), .nRES(w112), .D(w186), .C(w176) );
	io_DFFRPOS g_48 (.Q(w184), .nRES(w112), .D(w186), .C(w86) );
	io_DFFRPOS g_49 (.nRES(w112), .D(1'b0), .C(w176) );
	io_DFFRPOS g_50 (.nRES(w112), .D(1'b0), .C(w176) );
	io_DFFRPOS g_51 (.nRES(w112), .D(1'b0), .C(w137) );
	io_DFFRPOS g_52 (.nRES(w112), .D(1'b0), .C(w137) );
	io_DFFRPOS g_53 (.nRES(w112), .D(1'b0), .C(w137) );
	io_NAND4 g_54 (.B(w92), .C(w175), .A(w93), .D(w170) );
	io_NAND4 g_55 (.B(w94), .C(w93), .A(w92), .D(w170), .Z(w860) );
	io_NOT g_56 (.A(w2), .nZ(w168) );
	io_NAND4 g_57 (.B(w94), .C(w170), .A(w93), .D(w168) );
	io_NOT g_58 (.A(w170), .nZ(w95) );
	io_NAND4 g_59 (.B(w95), .C(w168), .A(w94), .D(w93) );
	io_NOT g_60 (.A(w175), .nZ(w94) );
	io_NAND4 g_61 (.B(w92), .C(w93), .A(w95), .D(w94) );
	io_NAND4 g_62 (.B(w95), .C(w175), .A(w92), .D(w93), .Z(w167) );
	io_NAND4 g_63 (.B(w95), .C(w175), .A(w93), .D(w168) );
	io_NOT g_64 (.A(w168), .nZ(w92) );
	io_NOT g_65 (.A(w96), .nZ(w46) );
	io_NOT g_66 (.A(w69), .nZ(w97) );
	io_AND3 g_67 (.Z(w192), .C(w237), .B(w236), .A(w879) );
	io_OR g_68 (.B(w291), .Z(w879), .A(w235) );
	io_NOT g_69 (.A(w268), .nZ(w235) );
	io_OR g_70 (.B(w268), .Z(w236), .A(w98) );
	io_OR g_71 (.B(w235), .Z(w234), .A(w98) );
	io_AND g_72 (.Z(w232), .B(w233), .A(w234) );
	io_OR g_73 (.B(w291), .Z(w233), .A(w268) );
	io_MUX4BIT g_74 (.S(w227), .Z0(w893), .A0(w198), .B0(w212), .A1(w197), .B1(w211), .Z1(w231), .Z2(w238), .B2(w210), .A2(w195), .A3(w191), .B3(w209), .Z3(w886) );
	io_NOT g_75 (.A(w814), .nZ(w931) );
	io_MUX4BIT g_76 (.S(w752), .Z0(w156), .A0(w198), .B0(w229), .A1(w197), .B1(w280), .Z1(w108), .Z2(w336), .B2(w228), .A2(w195), .A3(w191), .B3(w226), .Z3(w143) );
	io_MUX4BIT g_77 (.S(w53), .Z0(w213), .A0(w229), .B0(w902), .A1(w280), .B1(w901), .Z1(w196), .Z2(w194), .B2(w928), .A2(w228), .A3(w226), .B3(w225), .Z3(w193) );
	io_CNT_BIT g_78 (.nQ(w887), .C(w115), .nRES(1'b1), .D(1'b1), .nLD(w119), .CI(w218) );
	io_NOR4 g_79 (.Z(w394), .D(w887), .C(w910), .B(w888), .A(w889) );
	io_CNT_BIT g_80 (.nQ(w888), .C(w115), .nRES(1'b1), .D(1'b0), .nLD(w119), .CO(w890), .CI(w219) );
	io_CNT_BIT g_81 (.Q(w876), .nQ(w910), .C(w115), .nRES(1'b1), .D(1'b0), .nLD(w119), .CO(w218), .CI(w890) );
	io_DFFRPOS g_82 (.Q(w134), .nRES(w112), .D(w143), .C(w853) );
	io_DFFRPOS g_83 (.Q(w126), .nRES(1'b1), .D(w130), .C(w142) );
	io_DFFRPOS g_84 (.Q(w123), .nRES(1'b1), .D(w165), .C(w142) );
	io_DFFRPOS g_85 (.Q(w124), .nRES(1'b1), .D(w165), .C(w33) );
	io_NOT g_86 (.A(w241), .nZ(w146) );
	io_DFFRPOS g_87 (.Q(w254), .nRES(1'b1), .D(w138), .C(w142) );
	io_MUX4BIT g_88 (.S(w8), .Z0(w796), .A0(w63), .B0(w254), .A1(w65), .B1(w70), .Z1(w760), .Z2(w243), .B2(w71), .A2(w147), .A3(w73), .B3(w73), .Z3(w244) );
	io_MUX8TO1 g_89 (.S0(w250), .S2(w247), .S1(w251), .G(w252), .H(w253), .F(w134), .E(w249), .Z(w892), .C(w152), .D(w307), .B(w107), .A(w891) );
	io_MUX8TO1 g_90 (.S0(w250), .S2(w247), .S1(w251), .G(w255), .H(w248), .F(w221), .E(w77), .Z(w894), .C(w154), .D(w314), .B(w76), .A(w895) );
	io_MUX8TO1 g_91 (.S0(w250), .S2(w247), .S1(w251), .G(w477), .H(w650), .F(w166), .E(w139), .Z(w903), .C(w150), .D(w257), .B(w258), .A(w788) );
	io_DFFSPOS g_92 (.C(w366), .D(w71), .nSET(w276), .nQ(w260), .Q(w556) );
	io_DFFRPOS g_93 (.Q(w904), .nRES(w905), .D(w260), .C(w436) );
	io_MUX8TO1 g_94 (.S0(w250), .S2(w247), .S1(w251), .G(w925), .H(w265), .F(w676), .E(w270), .Z(w899), .C(w878), .D(w262), .B(w269), .A(w264) );
	io_DFFRPOS g_95 (.Q(w265), .nRES(w112), .D(w156), .C(w86) );
	io_NOR3 g_96 (.Z(w53), .C(w268), .B(w266), .A(w267) );
	io_AND g_97 (.Z(w272), .B(1'b1), .A(w556) );
	io_DFFRPOS g_98 (.Q(w839), .nRES(w905), .D(1'b1), .C(w436) );
	io_DFFRPOS g_99 (.Q(w264), .nRES(1'b1), .D(w920), .C(w436) );
	io_DFFRPOS g_100 (.Q(w823), .nRES(1'b1), .D(w908), .C(w436) );
	io_NOT g_101 (.A(w275), .nZ(w182) );
	io_SIPO_4BIT g_102 (.C(w355), .D(w272), .nRES(w276), .Q0(w921), .Q1(w274), .Q2(w850), .Q3(w909) );
	io_SIPO_4BIT g_103 (.C(w355), .D(w909), .nRES(w276), .Q0(w914), .Q1(w916), .Q2(w852), .Q3(w748) );
	io_AND g_104 (.Z(w905), .B(w859), .A(w171) );
	io_DFFRPOS g_105 (.Q(w919), .nRES(1'b1), .D(w915), .C(w436) );
	io_DFFRPOS g_106 (.Q(w838), .nRES(1'b1), .D(w917), .C(w436) );
	io_NOT g_107 (.A(w32), .nZ(w855) );
	io_OR g_108 (.B(w268), .Z(w277), .A(w266) );
	io_NOR g_109 (.Z(w47), .B(w46), .A(w189) );
	io_NOR g_110 (.Z(w48), .B(w49), .A(w47) );
	io_NAND g_111 (.B(w240), .A(w53), .Z(w237) );
	io_NOR g_112 (.Z(w40), .B(w8), .A(w48) );
	io_DFFSPOS g_113 (.C(w230), .D(w52), .nSET(w50), .Q(w45) );
	io_AND g_114 (.Z(w43), .B(w50), .A(w45) );
	io_NOT g_115 (.A(w51), .nZ(w44) );
	io_NOR g_116 (.Z(w239), .B(w189), .A(w44) );
	io_NOT g_117 (.A(w50), .nZ(w42) );
	io_AND g_118 (.Z(w13), .B(w42), .A(w931) );
	io_OR g_119 (.B(w41), .Z(w15), .A(w43) );
	io_AND g_120 (.B(w42), .Z(w41), .A(w29) );
	io_NOT g_121 (.A(w8), .nZ(w38) );
	io_NOR g_122 (.Z(w39), .B(w56), .A(w38) );
	io_NOR g_123 (.Z(w245), .B(w40), .A(w39) );
	io_BUF g_124 (.Z(w240), .A(w8) );
	io_AND g_125 (.Z(w227), .B(w36), .A(w240) );
	io_NOT g_126 (.A(w188), .nZ(w36) );
	io_MUX4BIT g_127 (.S(w8), .Z0(w222), .A0(w100), .B0(w101), .A1(w99), .B1(w100), .Z1(w55), .Z2(w223), .B2(w99), .A2(w35), .A3(w188), .B3(w35), .Z3(w224) );
	io_AND3 g_128 (.Z(w37), .C(1'b1), .B(w119), .A(1'b1) );
	io_CNT_BIT g_129 (.nQ(w109), .C(w115), .nRES(1'b1), .D(w121), .nLD(w119), .CO(w110), .CI(w37) );
	io_CNT_BIT g_130 (.nQ(w113), .C(w115), .nRES(1'b1), .D(1'b0), .nLD(w119), .CO(w111), .CI(w110) );
	io_AND g_131 (.Z(w112), .B(w8), .A(w127) );
	io_NOR4 g_132 (.Z(w523), .D(w113), .C(w109), .B(w117), .A(w116) );
	io_CNT_BIT g_133 (.nQ(w116), .C(w115), .nRES(1'b1), .D(1'b1), .nLD(w119), .CO(w118), .CI(w111) );
	io_CNT_BIT g_134 (.nQ(w117), .C(w115), .nRES(1'b1), .D(1'b1), .nLD(w119), .CI(w118) );
	io_BUF g_135 (.Z(w128), .A(w129) );
	io_BUF g_136 (.Z(w122), .A(w127) );
	io_NOR g_137 (.Z(w49), .B(w70), .A(w97) );
	io_NOT g_138 (.A(w817), .nZ(w164) );
	io_DFFSPOS g_139 (.C(w12), .D(w336), .nSET(w122), .Q(w125) );
	io_DFFSPOS g_140 (.C(w12), .D(w108), .nSET(w122), .Q(w136) );
	io_MUX4BIT g_141 (.S(w8), .Z0(w96), .A0(w135), .B0(w146), .A1(w136), .B1(w180), .Z1(w25), .Z2(w69), .B2(w164), .A2(w125), .A3(w144), .B3(w148), .Z3(w72) );
	io_DFFSPOS g_142 (.C(w12), .D(w143), .nSET(w122), .Q(w144) );
	io_DFFSPOS g_143 (.C(w12), .D(w156), .nSET(w122), .Q(w135) );
	io_BUF g_144 (.Z(w251), .A(w129) );
	io_DFFRPOS g_145 (.Q(w249), .nRES(w112), .D(w143), .C(w140) );
	io_DFFRPOS g_146 (.Q(w77), .nRES(w112), .D(w156), .C(w140) );
	io_MUX8TO1 g_147 (.SO(w250), .S1(w251), .S2(w247), .G(w351), .H(w159), .F(w120), .E(w141), .Z(w158), .C(w149), .D(w157), .B(w160), .A(w256) );
	io_NOT g_148 (.A(w139), .nZ(w80) );
	io_NOT g_149 (.A(w141), .nZ(w79) );
	io_DFFRPOS g_150 (.Q(w139), .nRES(w112), .D(w108), .C(w140) );
	io_DFFRPOS g_151 (.Q(w787), .nRES(w112), .D(w138), .C(w137) );
	io_DFFRPOS g_152 (.Q(w261), .nRES(w112), .D(w186), .C(w137) );
	io_DFFRPOS g_153 (.Q(w141), .nRES(w112), .D(w336), .C(w140) );
	io_DFFRPOS g_154 (.nRES(w112), .D(1'b0), .C(w86) );
	io_DFFRPOS g_155 (.Q(w269), .nRES(w112), .D(w156), .C(w137) );
	io_DFFRPOS g_156 (.Q(w270), .nRES(w112), .D(w156), .C(w176) );
	io_OR g_157 (.A(w178), .Z(w180), .B(w179) );
	io_NOT g_158 (.A(w263), .nZ(w179) );
	io_DFFRPOS g_159 (.Q(w271), .nRES(w112), .D(w165), .C(w86) );
	io_DFFRPOS g_160 (.Q(w275), .nRES(w112), .D(w165), .C(w140) );
	io_OR g_161 (.B(w276), .Z(w148), .A(w182) );
	io_BUF g_162 (.Z(w247), .A(w181) );
	io_BUF g_163 (.Z(w183), .A(w181) );
	io_DFFRPOS g_164 (.nRES(w112), .D(1'b0), .C(w176) );
	io_DFFRPOS g_165 (.Q(w178), .nRES(w112), .D(w165), .C(w176) );
	io_DFFRPOS g_166 (.Q(w276), .nRES(w112), .D(w165), .C(w137) );
	io_AND g_167 (.Z(w181), .B(w17), .A(w8) );
	io_NOT g_168 (.A(w17), .nZ(w170) );
	io_NAND g_169 (.A(w8), .B(w174), .Z(w172) );
	io_AND g_170 (.Z(w267), .B(w173), .A(w172) );
	io_NOT g_171 (.A(w9), .nZ(w175) );
	io_NAND4 g_172 (.B(w175), .C(w170), .A(w168), .D(w93), .Z(w171) );
	io_NOR3 g_173 (.Z(w93), .C(w172), .B(w277), .A(w169) );
	io_NOT g_174 (.A(w32), .nZ(w169) );
	io_AND g_175 (.Z(w52), .B(w589), .A(w880) );
	io_NOT g_176 (.A(w881), .nZ(w880) );
	io_DFFRPOS g_177 (.Q(w881), .nRES(w50), .D(w882), .C(w727) );
	io_AON22 g_178 (.Z(w882), .B2(w731), .A2(w728), .B1(w883), .A1(w874) );
	io_DFFRPOS g_179 (.Q(w883), .nRES(w50), .D(w884), .C(w727) );
	io_NOT g_180 (.A(w728), .Z(w731) );
	io_AON22 g_181 (.Z(w884), .B2(w731), .A2(w728), .B1(w885), .A1(w765) );
	io_DFFRPOS g_182 (.Q(w885), .nRES(w50), .D(w875), .C(w727) );
	io_DFFRPOS g_183 (.Q(w221), .nRES(w112), .D(w156), .C(w853) );
	io_DFFRPOS g_184 (.Q(w166), .nRES(w112), .D(w108), .C(w853) );
	io_DFFRPOS g_185 (.Q(w120), .nRES(w112), .D(w336), .C(w853) );
	io_DFFRPOS g_186 (.Q(w51), .nRES(w112), .D(w138), .C(w853) );
	io_AND g_187 (.Z(w895), .B(w230), .A(w324) );
	io_CNT_BIT g_188 (.nQ(w889), .C(w115), .nRES(1'b1), .D(1'b1), .nLD(w119), .CO(w219), .CI(w877) );
	io_DFFRPOS g_189 (.Q(w814), .nRES(w112), .D(w186), .C(w853) );
	io_DFFRPOS g_190 (.Q(w241), .nRES(w112), .D(w130), .C(w853) );
	io_DFFRPOS g_191 (.Q(w133), .nRES(1'b1), .D(w130), .C(w33) );
	io_DFFRPOS g_192 (.Q(w822), .nRES(1'b1), .D(w138), .C(w33) );
	io_DFFRPOS g_193 (.Q(w817), .nRES(w112), .D(w130), .C(w140) );
	io_DFFRPOS g_194 (.Q(w813), .nRES(w112), .D(w186), .C(w140) );
	io_DFFRPOS g_195 (.Q(w803), .nRES(w112), .D(w138), .C(w140) );
	io_AND g_196 (.Z(w891), .B(w366), .A(w324) );
	io_DFFRPOS g_197 (.Q(w867), .nRES(1'b1), .D(w186), .C(w142) );
	io_AND g_198 (.Z(w871), .B(w32), .A(w8) );
	io_MUX4BIT g_199 (.S(w53), .Z0(w278), .A0(w893), .B0(w902), .A1(w231), .B1(w901), .Z1(w279), .Z2(w281), .B2(w928), .A2(w238), .A3(w886), .B3(w225), .Z3(w282) );
	io_DFFRPOS g_200 (.Q(w263), .nRES(w112), .D(w165), .C(w853) );
	io_MUX4BIT g_201 (.S(w871), .Z0(w902), .A0(w894), .B0(w899), .A1(w903), .B1(w897), .Z1(w901), .Z2(w928), .B2(w827), .A2(w158), .A3(w892), .B3(w670), .Z3(w225) );
	io_DFFRPOS g_202 (.Q(w896), .nRES(1'b1), .D(w900), .C(w712) );
	io_NOR6 g_203 (.Z(w56), .F(w794), .E(w239), .D(w868), .C(w907), .B(w906), .A(w870) );
	io_MUX8TO1 g_204 (.S0(w250), .S2(w247), .S1(w251), .G(w858), .H(w866), .F(w747), .E(w898), .Z(w897), .C(w869), .D(w896), .B(w904), .A(w919) );
	io_AND g_205 (.Z(w907), .B(w829), .A(w265) );
	io_AND g_206 (.Z(w870), .B(w839), .A(w269) );
	io_AND g_207 (.Z(w906), .B(w828), .A(w270) );
	io_DFFRPOS g_208 (.Q(w671), .nRES(1'b1), .D(w927), .C(w712) );
	io_SIPO_4BIT g_209 (.C(w362), .D(w751), .nRES(w178), .Q0(w922), .Q1(w924), .Q2(w842), .Q3(w865) );
	io_DFFRPOS g_210 (.Q(w925), .nRES(1'b1), .D(w864), .C(w637) );
	io_DFFRPOS g_211 (.Q(w898), .nRES(w918), .D(w926), .C(w712) );
	io_DFFSPOS g_212 (.C(w623), .D(w23), .nSET(w178), .nQ(w926), .Q(w844) );
	io_DFFRPOS g_213 (.Q(w845), .nRES(1'b1), .D(w273), .C(w436) );
	io_DFFRPOS g_214 (.Q(w863), .nRES(1'b1), .D(w862), .C(w436) );
	io_DFFRPOS g_215 (.Q(w828), .nRES(w918), .D(1'b1), .C(w712) );
	io_DFFRPOS g_216 (.Q(w262), .nRES(1'b1), .D(w861), .C(w712) );
	io_AND g_217 (.Z(w918), .B(w859), .A(w860) );
	io_NAND4 g_218 (.A(w856), .D(w737), .B(w913), .C(w446), .Z(w364) );
	io_AND g_219 (.Z(w857), .B(w737), .A(w446) );
	io_DFFRPOS g_220 (.nQ(w913), .nRES(w461), .D(w854), .C(w623) );
	io_NAND g_221 (.A(w872), .B(w912), .Z(w854) );
	io_OR g_222 (.A(w913), .Z(w912), .B(w700) );
	io_OR g_223 (.A(w699), .Z(w872), .B(w700) );
	io_NOR3 g_224 (.Z(w700), .C(w913), .B(w844), .A(w911) );
	io_NOT g_225 (.A(w857), .nZ(w911) );
	io_NOT g_226 (.A(w844), .nZ(w856) );
	io_NOT g_227 (.A(w855), .nZ(w849) );
	io_NOT g_228 (.A(w589), .nZ(w728) );
	io_DFFRPOS g_229 (.Q(w777), .nRES(w50), .D(w778), .C(w727) );
	io_AON22 g_230 (.Z(w778), .B2(w731), .A2(w728), .B1(w779), .A1(w768) );
	io_DFFRPOS g_231 (.Q(w779), .nRES(w50), .D(w776), .C(w727) );
	io_AON22 g_232 (.Z(w875), .B2(w731), .A2(w770), .B1(w777), .A1(w728) );
	io_AON22 g_233 (.Z(w776), .B2(w731), .A2(w728), .B1(w775), .A1(w772) );
	io_DFFRPOS g_234 (.Q(w775), .nRES(w50), .D(w774), .C(w727) );
	io_AON22 g_235 (.Z(w774), .B2(w773), .A2(w728), .B1(w731), .A1(w757) );
	io_DFFRPOS g_236 (.Q(w773), .nRES(w50), .D(w755), .C(w727) );
	io_BUF g_237 (.Z(w609), .A(w127) );
	io_TFF g_238 (.Q(w615), .T(w609), .C(w769) );
	io_TFF g_239 (.Q(w759), .T(w609), .C(w758) );
	io_TFF g_240 (.Q(w722), .T(w609), .C(w759) );
	io_DFFSPOS g_241 (.C(w412), .D(w614), .nSET(w261), .Q(w761) );
	io_AND3 g_242 (.Z(w877), .C(1'b1), .B(w119), .A(w390) );
	io_TFF g_243 (.Q(w769), .T(w609), .C(w762) );
	io_TFF g_244 (.Q(w762), .T(w609), .C(w722) );
	io_MUX g_245 (.C(w324), .Z(w767), .A(w121), .B(w876) );
	io_SLATCH g_246 (.nQ(w768), .C(w673), .Q(w878), .D(w156) );
	io_AND g_247 (.Z(w763), .B(w261), .A(w761) );
	io_MUX g_248 (.C(w324), .Z(w758), .A(w876), .B(w115) );
	io_SLATCH g_249 (.nQ(w874), .C(w673), .Q(w672), .D(w143) );
	io_SLATCH g_250 (.nQ(w770), .C(w673), .Q(w869), .D(w108) );
	io_SLATCH g_251 (.nQ(w771), .C(w673), .Q(w764), .D(w130) );
	io_SLATCH g_252 (.nQ(w772), .C(w673), .Q(w821), .D(w186) );
	io_MUX4BIT g_253 (.S(w871), .Z0(w753), .A0(w807), .B0(w809), .A1(w766), .B1(w818), .Z1(w756), .Z2(w819), .B2(w820), .A2(w806), .A3(w812), .B3(w805), .Z3(w725) );
	io_OR g_254 (.A(w96), .Z(w804), .B(w153) );
	io_AND g_255 (.Z(w802), .B(w189), .A(w804) );
	io_MUX4BIT g_256 (.S(w8), .Z0(w934), .A0(w802), .B0(w822), .A1(w801), .B1(w189), .Z1(w800), .Z2(w795), .B2(w23), .A2(1'b0), .A3(1'b1), .B3(w242), .Z3(w793) );
	io_MUX8TO1 g_257 (.S0(w797), .S2(w183), .S1(w128), .G(w678), .H(w734), .F(w263), .E(w275), .Z(w806), .C(w795), .D(w318), .B(w243), .A(w346) );
	io_OR g_258 (.B(w69), .Z(w785), .A(w153) );
	io_AND g_259 (.Z(w801), .B(w70), .A(w785) );
	io_NOT g_260 (.A(w813), .nZ(w783) );
	io_DFFRPOS g_261 (.Q(w790), .nRES(w112), .D(w186), .C(w430) );
	io_BUF g_262 (.Z(w859), .A(w127) );
	io_NOT g_263 (.A(w803), .nZ(w786) );
	io_NOR g_264 (.Z(w868), .B(w786), .A(w70) );
	io_AND g_265 (.Z(w155), .B(w783), .A(w784) );
	io_AND g_266 (.Z(w788), .B(w324), .A(w623) );
	io_NOT g_267 (.A(w261), .nZ(w784) );
	io_AND g_268 (.Z(w782), .B(w867), .A(w784) );
	io_AND g_269 (.Z(w256), .B(w324), .A(w412) );
	io_OR g_270 (.B(w782), .Z(w74), .A(w763) );
	io_MUX8TO1 g_271 (.S0(w797), .S2(w183), .S1(w128), .G(w653), .H(w816), .F(w746), .E(w721), .Z(w818), .C(w764), .D(w835), .B(w815), .A(w838) );
	io_DFFRPOS g_272 (.Q(w866), .nRES(w836), .D(w677), .C(w637) );
	io_DFFRPOS g_273 (.Q(w815), .nRES(w112), .D(w130), .C(w137) );
	io_DFFRPOS g_274 (.Q(w835), .nRES(1'b1), .D(w837), .C(w712) );
	io_SIPO_4BIT g_275 (.C(w379), .D(w655), .nRES(w271), .Q0(w873), .Q1(w834), .Q2(w840), .Q3(w667) );
	io_MUX8TO1 g_276 (.S0(w797), .S2(w183), .S1(w128), .G(w702), .H(w271), .F(w557), .E(w178), .Z(w820), .C(w833), .D(w716), .B(w276), .A(w863) );
	io_DFFRPOS g_277 (.Q(w721), .nRES(w112), .D(w130), .C(w176) );
	io_DFFRPOS g_278 (.Q(w858), .nRES(1'b1), .D(w847), .C(w637) );
	io_AND g_279 (.Z(w836), .B(w167), .A(w859) );
	io_DFFRPOS g_280 (.Q(w829), .nRES(w836), .D(1'b1), .C(w637) );
	io_DFFRPOS g_281 (.Q(w825), .nRES(1'b1), .D(w851), .C(w436) );
	io_NOR3 g_282 (.Z(w739), .C(w849), .B(w172), .A(w16) );
	io_NAND4 g_283 (.A(w739), .D(w738), .B(w741), .C(w740), .Z(w333) );
	io_NAND4 g_284 (.A(w740), .D(w742), .B(w739), .C(w743), .Z(w853) );
	io_NAND4 g_285 (.A(w739), .D(w744), .B(w741), .C(w738), .Z(w33) );
	io_NAND4 g_286 (.B(w741), .C(w740), .A(w739), .D(w743), .Z(w142) );
	io_NAND4 g_287 (.B(w742), .C(w744), .A(w739), .D(w743), .Z(w140) );
	io_NOT g_288 (.A(w240), .nZ(w752) );
	io_MUX4BIT g_289 (.S(w53), .Z0(w205), .A0(w289), .B0(w753), .A1(w288), .B1(w756), .Z1(w203), .Z2(w201), .B2(w819), .A2(w286), .A3(w283), .B3(w725), .Z3(w200) );
	io_MUX4BIT g_290 (.S(w227), .Z0(w726), .A0(w206), .B0(w217), .A1(w204), .B1(w216), .Z1(w754), .Z2(w723), .B2(w215), .A2(w202), .A3(w199), .B3(w214), .Z3(w724) );
	io_AON22 g_291 (.Z(w755), .B2(w731), .A2(w728), .B1(w730), .A1(w771) );
	io_MUX4BIT g_292 (.S(w752), .Z0(w138), .A0(w206), .B0(w289), .A1(w204), .B1(w288), .Z1(w130), .Z2(w165), .B2(w286), .A2(w202), .A3(w199), .B3(w283), .Z3(w186) );
	io_MUX4BIT g_293 (.S(w53), .Z0(w290), .A0(w726), .B0(w753), .A1(w754), .B1(w756), .Z1(w287), .Z2(w285), .B2(w819), .A2(w723), .A3(w724), .B3(w725), .Z3(w284) );
	io_MUX2BIT4TO1 g_294 (.A0(w769), .A1(w611), .ZA(w412), .A3(w720), .A2(w615), .B0(w758), .B1(w722), .ZB(w366), .B3(w769), .B2(w759), .S1(w815), .S0(w787) );
	io_MUX2BIT4TO1 g_295 (.A0(w769), .A1(w611), .ZA(w230), .A3(w720), .A2(w615), .B0(w758), .B1(w722), .ZB(w623), .B3(w769), .B2(w759), .S1(w721), .S0(w808) );
	io_MUX2BIT4TO1 g_296 (.A0(w769), .A1(w611), .ZA(w345), .A3(w720), .A2(w615), .B0(w758), .B1(w722), .ZB(w426), .B3(w769), .B2(w759), .S1(w816), .S0(w791) );
	io_SLATCH g_297 (.nQ(w719), .C(w673), .Q(w789), .D(w138) );
	io_MUX8TO1 g_298 (.S0(w797), .S2(w183), .S1(w128), .G(w352), .H(w729), .F(w241), .E(w817), .Z(w766), .C(w800), .D(w321), .B(w760), .A(w767) );
	io_MUX8TO1 g_299 (.S0(w797), .S2(w183), .S1(w128), .G(w790), .H(w718), .F(w814), .E(w813), .Z(w812), .C(w793), .D(w317), .B(w244), .A(w604) );
	io_NOT g_300 (.A(w733), .nZ(w792) );
	io_NOR g_301 (.Z(w794), .B(w321), .A(w792) );
	io_DFFRPOS g_302 (.Q(w733), .nRES(w112), .D(w138), .C(w430) );
	io_MUX8TO1 g_303 (.S0(w797), .S2(w183), .S1(w128), .G(w733), .H(w732), .F(w51), .E(w803), .Z(w807), .C(w934), .D(w368), .B(w796), .A(w153) );
	io_SLATCH g_304 (.nQ(w765), .C(w673), .Q(w811), .D(w336) );
	io_NOT g_305 (.A(w790), .nZ(w810) );
	io_AND g_306 (.Z(w316), .B(w781), .A(w810) );
	io_NOT g_307 (.A(w184), .nZ(w781) );
	io_AND g_308 (.Z(w780), .B(w781), .A(w350) );
	io_MUX8TO1 g_309 (.S0(w797), .S2(w183), .S1(w128), .G(w462), .H(w791), .F(w564), .E(w808), .Z(w809), .C(w789), .D(w713), .B(w787), .A(w823) );
	io_AND g_310 (.Z(w824), .B(w184), .A(w735) );
	io_OR g_311 (.B(w780), .Z(w315), .A(w824) );
	io_DFFRPOS g_312 (.Q(w791), .nRES(w112), .D(w138), .C(w86) );
	io_MUX8TO1 g_313 (.S0(w250), .S2(w247), .S1(w251), .G(w830), .H(w829), .F(w717), .E(w828), .Z(w827), .C(w811), .D(w826), .B(w839), .A(w825) );
	io_DFFRPOS g_314 (.Q(w816), .nRES(w112), .D(w130), .C(w86) );
	io_DFFRPOS g_315 (.Q(w826), .nRES(1'b1), .D(w841), .C(w712) );
	io_DFFRPOS g_316 (.Q(w830), .nRES(1'b1), .D(w846), .C(w637) );
	io_MUX8TO1 g_317 (.S0(w797), .S2(w183), .S1(w128), .G(w832), .H(w184), .F(w680), .E(w50), .Z(w805), .C(w821), .D(w831), .B(w261), .A(w845) );
	io_DFFRPOS g_318 (.Q(w831), .nRES(1'b1), .D(w750), .C(w712) );
	io_SLATCH g_319 (.nQ(w757), .C(w673), .Q(w833), .D(w165) );
	io_DFFRPOS g_320 (.Q(w832), .nRES(1'b1), .D(w843), .C(w637) );
	io_DFFRPOS g_321 (.Q(w808), .nRES(w112), .D(w138), .C(w176) );
	io_BUF g_322 (.Z(w250), .A(w848) );
	io_BUF g_323 (.Z(w797), .A(w848) );
	io_XNOR g_324 (.A(w9), .B(w8), .Z(w848) );
	io_NOT g_325 (.A(w2), .nZ(w711) );
	io_NOT g_326 (.A(w17), .nZ(w710) );
	io_NOT g_327 (.A(w17), .nZ(w741) );
	io_NOT g_328 (.A(w9), .nZ(w744) );
	io_NAND4 g_329 (.B(w744), .C(w738), .A(w742), .D(w739), .Z(w430) );
	io_NOT g_330 (.A(w2), .nZ(w743) );
	io_NAND4 g_331 (.B(w739), .C(w740), .A(w738), .D(w742), .Z(w569) );
	io_NOT g_332 (.A(w743), .nZ(w738) );
	io_NAND4 g_333 (.B(w744), .C(w739), .A(w743), .D(w741) );
	io_NOT g_334 (.A(w741), .nZ(w742) );
	io_NOR3 g_335 (.Z(w708), .C(w16), .B(w172), .A(w745) );
	io_NOT g_336 (.A(w744), .nZ(w740) );
	io_NOT g_337 (.A(w32), .nZ(w745) );
	io_AND g_338 (.Z(w208), .B(w240), .A(w192) );
	io_MUX g_339 (.C(w240), .Z(w207), .A(w608), .B(w193) );
	io_DFFRPOS g_340 (.Q(w608), .nRES(w127), .D(w199), .C(w607) );
	io_OR g_341 (.B(w9), .Z(w607), .A(w6) );
	io_OR g_342 (.A(w230), .Z(w727), .B(1'b0) );
	io_AON22 g_343 (.Z(w605), .B2(w731), .A2(w719), .B1(1'b0), .A1(w728) );
	io_DFFRPOS g_344 (.Q(w730), .nRES(w50), .D(w605), .C(w727) );
	io_TFF g_345 (.Q(w720), .T(w609), .C(w610) );
	io_TFF g_346 (.Q(w610), .T(w609), .C(w611) );
	io_TFF g_347 (.Q(w611), .T(w609), .C(w615) );
	io_NOT g_348 (.A(w589), .nZ(w613) );
	io_NOT g_349 (.A(w230), .nZ(w612) );
	io_NOT g_350 (.A(w663), .nZ(w619) );
	io_AND g_351 (.Z(w614), .B(w506), .A(w617) );
	io_NOT g_352 (.A(w618), .nZ(w617) );
	io_DFFRPOS g_353 (.Q(w618), .nRES(w261), .D(w620), .C(w601) );
	io_JKFFSRNEG g_354 (.C(w612), .K(1'b0), .J(w613), .nSET(w628), .nRES(w533), .Q(w625), .nQ(w621) );
	io_DFFRPOS g_355 (.Q(w627), .nRES(w261), .D(w626), .C(w601) );
	io_AON22 g_356 (.Z(w620), .B2(w624), .A2(w629), .B1(w627), .A1(w597) );
	io_AON22 g_357 (.Z(w626), .B2(w624), .A2(w597), .B1(w630), .A1(w631) );
	io_DFFRPOS g_358 (.Q(w630), .nRES(w261), .D(w640), .C(w601) );
	io_AON22 g_359 (.Z(w641), .B2(w624), .A2(w642), .B1(w633), .A1(w597) );
	io_DFFRPOS g_360 (.Q(w639), .nRES(w261), .D(w641), .C(w601) );
	io_AON22 g_361 (.Z(w640), .B1(w624), .A2(w597), .B2(w639), .A1(w638) );
	io_SLATCH g_362 (.nQ(w634), .C(w643), .Q(w718), .D(w186) );
	io_NOT g_363 (.A(w569), .nZ(w643) );
	io_SLATCH g_364 (.nQ(w645), .C(w643), .Q(w729), .D(w130) );
	io_SLATCH g_365 (.nQ(w644), .C(w643), .Q(w734), .D(w165) );
	io_SLATCH g_366 (.nQ(w638), .C(w643), .Q(w650), .D(w108) );
	io_SLATCH g_367 (.nQ(w642), .C(w643), .Q(w248), .D(w156) );
	io_SLATCH g_368 (.nQ(w629), .C(w643), .Q(w253), .D(w143) );
	io_SLATCH g_369 (.nQ(w631), .C(w643), .Q(w159), .D(w336) );
	io_SLATCH g_370 (.nQ(w649), .C(w643), .Q(w732), .D(w138) );
	io_DFFSPOS g_371 (.C(w345), .D(w651), .nSET(w184), .Q(w735) );
	io_AND g_372 (.Z(w651), .B(w387), .A(w685) );
	io_SLATCH g_373 (.nQ(w568), .C(w567), .Q(w746), .D(w130) );
	io_NOT g_374 (.A(w682), .nZ(w685) );
	io_SLATCH g_375 (.nQ(w679), .C(w567), .Q(w747), .D(w108) );
	io_BUF g_376 (.Z(w431), .A(w127) );
	io_DFFRPOS g_377 (.Q(w682), .nRES(w184), .D(w681), .C(w538) );
	io_SLATCH g_378 (.nQ(w933), .C(w567), .Q(w680), .D(w186) );
	io_DFFRPOS g_379 (.Q(w678), .nRES(w112), .D(w165), .C(w430) );
	io_NOT g_380 (.A(w678), .nZ(w674) );
	io_DFFSPOS g_381 (.C(w426), .D(w318), .nSET(w271), .nQ(w677), .Q(w663) );
	io_OR g_382 (.A(w674), .Z(w319), .B(w271) );
	io_SLATCH g_383 (.nQ(w688), .C(w567), .Q(w717), .D(w336) );
	io_SLATCH g_384 (.nQ(w560), .C(w567), .Q(w676), .D(w156) );
	io_SLATCH g_385 (.nQ(w675), .C(w567), .Q(w668), .D(w143) );
	io_NOT g_386 (.A(w666), .nZ(w567) );
	io_MUX8TO1 g_387 (.S0(w250), .S2(w247), .S1(w251), .G(w660), .H(w665), .F(w668), .E(w625), .Z(w670), .C(w672), .D(w671), .B(w566), .A(w669) );
	io_NOT g_388 (.A(w628), .nZ(w673) );
	io_DFFRPOS g_389 (.Q(w669), .nRES(1'b1), .D(w736), .C(w436) );
	io_DFFRPOS g_390 (.Q(w713), .nRES(1'b1), .D(w689), .C(w712) );
	io_DFFRPOS g_391 (.Q(w716), .nRES(1'b1), .D(w691), .C(w712) );
	io_SIPO_4BIT g_392 (.C(w362), .D(w693), .nRES(w178), .Q0(w692), .Q1(w749), .Q2(w690), .Q3(w751) );
	io_BUF g_393 (.Z(w435), .A(w431) );
	io_AND g_394 (.Z(w693), .B(w844), .A(1'b1) );
	io_BUF g_395 (.Z(w461), .A(w431) );
	io_NAND4 g_396 (.B(w711), .C(w707), .A(w708), .D(w709), .Z(w666) );
	io_NAND4 g_397 (.B(w709), .C(w705), .A(w708), .D(w707), .Z(w86) );
	io_NOT g_398 (.A(w711), .nZ(w705) );
	io_NAND4 g_399 (.B(w708), .C(w709), .A(w710), .D(w705) );
	io_NAND4 g_400 (.B(w711), .C(w708), .A(w710), .D(w709), .Z(w137) );
	io_NOT g_401 (.A(w706), .nZ(w709) );
	io_NAND4 g_402 (.B(w711), .C(w706), .A(w710), .D(w708) );
	io_NAND4 g_403 (.B(w711), .C(w706), .A(w708), .D(w707), .Z(w176) );
	io_NAND4 g_404 (.B(w710), .C(w705), .A(w708), .D(w706), .Z(w628) );
	io_NAND4 g_405 (.B(w705), .C(w706), .A(w708), .D(w707) );
	io_NOT g_406 (.A(w710), .nZ(w707) );
	io_NOT g_407 (.A(w9), .nZ(w706) );
	io_DFFSPOS g_408 (.C(w362), .D(w363), .nSET(w435), .Q(w704) );
	io_OR g_409 (.B(w362), .Z(w712), .A(w704) );
	io_DFFSPOS g_410 (.C(w623), .D(w698), .nSET(w461), .nQ(w362), .Q(w699) );
	io_DFFRPOS g_411 (.nQ(w580), .Q(w574), .nRES(w588), .D(w584), .C(w230) );
	io_NAND6 g_412 (.C(w587), .D(w582), .B(w586), .E(w581), .A(1'b1), .F(w580), .Z(w589) );
	io_NAND3 g_413 (.A(w582), .B(w581), .C(w580), .Z(w572) );
	io_DFFRPOS g_414 (.nQ(w586), .Q(w571), .nRES(w588), .D(w577), .C(w230) );
	io_NAND4 g_415 (.B(w574), .C(w581), .A(w586), .D(w583), .Z(w570) );
	io_DFFRPOS g_416 (.nQ(w587), .Q(w583), .nRES(w588), .D(w578), .C(w230) );
	io_NAND4 g_417 (.B(w586), .C(w574), .A(w587), .D(w581), .Z(w590) );
	io_DFFRPOS g_418 (.nQ(w581), .Q(w575), .nRES(w588), .D(w579), .C(w230) );
	io_DFFSPOS g_419 (.C(w230), .D(w590), .nSET(w588), .Q(w595) );
	io_BUF g_420 (.Z(w588), .A(w431) );
	io_NOT g_421 (.A(w594), .nZ(w593) );
	io_NOR3 g_422 (.Z(w591), .C(w593), .B(w663), .A(w596) );
	io_OR g_423 (.A(w591), .Z(w599), .B(w596) );
	io_NAND g_424 (.A(w599), .B(w592), .Z(w598) );
	io_DFFRPOS g_425 (.nQ(w596), .nRES(w500), .D(w598), .C(w426) );
	io_DFFSRPOS g_426 (.C(w595), .D(1'b0), .nRES(w533), .nSET(w621), .Q(w622) );
	io_AND g_427 (.Z(w594), .B(w388), .A(w377) );
	io_NAND4 g_428 (.B(w596), .C(w377), .A(w619), .D(w388), .Z(w378) );
	io_DFFPOS g_429 (.Q(w582), .D(w622), .C(w623) );
	io_NOT g_430 (.A(w597), .nZ(w624) );
	io_BUF g_431 (.Z(w374), .A(w431) );
	io_BUF g_432 (.Z(w533), .A(w127) );
	io_OR g_433 (.B(1'b0), .Z(w601), .A(w412) );
	io_DFFRPOS g_434 (.Q(w633), .nRES(w261), .D(w632), .C(w601) );
	io_AON22 g_435 (.Z(w632), .B2(w624), .A2(w597), .B1(w635), .A1(w634) );
	io_DFFSPOS g_436 (.C(w379), .D(w299), .nSET(w374), .Q(w636) );
	io_OR g_437 (.A(w379), .Z(w637), .B(w636) );
	io_DFFRPOS g_438 (.Q(w635), .nRES(w261), .D(w684), .C(w601) );
	io_AON22 g_439 (.Z(w684), .B2(w624), .A2(w644), .B1(w646), .A1(w597) );
	io_AON22 g_440 (.Z(w647), .B2(w624), .A2(w649), .B1(1'b0), .A1(w597) );
	io_AON22 g_441 (.Z(w602), .B2(w624), .A2(w645), .B1(w648), .A1(w597) );
	io_DFFRPOS g_442 (.Q(w648), .nRES(w261), .D(w647), .C(w601) );
	io_DFFRPOS g_443 (.Q(w646), .nRES(w261), .D(w602), .C(w601) );
	io_NOT g_444 (.A(w387), .nZ(w548) );
	io_NOT g_445 (.A(w387), .nZ(w563) );
	io_DFFRPOS g_446 (.Q(w603), .nRES(w184), .D(w600), .C(w538) );
	io_AON22 g_447 (.Z(w600), .B2(w547), .A2(w679), .B1(w683), .A1(w548) );
	io_DFFRPOS g_448 (.Q(w683), .nRES(w184), .D(w565), .C(w538) );
	io_AON22 g_449 (.Z(w565), .B2(w547), .A2(w548), .B1(w558), .A1(w560) );
	io_AON22 g_450 (.Z(w561), .B2(w547), .A2(w933), .B1(w549), .A1(w548) );
	io_DFFRPOS g_451 (.Q(w558), .nRES(w184), .D(w561), .C(w538) );
	io_DFFRPOS g_452 (.Q(w559), .nRES(w184), .D(w687), .C(w538) );
	io_AON22 g_453 (.Z(w687), .B2(w547), .A2(w688), .B1(w603), .A1(w548) );
	io_AON22 g_454 (.Z(w681), .B2(w547), .A2(w548), .B1(w559), .A1(w675) );
	io_NOT g_455 (.A(w345), .nZ(w686) );
	io_JKFFSRNEG g_456 (.C(w686), .K(1'b0), .J(w563), .nSET(w666), .nRES(w533), .Q(w665), .nQ(w664) );
	io_DFFSRPOS g_457 (.C(w513), .D(1'b0), .nRES(w533), .nSET(w664), .Q(w555) );
	io_AND g_458 (.Z(w658), .B(1'b1), .A(w663) );
	io_DFFRPOS g_459 (.Q(w660), .nRES(1'b1), .D(w659), .C(w637) );
	io_SIPO_4BIT g_460 (.C(w379), .D(w658), .nRES(w271), .Q0(w656), .Q1(w657), .Q2(w661), .Q3(w655) );
	io_DFFRPOS g_461 (.Q(w653), .nRES(1'b1), .D(w654), .C(w637) );
	io_DFFRPOS g_462 (.Q(w462), .nRES(1'b1), .D(w652), .C(w637) );
	io_DFFSPOS g_463 (.C(w623), .D(w451), .nSET(w461), .nQ(w456), .Q(w453) );
	io_DFFSPOS g_464 (.C(w623), .D(w459), .nSET(w461), .nQ(w445), .Q(w457) );
	io_NAND4 g_465 (.B(w445), .C(w456), .A(w362), .D(w455), .Z(w463) );
	io_DFFRPOS g_466 (.nQ(w737), .Q(w433), .nRES(w435), .D(w443), .C(w362) );
	io_DFFRPOS g_467 (.Q(w702), .nRES(1'b1), .D(w703), .C(w637) );
	io_DFFRPOS g_468 (.nQ(w454), .Q(w455), .nRES(w461), .D(w701), .C(w623) );
	io_NOR g_469 (.Z(w701), .B(w455), .A(w700) );
	io_NOT g_470 (.A(w700), .nZ(w452) );
	io_NAND6 g_471 (.C(w696), .D(w465), .B(w695), .E(w463), .A(1'b1), .F(w452), .Z(w698) );
	io_NAND g_472 (.A(w699), .B(w457), .Z(w465) );
	io_NAND g_473 (.A(w699), .B(w453), .Z(w696) );
	io_NAND g_474 (.A(w454), .B(w699), .Z(w695) );
	io_NAND3 g_475 (.A(w485), .B(w570), .C(w572), .Z(w577) );
	io_NAND4 g_476 (.B(w576), .C(w486), .A(w570), .D(w485), .Z(w584) );
	io_NAND g_477 (.A(w575), .B(w574), .Z(w486) );
	io_NAND g_478 (.A(w571), .B(w574), .Z(w576) );
	io_NAND g_479 (.A(w575), .B(w571), .Z(w485) );
	io_NAND3 g_480 (.A(w575), .B(w571), .C(w580), .Z(w488) );
	io_NAND g_481 (.A(w581), .B(w574), .Z(w487) );
	io_NAND3 g_482 (.A(w487), .B(w572), .C(w488), .Z(w579) );
	io_NAND4 g_483 (.B(w572), .C(w488), .A(w573), .D(w489), .Z(w578) );
	io_NAND3 g_484 (.A(w583), .B(w575), .C(w574), .Z(w489) );
	io_NAND3 g_485 (.A(w574), .B(w583), .C(w571), .Z(w573) );
	io_NAND4 g_486 (.B(w492), .C(w491), .A(w379), .D(w501), .Z(w519) );
	io_NOT g_487 (.A(w591), .nZ(w498) );
	io_NOR g_488 (.Z(w508), .B(w501), .A(w591) );
	io_DFFRPOS g_489 (.nQ(w507), .Q(w501), .nRES(w500), .D(w508), .C(w426) );
	io_BUF g_490 (.Z(w500), .A(w431) );
	io_BUF g_491 (.Z(w410), .A(w431) );
	io_DFFSPOS g_492 (.C(w426), .D(w509), .nSET(w500), .nQ(w379), .Q(w514) );
	io_NAND g_493 (.A(w507), .B(w514), .Z(w515) );
	io_NAND6 g_494 (.C(1'b1), .D(w516), .B(w520), .E(w515), .A(w519), .F(w498), .Z(w509) );
	io_NAND g_495 (.A(w514), .B(w495), .Z(w520) );
	io_NAND g_496 (.A(w514), .B(w490), .Z(w516) );
	io_OR g_497 (.A(w514), .Z(w592), .B(w591) );
	io_DFFSPOS g_498 (.C(w412), .D(w505), .nSET(w410), .Q(w511) );
	io_NOT g_499 (.A(w506), .nZ(w597) );
	io_NOT g_500 (.A(w506), .nZ(w512) );
	io_BUF g_501 (.Z(w401), .A(w431) );
	io_DFFSPOS g_502 (.C(w345), .D(w510), .nSET(w401), .Q(w513) );
	io_NAND4 g_503 (.B(w386), .C(w383), .A(w393), .D(w382), .Z(w510) );
	io_DFFSRPOS g_504 (.C(w511), .D(1'b0), .nRES(w533), .nSET(w526), .Q(w517) );
	io_JKFFSRNEG g_505 (.c(w534), .K(1'b0), .J(w512), .nSET(w569), .nRES(w533), .Q(w566), .nQ(w526) );
	io_NOT g_506 (.A(w412), .nZ(w534) );
	io_DFFPOS g_507 (.Q(w527), .D(w555), .C(w426) );
	io_AND g_508 (.Z(w604), .B(w426), .A(w324) );
	io_DFFRPOS g_509 (.Q(w528), .nRES(w184), .D(w529), .C(w538) );
	io_BUF g_510 (.Z(w365), .A(w431) );
	io_AON22 g_511 (.Z(w529), .B2(w536), .A2(w568), .B1(w547), .A1(w548) );
	io_NOT g_512 (.A(w548), .nZ(w547) );
	io_DFFRPOS g_513 (.Q(w536), .nRES(w184), .D(w539), .C(w538) );
	io_AON22 g_514 (.Z(w539), .B2(w547), .A2(w548), .B1(1'b0), .A1(w540) );
	io_OR g_515 (.B(w345), .Z(w538), .A(1'b0) );
	io_AON22 g_516 (.Z(w546), .B2(w547), .A2(w482), .B1(w528), .A1(w548) );
	io_DFFRPOS g_517 (.Q(w549), .nRES(w184), .D(w546), .C(w538) );
	io_SLATCH g_518 (.nQ(w540), .C(w567), .Q(w564), .D(w138) );
	io_SLATCH g_519 (.nQ(w482), .C(w567), .Q(w557), .D(w165) );
	io_NOT g_520 (.A(w474), .nZ(w481) );
	io_NOR3 g_521 (.Z(w373), .C(w478), .B(w556), .A(w481) );
	io_DFFRPOS g_522 (.nQ(w478), .nRES(w365), .D(w479), .C(w366) );
	io_OR g_523 (.B(w480), .Z(w483), .A(w373) );
	io_NAND g_524 (.A(w484), .B(w483), .Z(w479) );
	io_OR g_525 (.B(w478), .Z(w484), .A(w373) );
	io_DFFRPOS g_526 (.Q(w477), .nRES(w112), .D(w108), .C(w430) );
	io_NOT g_527 (.A(w477), .nZ(w331) );
	io_DFFRPOS g_528 (.Q(w255), .nRES(w112), .D(w156), .C(w430) );
	io_NOT g_529 (.A(w556), .nZ(w554) );
	io_AND g_530 (.Z(w474), .B(w354), .A(w466) );
	io_NAND4 g_531 (.B(w478), .C(w466), .A(w554), .D(w354), .Z(w476) );
	io_NOT g_532 (.A(w255), .nZ(w313) );
	io_NAND4 g_533 (.B(w553), .C(w473), .A(w476), .D(w472), .Z(w432) );
	io_NAND g_534 (.A(w469), .B(w353), .Z(w473) );
	io_DFFRPOS g_535 (.nQ(w466), .Q(w469), .nRES(w357), .D(w475), .C(w355) );
	io_NAND4 g_536 (.B(w553), .C(w472), .A(w476), .D(w356), .Z(w475) );
	io_NAND3 g_537 (.A(w470), .B(w466), .C(w353), .Z(w472) );
	io_DFFRPOS g_538 (.nQ(w551), .Q(w470), .nRES(w357), .D(w429), .C(w355) );
	io_NAND4 g_539 (.B(w553), .C(w471), .A(w476), .D(w356), .Z(w429) );
	io_NAND3 g_540 (.A(w469), .B(w470), .C(w353), .Z(w471) );
	io_NAND4 g_541 (.B(w551), .C(w466), .A(w550), .D(w353), .Z(w553) );
	io_NAND4 g_542 (.B(w551), .C(w466), .A(w552), .D(w353), .Z(w356) );
	io_DFFRPOS g_543 (.nQ(w552), .Q(w550), .nRES(w357), .D(w467), .C(w355) );
	io_NAND4 g_544 (.B(w460), .C(w468), .A(w476), .D(w356), .Z(w467) );
	io_NAND3 g_545 (.A(w353), .B(w550), .C(w470), .Z(w468) );
	io_NAND3 g_546 (.A(w469), .B(w550), .C(w353), .Z(w460) );
	io_NAND4 g_547 (.A(w458), .D(w450), .B(w452), .C(w448), .Z(w459) );
	io_NAND g_548 (.A(w453), .B(w457), .Z(w458) );
	io_NAND g_549 (.A(w454), .B(w457), .Z(w450) );
	io_NAND3 g_550 (.A(w455), .B(w456), .C(w445), .Z(w448) );
	io_NAND g_551 (.A(w455), .B(w456), .Z(w449) );
	io_NAND g_552 (.A(w454), .B(w453), .Z(w447) );
	io_NAND3 g_553 (.A(w449), .B(w447), .C(w452), .Z(w451) );
	io_NAND4 g_554 (.B(w446), .C(w359), .A(w433), .D(w440), .Z(w363) );
	io_NAND4 g_555 (.B(w446), .C(w360), .A(w433), .D(w440), .Z(w442) );
	io_NAND3 g_556 (.A(w433), .B(w434), .C(w446), .Z(w438) );
	io_DFFRPOS g_557 (.nQ(w446), .Q(w428), .nRES(w435), .D(w444), .C(w362) );
	io_NAND4 g_558 (.B(w442), .C(w438), .A(w363), .D(w364), .Z(w444) );
	io_DFFRPOS g_559 (.nQ(w440), .Q(w434), .nRES(w435), .D(w441), .C(w362) );
	io_NAND4 g_560 (.B(w442), .C(w439), .A(w363), .D(w364), .Z(w441) );
	io_NAND4 g_561 (.B(w364), .C(w437), .A(w442), .D(w438), .Z(w443) );
	io_NAND3 g_562 (.A(w433), .B(w428), .C(w434), .Z(w439) );
	io_NAND g_563 (.A(w428), .B(w433), .Z(w437) );
	io_NAND g_564 (.A(w507), .B(w495), .Z(w493) );
	io_NAND g_565 (.A(w507), .B(w490), .Z(w494) );
	io_NAND g_566 (.A(w490), .B(w495), .Z(w421) );
	io_NAND4 g_567 (.B(w493), .C(w421), .A(w498), .D(w422), .Z(w499) );
	io_NAND3 g_568 (.A(w494), .B(w498), .C(w497), .Z(w496) );
	io_NAND g_569 (.A(w501), .B(w491), .Z(w497) );
	io_NAND3 g_570 (.A(w492), .B(w501), .C(w491), .Z(w422) );
	io_DFFSPOS g_571 (.C(w426), .D(w496), .nSET(w500), .nQ(w491), .Q(w490) );
	io_DFFSPOS g_572 (.C(w426), .D(w499), .nSET(w500), .nQ(w492), .Q(w495) );
	io_NAND3 g_573 (.A(w503), .B(w418), .C(w415), .Z(w420) );
	io_NAND4 g_574 (.A(w502), .D(w409), .B(w296), .C(w418), .Z(w505) );
	io_NAND6 g_575 (.C(w503), .D(w409), .B(w502), .E(w415), .A(1'b1), .F(w418), .Z(w506) );
	io_DFFRPOS g_576 (.nQ(w502), .Q(w329), .nRES(w410), .D(w425), .C(w412) );
	io_DFFPOS g_577 (.Q(w503), .D(w517), .C(w366) );
	io_NAND g_578 (.A(w404), .B(w393), .Z(w408) );
	io_NAND g_579 (.A(w397), .B(w393), .Z(w518) );
	io_NAND4 g_580 (.A(w408), .D(w403), .B(w518), .C(w402), .Z(w407) );
	io_DFFRPOS g_581 (.nQ(w384), .Q(w393), .nRES(w401), .D(w407), .C(w345) );
	io_NAND4 g_582 (.B(w405), .C(w383), .A(w393), .D(w382), .Z(w403) );
	io_NAND3 g_583 (.A(w397), .B(w404), .C(w384), .Z(w398) );
	io_NAND3 g_584 (.A(w393), .B(w405), .C(w397), .Z(w406) );
	io_NAND3 g_585 (.A(w404), .B(w405), .C(w522), .Z(w524) );
	io_NAND4 g_586 (.B(w406), .C(w395), .A(w524), .D(w398), .Z(w522) );
	io_DFFRPOS g_587 (.nQ(w386), .Q(w405), .nRES(w401), .D(w522), .C(w345) );
	io_NAND3 g_588 (.A(w383), .B(w384), .C(w527), .Z(w395) );
	io_NAND6 g_589 (.C(w386), .D(w382), .B(1'b1), .E(w383), .A(w527), .F(w384), .Z(w387) );
	io_DFFRPOS g_590 (.nQ(w388), .Q(w371), .nRES(w374), .D(w531), .C(w379) );
	io_NAND g_591 (.A(w372), .B(w371), .Z(w532) );
	io_NAND4 g_592 (.B(w532), .C(w375), .A(w378), .D(w376), .Z(w531) );
	io_NAND4 g_593 (.B(w378), .C(w375), .A(w299), .D(w376), .Z(w530) );
	io_DFFRPOS g_594 (.nQ(w377), .Q(w372), .nRES(w374), .D(w530), .C(w379) );
	io_DFFPOS g_595 (.nQ(w300), .Q(w127), .D(w292), .C(w115) );
	io_NOT g_596 (.A(w373), .nZ(w338) );
	io_NOR g_597 (.Z(w541), .B(w341), .A(w373) );
	io_DFFRPOS g_598 (.nQ(w344), .Q(w341), .nRES(w365), .D(w541), .C(w366) );
	io_NAND4 g_599 (.B(w367), .C(w341), .A(w355), .D(w342), .Z(w347) );
	io_DFFRPOS g_600 (.Q(w368), .nRES(1'b1), .D(w138), .C(w333) );
	io_NAND g_601 (.A(w344), .B(w480), .Z(w542) );
	io_DFFRPOS g_602 (.Q(w252), .nRES(w112), .D(w143), .C(w430) );
	io_NAND g_603 (.A(w343), .B(w480), .Z(w543) );
	io_NAND6 g_604 (.C(w543), .D(w347), .B(w542), .E(w338), .A(w544), .F(1'b1), .Z(w545) );
	io_NAND g_605 (.A(w480), .B(w349), .Z(w544) );
	io_DFFSPOS g_606 (.C(w366), .D(w545), .nSET(w365), .nQ(w355), .Q(w480) );
	io_DFFRPOS g_607 (.Q(w350), .nRES(1'b1), .D(w186), .C(w333) );
	io_NOT g_608 (.A(w351), .nZ(w310) );
	io_DFFRPOS g_609 (.Q(w351), .nRES(w112), .D(w336), .C(w430) );
	io_DFFRPOS g_610 (.Q(w352), .nRES(w112), .D(w130), .C(w430) );
	io_NOT g_611 (.A(w352), .nZ(w322) );
	io_BUF g_612 (.Z(w357), .A(w431) );
	io_DFFRPOS g_613 (.nQ(w354), .Q(w353), .nRES(w357), .D(w432), .C(w355) );
	io_DFFSPOS g_614 (.C(w355), .D(w356), .nSET(w357), .Q(w358) );
	io_OR g_615 (.A(w358), .Z(w436), .B(w355) );
	io_DFFRPOS g_616 (.nQ(w359), .Q(w360), .nRES(w435), .D(w361), .C(w362) );
	io_NAND4 g_617 (.B(w364), .C(w334), .A(w363), .D(w335), .Z(w361) );
	io_NAND3 g_618 (.A(w433), .B(w434), .C(w360), .Z(w335) );
	io_NAND3 g_619 (.A(w428), .B(w360), .C(w433), .Z(w334) );
	io_OR g_620 (.A(w325), .Z(w16), .B(w266) );
	io_DFFRPOS g_621 (.nQ(w409), .Q(w411), .nRES(w410), .D(w414), .C(w412) );
	io_DFFRPOS g_622 (.nQ(w415), .Q(w296), .nRES(w410), .D(w413), .C(w412) );
	io_NAND g_623 (.A(w411), .B(w296), .Z(w295) );
	io_NAND4 g_624 (.B(w417), .C(w294), .A(w416), .D(w295), .Z(w413) );
	io_NAND3 g_625 (.A(w420), .B(w417), .C(w294), .Z(w414) );
	io_NAND g_626 (.A(w419), .B(w411), .Z(w417) );
	io_NAND g_627 (.A(w419), .B(w296), .Z(w416) );
	io_NAND4 g_628 (.B(w418), .C(w329), .A(w409), .D(w296), .Z(w294) );
	io_DFFRPOS g_629 (.nQ(w418), .Q(w419), .nRES(w410), .D(w424), .C(w412) );
	io_NAND3 g_630 (.A(w415), .B(w411), .C(w419), .Z(w423) );
	io_NAND g_631 (.A(w418), .B(w296), .Z(w427) );
	io_NAND3 g_632 (.A(w423), .B(w420), .C(w427), .Z(w424) );
	io_NAND3 g_633 (.A(w419), .B(w329), .C(w296), .Z(w297) );
	io_NAND4 g_634 (.B(w423), .C(w298), .A(w420), .D(w297), .Z(w425) );
	io_NAND3 g_635 (.A(w411), .B(w329), .C(w296), .Z(w298) );
	io_DFFRPOS g_636 (.nQ(w382), .Q(w404), .nRES(w401), .D(w400), .C(w345) );
	io_NAND g_637 (.A(w397), .B(w404), .Z(w402) );
	io_NAND3 g_638 (.A(w402), .B(w403), .C(w395), .Z(w400) );
	io_DFFRPOS g_639 (.nQ(w383), .Q(w397), .nRES(w401), .D(w396), .C(w345) );
	io_NAND3 g_640 (.A(w392), .B(w398), .C(w395), .Z(w396) );
	io_NAND g_641 (.A(w383), .B(w393), .Z(w392) );
	io_AND g_642 (.Z(w399), .B(w390), .A(w394) );
	io_NOR g_643 (.Z(w391), .B(w300), .A(w399) );
	io_BUF g_644 (.Z(w119), .A(w391) );
	io_AND g_645 (.Z(w390), .B(1'b1), .A(w523) );
	io_DFFRPOS g_646 (.nQ(w326), .Q(w389), .nRES(w374), .D(w380), .C(w379) );
	io_DFFRPOS g_647 (.nQ(w328), .Q(w327), .nRES(w374), .D(w381), .C(w379) );
	io_NAND3 g_648 (.A(w372), .B(w389), .C(w371), .Z(w301) );
	io_NAND4 g_649 (.B(w376), .C(w301), .A(w378), .D(w299), .Z(w380) );
	io_NAND4 g_650 (.B(w371), .C(w326), .A(w377), .D(w327), .Z(w376) );
	io_NAND4 g_651 (.B(w299), .C(w302), .A(w378), .D(w303), .Z(w381) );
	io_NAND4 g_652 (.B(w377), .C(w326), .A(w371), .D(w328), .Z(w299) );
	io_NAND3 g_653 (.A(w377), .B(w389), .C(w371), .Z(w375) );
	io_NAND3 g_654 (.A(w371), .B(w327), .C(w389), .Z(w303) );
	io_NAND3 g_655 (.A(w372), .B(w327), .C(w371), .Z(w302) );
	io_NAND g_656 (.A(w343), .B(w349), .Z(w304) );
	io_NAND g_657 (.A(w349), .B(w344), .Z(w370) );
	io_NAND4 g_658 (.B(w370), .C(w304), .A(w338), .D(w305), .Z(w369) );
	io_DFFSPOS g_659 (.C(w366), .D(w369), .nSET(w365), .nQ(w367), .Q(w349) );
	io_NAND3 g_660 (.A(w342), .B(w341), .C(w367), .Z(w305) );
	io_DFFSPOS g_661 (.C(w366), .D(w339), .nSET(w365), .nQ(w342), .Q(w343) );
	io_NAND g_662 (.A(w341), .B(w342), .Z(w340) );
	io_NAND3 g_663 (.A(w337), .B(w338), .C(w340), .Z(w339) );
	io_NAND g_664 (.A(w344), .B(w343), .Z(w337) );
	io_MUX g_665 (.C(w324), .Z(w346), .A(w306), .B(w345) );
	io_NOT g_666 (.A(w293), .nZ(w121) );
	io_NOT g_667 (.A(w252), .nZ(w308) );
	io_DFFRPOS g_668 (.Q(w330), .nRES(1'b1), .D(w143), .C(w333) );
	io_DFFRPOS g_669 (.Q(w309), .nRES(1'b1), .D(w336), .C(w333) );
	io_DFFRPOS g_670 (.Q(w323), .nRES(1'b1), .D(w130), .C(w333) );
	io_DFFRPOS g_671 (.Q(w311), .nRES(1'b1), .D(w108), .C(w333) );
	io_DFFRPOS g_672 (.Q(w320), .nRES(1'b1), .D(w165), .C(w333) );
	io_DFFRPOS g_673 (.Q(w312), .nRES(1'b1), .D(w156), .C(w333) );
	io_DFFSPOS g_674 (.C(w12), .D(w186), .nSET(w122), .Q(w132) );
	io_RCDELAY g_675 (.A(w657), .Z(w654) );
	io_RCDELAY g_676 (.A(w690), .Z(w691) );
	io_RCDELAY g_677 (.A(w692), .Z(w689) );
	io_RCDELAY g_678 (.A(w656), .Z(w652) );
	io_RCDELAY g_679 (.A(w661), .Z(w703) );
	io_RCDELAY g_680 (.A(w748), .Z(w736) );
	io_RCDELAY g_681 (.A(w751), .Z(w750) );
	io_RCDELAY g_682 (.A(w842), .Z(w841) );
	io_RCDELAY g_683 (.A(w840), .Z(w846) );
	io_RCDELAY g_684 (.A(w749), .Z(w837) );
	io_RCDELAY g_685 (.A(w655), .Z(w843) );
	io_RCDELAY g_686 (.A(w834), .Z(w847) );
	io_RCDELAY g_687 (.A(w873), .Z(w864) );
	io_RCDELAY g_688 (.A(w850), .Z(w862) );
	io_RCDELAY g_689 (.A(w852), .Z(w851) );
	io_RCDELAY g_690 (.A(w274), .Z(w917) );
	io_RCDELAY g_691 (.A(w916), .Z(w915) );
	io_RCDELAY g_692 (.A(w914), .Z(w920) );
	io_RCDELAY g_693 (.A(w921), .Z(w908) );
	io_RCDELAY g_694 (.A(w922), .Z(w861) );
	io_RCDELAY g_695 (.A(w865), .Z(w927) );
	io_RCDELAY g_696 (.A(w909), .Z(w273) );
	io_RCDELAY g_697 (.A(w924), .Z(w900) );
	io_RCDELAY g_698 (.A(w667), .Z(w659) );
endmodule // IO

// Module Definitions [It is possible to wrap here on your primitives]

module io_AND (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // io_AND

module io_OR (  A, Z, B);

	input wire A;
	output wire Z;
	input wire B;

endmodule // io_OR

module io_NOR (  Z, B, A);

	output wire Z;
	input wire B;
	input wire A;

endmodule // io_NOR

module io_NOT (  A, nZ);

	input wire A;
	output wire nZ;

endmodule // io_NOT

module io_OR4 (  Z, D, C, B, A);

	output wire Z;
	input wire D;
	input wire C;
	input wire B;
	input wire A;

endmodule // io_OR4

module io_OR3 (  Z, C, B, A);

	output wire Z;
	input wire C;
	input wire B;
	input wire A;

endmodule // io_OR3

module io_NAND (  A, B, Z);

	input wire A;
	input wire B;
	output wire Z;

endmodule // io_NAND

module io_NAND8 (  Z, D, C, B, A, E, F, G, H);

	output wire Z;
	input wire D;
	input wire C;
	input wire B;
	input wire A;
	input wire E;
	input wire F;
	input wire G;
	input wire H;

endmodule // io_NAND8

module io_AND3 (  Z, C, B, A);

	output wire Z;
	input wire C;
	input wire B;
	input wire A;

endmodule // io_AND3

module io_NOR3 (  Z, C, B, A);

	output wire Z;
	input wire C;
	input wire B;
	input wire A;

endmodule // io_NOR3

module io_DFFRPOS (  nQ, Q, nRES, D, C);

	output wire nQ;
	output wire Q;
	input wire nRES;
	input wire D;
	input wire C;

endmodule // io_DFFRPOS

module io_MUX4BIT (  S, Z0, A0, B0, A1, B1, Z1, Z2, B2, A2, A3, B3, Z3);

	input wire S;
	output wire Z0;
	input wire A0;
	input wire B0;
	input wire A1;
	input wire B1;
	output wire Z1;
	output wire Z2;
	input wire B2;
	input wire A2;
	input wire A3;
	input wire B3;
	output wire Z3;

endmodule // io_MUX4BIT

module io_DFFSPOS (  C, D, nSET, nQ, Q);

	input wire C;
	input wire D;
	input wire nSET;
	output wire nQ;
	output wire Q;

endmodule // io_DFFSPOS

module io_NOR4 (  Z, D, C, B, A);

	output wire Z;
	input wire D;
	input wire C;
	input wire B;
	input wire A;

endmodule // io_NOR4

module io_NAND4 (  B, C, A, D, Z);

	input wire B;
	input wire C;
	input wire A;
	input wire D;
	output wire Z;

endmodule // io_NAND4

module io_CNT_BIT (  Q, nQ, C, nRES, D, nLD, CO, CI);

	output wire Q;
	output wire nQ;
	input wire C;
	input wire nRES;
	input wire D;
	input wire nLD;
	output wire CO;
	input wire CI;

endmodule // io_CNT_BIT

module io_MUX8TO1 (  S0, S2, S1, G, H, F, E, Z, C, D, B, A);

	input wire S0;
	input wire S2;
	input wire S1;
	input wire G;
	input wire H;
	input wire F;
	input wire E;
	output wire Z;
	input wire C;
	input wire D;
	input wire B;
	input wire A;

endmodule // io_MUX8TO1

module io_SIPO_4BIT (  C, D, nRES, Q0, Q1, Q2, Q3);

	input wire C;
	input wire D;
	input wire nRES;
	output wire Q0;
	output wire Q1;
	output wire Q2;
	output wire Q3;

endmodule // io_SIPO_4BIT

module io_BUF (  Z, A);

	output wire Z;
	input wire A;

endmodule // io_BUF

module io_AON22 (  Z, B2, A2, B1, A1);

	output wire Z;
	input wire B2;
	input wire A2;
	input wire B1;
	input wire A1;

endmodule // io_AON22

module io_NOR6 (  Z, F, E, D, C, B, A);

	output wire Z;
	input wire F;
	input wire E;
	input wire D;
	input wire C;
	input wire B;
	input wire A;

endmodule // io_NOR6

module io_TFF (  nQ, Q, T, C);

	output wire nQ;
	output wire Q;
	input wire T;
	input wire C;

endmodule // io_TFF

module io_MUX (  C, Z, A, B);

	input wire C;
	output wire Z;
	input wire A;
	input wire B;

endmodule // io_MUX

module io_SLATCH (  nQ, C, Q, D);

	output wire nQ;
	input wire C;
	output wire Q;
	input wire D;

endmodule // io_SLATCH

module io_MUX2BIT4TO1 (  A0, A1, ZA, A3, A2, B0, B1, ZB, B3, B2, S1, S0);

	input wire A0;
	input wire A1;
	output wire ZA;
	input wire A3;
	input wire A2;
	input wire B0;
	input wire B1;
	output wire ZB;
	input wire B3;
	input wire B2;
	input wire S1;
	input wire S0;

endmodule // io_MUX2BIT4TO1

module io_XNOR (  A, B, Z);

	input wire A;
	input wire B;
	output wire Z;

endmodule // io_XNOR

module io_JKFFSRNEG (  C, K, J, nSET, nRES, Q, nQ);

	input wire C;
	input wire K;
	input wire J;
	input wire nSET;
	input wire nRES;
	output wire Q;
	output wire nQ;

endmodule // io_JKFFSRNEG

module io_NAND6 (  C, D, B, E, A, F, Z);

	input wire C;
	input wire D;
	input wire B;
	input wire E;
	input wire A;
	input wire F;
	output wire Z;

endmodule // io_NAND6

module io_NAND3 (  A, B, C, Z);

	input wire A;
	input wire B;
	input wire C;
	output wire Z;

endmodule // io_NAND3

module io_DFFSRPOS (  C, D, nRES, nQ, nSET, Q);

	input wire C;
	input wire D;
	input wire nRES;
	output wire nQ;
	input wire nSET;
	output wire Q;

endmodule // io_DFFSRPOS

module io_DFFPOS (  nQ, Q, D, C);

	output wire nQ;
	output wire Q;
	input wire D;
	input wire C;

endmodule // io_DFFPOS

module io_RCDELAY (  A, Z);

	input wire A;
	output wire Z;

endmodule // io_RCDELAY



// ERROR: floating wire w19
// ERROR: floating wire w34
// ERROR: floating wire w78
// ERROR: floating wire w87
// ERROR: floating wire w89
// ERROR: floating wire w114
// ERROR: floating wire w177
// ERROR: floating wire w185
// ERROR: floating wire w187
// ERROR: floating wire w220
// ERROR: floating wire w332
// ERROR: floating wire w348
// ERROR: floating wire w385
// ERROR: floating wire w464
// ERROR: floating wire w504
// ERROR: floating wire w521
// ERROR: floating wire w525
// ERROR: floating wire w535
// ERROR: floating wire w537
// ERROR: floating wire w562
// ERROR: floating wire w585
// ERROR: floating wire w606
// ERROR: floating wire w616
// ERROR: floating wire w662
// ERROR: floating wire w694
// ERROR: floating wire w697
// ERROR: floating wire w714
// ERROR: floating wire w715
// ERROR: floating wire w798
// ERROR: floating wire w799
// ERROR: floating wire w923
// WARNING: Cell io_DFFRPOS:g_17 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_18 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_20 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_21 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_26 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_27 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_29 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_30 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_36 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_38 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_39 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_40 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_42 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_42 port Q not connected.
// WARNING: Cell io_MUX4BIT:g_43 port Z0 not connected.
// WARNING: Cell io_DFFRPOS:g_44 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_44 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_47 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_48 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_49 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_49 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_50 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_50 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_51 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_51 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_52 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_52 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_53 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_53 port Q not connected.
// WARNING: Cell io_NAND4:g_54 port Z not connected.
// WARNING: Cell io_NAND4:g_57 port Z not connected.
// WARNING: Cell io_NAND4:g_59 port Z not connected.
// WARNING: Cell io_NAND4:g_61 port Z not connected.
// WARNING: Cell io_NAND4:g_63 port Z not connected.
// WARNING: Cell io_CNT_BIT:g_78 port Q not connected.
// WARNING: Cell io_CNT_BIT:g_78 port CO not connected.
// WARNING: Cell io_CNT_BIT:g_80 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_82 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_83 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_84 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_85 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_87 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_93 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_95 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_98 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_99 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_100 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_105 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_106 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_113 port nQ not connected.
// WARNING: Cell io_CNT_BIT:g_129 port Q not connected.
// WARNING: Cell io_CNT_BIT:g_130 port Q not connected.
// WARNING: Cell io_CNT_BIT:g_133 port Q not connected.
// WARNING: Cell io_CNT_BIT:g_134 port Q not connected.
// WARNING: Cell io_CNT_BIT:g_134 port CO not connected.
// WARNING: Cell io_DFFSPOS:g_139 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_140 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_142 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_143 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_145 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_146 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_150 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_151 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_152 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_153 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_154 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_154 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_155 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_156 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_159 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_160 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_164 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_164 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_165 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_166 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_177 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_179 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_182 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_183 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_184 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_185 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_186 port nQ not connected.
// WARNING: Cell io_CNT_BIT:g_188 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_189 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_190 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_191 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_192 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_193 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_194 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_195 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_197 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_200 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_202 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_208 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_210 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_211 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_213 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_214 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_215 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_216 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_220 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_229 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_231 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_234 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_236 port nQ not connected.
// WARNING: Cell io_TFF:g_238 port nQ not connected.
// WARNING: Cell io_TFF:g_239 port nQ not connected.
// WARNING: Cell io_TFF:g_240 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_241 port nQ not connected.
// WARNING: Cell io_TFF:g_243 port nQ not connected.
// WARNING: Cell io_TFF:g_244 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_261 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_272 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_273 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_274 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_277 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_278 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_280 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_281 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_302 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_312 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_314 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_315 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_316 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_318 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_320 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_321 port nQ not connected.
// WARNING: Cell io_NAND4:g_333 port Z not connected.
// WARNING: Cell io_DFFRPOS:g_340 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_344 port nQ not connected.
// WARNING: Cell io_TFF:g_345 port nQ not connected.
// WARNING: Cell io_TFF:g_346 port nQ not connected.
// WARNING: Cell io_TFF:g_347 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_353 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_355 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_358 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_360 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_371 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_377 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_379 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_389 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_390 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_391 port nQ not connected.
// WARNING: Cell io_NAND4:g_399 port Z not connected.
// WARNING: Cell io_NAND4:g_402 port Z not connected.
// WARNING: Cell io_NAND4:g_405 port Z not connected.
// WARNING: Cell io_DFFSPOS:g_408 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_419 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_425 port Q not connected.
// WARNING: Cell io_DFFSRPOS:g_426 port nQ not connected.
// WARNING: Cell io_DFFPOS:g_429 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_434 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_436 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_438 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_442 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_443 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_446 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_448 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_451 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_452 port nQ not connected.
// WARNING: Cell io_DFFSRPOS:g_457 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_459 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_461 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_462 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_467 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_498 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_502 port nQ not connected.
// WARNING: Cell io_DFFSRPOS:g_504 port nQ not connected.
// WARNING: Cell io_DFFPOS:g_507 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_509 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_513 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_517 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_522 port Q not connected.
// WARNING: Cell io_DFFRPOS:g_526 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_528 port nQ not connected.
// WARNING: Cell io_DFFPOS:g_577 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_600 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_602 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_607 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_609 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_610 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_614 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_668 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_669 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_670 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_671 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_672 port nQ not connected.
// WARNING: Cell io_DFFRPOS:g_673 port nQ not connected.
// WARNING: Cell io_DFFSPOS:g_674 port nQ not connected.
